/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sat Apr 25 22:33:22 2020
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 2363246184 */

module datapath(R, L, plus);
   input [30:0]R;
   input [30:0]L;
   output [30:0]plus;

   HA_X1 i_1 (.A(R[0]), .B(L[0]), .CO(n_2), .S(n_1));
   FA_X1 i_2 (.A(R[1]), .B(L[1]), .CI(n_2), .CO(n_3), .S(plus[1]));
   FA_X1 i_3 (.A(R[2]), .B(L[2]), .CI(n_3), .CO(n_4), .S(plus[2]));
   FA_X1 i_4 (.A(R[3]), .B(L[3]), .CI(n_4), .CO(n_5), .S(plus[3]));
   FA_X1 i_5 (.A(R[4]), .B(L[4]), .CI(n_5), .CO(n_6), .S(plus[4]));
   FA_X1 i_6 (.A(R[5]), .B(L[5]), .CI(n_6), .CO(n_7), .S(plus[5]));
   FA_X1 i_7 (.A(R[6]), .B(L[6]), .CI(n_7), .CO(n_8), .S(plus[6]));
   FA_X1 i_8 (.A(R[7]), .B(L[7]), .CI(n_8), .CO(n_9), .S(plus[7]));
   FA_X1 i_9 (.A(R[8]), .B(L[8]), .CI(n_9), .CO(n_10), .S(plus[8]));
   FA_X1 i_10 (.A(R[9]), .B(L[9]), .CI(n_10), .CO(n_11), .S(plus[9]));
   FA_X1 i_11 (.A(R[10]), .B(L[10]), .CI(n_11), .CO(n_12), .S(plus[10]));
   FA_X1 i_12 (.A(R[11]), .B(L[11]), .CI(n_12), .CO(n_13), .S(plus[11]));
   FA_X1 i_13 (.A(R[12]), .B(L[12]), .CI(n_13), .CO(n_14), .S(plus[12]));
   FA_X1 i_14 (.A(R[13]), .B(L[13]), .CI(n_14), .CO(n_15), .S(plus[13]));
   XNOR2_X1 i_0 (.A(n_15), .B(n_0), .ZN(plus[14]));
   XNOR2_X1 i_15 (.A(R[14]), .B(L[14]), .ZN(n_0));
   XOR2_X1 i_16 (.A(R[15]), .B(n_16), .Z(plus[15]));
   NAND2_X1 i_17 (.A1(n_19), .A2(n_18), .ZN(n_16));
   NAND2_X1 i_18 (.A1(n_18), .A2(n_17), .ZN(plus[30]));
   NAND2_X1 i_19 (.A1(n_19), .A2(R[15]), .ZN(n_17));
   OR3_X1 i_20 (.A1(n_20), .A2(n_15), .A3(R[14]), .ZN(n_18));
   NAND3_X1 i_21 (.A1(n_20), .A2(n_15), .A3(R[14]), .ZN(n_19));
   INV_X1 i_22 (.A(L[14]), .ZN(n_20));
endmodule

module datapath__0_9(R, L, plus);
   input [29:0]R;
   input [29:0]L;
   output [29:0]plus;

   INV_X1 i_0 (.A(R[15]), .ZN(n_0));
   INV_X1 i_1 (.A(L[29]), .ZN(n_1));
   HA_X1 i_2 (.A(R[0]), .B(L[0]), .CO(n_3), .S(n_2));
   FA_X1 i_3 (.A(R[1]), .B(L[1]), .CI(n_3), .CO(n_4), .S(plus[1]));
   FA_X1 i_4 (.A(R[2]), .B(L[2]), .CI(n_4), .CO(n_5), .S(plus[2]));
   FA_X1 i_5 (.A(R[3]), .B(L[3]), .CI(n_5), .CO(n_6), .S(plus[3]));
   FA_X1 i_6 (.A(R[4]), .B(L[4]), .CI(n_6), .CO(n_7), .S(plus[4]));
   FA_X1 i_7 (.A(R[5]), .B(L[5]), .CI(n_7), .CO(n_8), .S(plus[5]));
   FA_X1 i_8 (.A(R[6]), .B(L[6]), .CI(n_8), .CO(n_9), .S(plus[6]));
   FA_X1 i_9 (.A(R[7]), .B(L[7]), .CI(n_9), .CO(n_10), .S(plus[7]));
   FA_X1 i_10 (.A(R[8]), .B(L[8]), .CI(n_10), .CO(n_11), .S(plus[8]));
   FA_X1 i_11 (.A(R[9]), .B(L[9]), .CI(n_11), .CO(n_12), .S(plus[9]));
   FA_X1 i_12 (.A(R[10]), .B(L[10]), .CI(n_12), .CO(n_13), .S(plus[10]));
   FA_X1 i_13 (.A(R[11]), .B(L[11]), .CI(n_13), .CO(n_14), .S(plus[11]));
   FA_X1 i_14 (.A(R[12]), .B(L[12]), .CI(n_14), .CO(n_15), .S(plus[12]));
   FA_X1 i_15 (.A(R[13]), .B(L[13]), .CI(n_15), .CO(n_16), .S(plus[13]));
   FA_X1 i_16 (.A(R[14]), .B(L[14]), .CI(n_16), .CO(n_17), .S(plus[14]));
   FA_X1 i_17 (.A(L[29]), .B(R[15]), .CI(n_17), .CO(n_18), .S(plus[15]));
   FA_X1 i_18 (.A(n_0), .B(n_1), .CI(n_18), .CO(n_19), .S(plus[16]));
   INV_X1 i_19 (.A(n_19), .ZN(plus[29]));
endmodule

module datapath__0_13(R, L, plus);
   input [28:0]R;
   input [28:0]L;
   output [28:0]plus;

   INV_X1 i_0 (.A(R[15]), .ZN(n_0));
   INV_X1 i_1 (.A(L[28]), .ZN(n_1));
   HA_X1 i_2 (.A(R[0]), .B(L[0]), .CO(n_3), .S(n_2));
   FA_X1 i_3 (.A(R[1]), .B(L[1]), .CI(n_3), .CO(n_4), .S(plus[1]));
   FA_X1 i_4 (.A(R[2]), .B(L[2]), .CI(n_4), .CO(n_5), .S(plus[2]));
   FA_X1 i_5 (.A(R[3]), .B(L[3]), .CI(n_5), .CO(n_6), .S(plus[3]));
   FA_X1 i_6 (.A(R[4]), .B(L[4]), .CI(n_6), .CO(n_7), .S(plus[4]));
   FA_X1 i_7 (.A(R[5]), .B(L[5]), .CI(n_7), .CO(n_8), .S(plus[5]));
   FA_X1 i_8 (.A(R[6]), .B(L[6]), .CI(n_8), .CO(n_9), .S(plus[6]));
   FA_X1 i_9 (.A(R[7]), .B(L[7]), .CI(n_9), .CO(n_10), .S(plus[7]));
   FA_X1 i_10 (.A(R[8]), .B(L[8]), .CI(n_10), .CO(n_11), .S(plus[8]));
   FA_X1 i_11 (.A(R[9]), .B(L[9]), .CI(n_11), .CO(n_12), .S(plus[9]));
   FA_X1 i_12 (.A(R[10]), .B(L[10]), .CI(n_12), .CO(n_13), .S(plus[10]));
   FA_X1 i_13 (.A(R[11]), .B(L[11]), .CI(n_13), .CO(n_14), .S(plus[11]));
   FA_X1 i_14 (.A(R[12]), .B(L[12]), .CI(n_14), .CO(n_15), .S(plus[12]));
   FA_X1 i_15 (.A(R[13]), .B(L[13]), .CI(n_15), .CO(n_16), .S(plus[13]));
   FA_X1 i_16 (.A(R[14]), .B(L[14]), .CI(n_16), .CO(n_17), .S(plus[14]));
   FA_X1 i_17 (.A(L[15]), .B(R[15]), .CI(n_17), .CO(n_18), .S(plus[15]));
   FA_X1 i_18 (.A(n_0), .B(n_1), .CI(n_18), .CO(n_19), .S(plus[16]));
   INV_X1 i_19 (.A(n_19), .ZN(plus[28]));
endmodule

module datapath__0_17(R, L, plus);
   input [27:0]R;
   input [27:0]L;
   output [27:0]plus;

   INV_X1 i_0 (.A(R[15]), .ZN(n_0));
   INV_X1 i_1 (.A(L[27]), .ZN(n_1));
   HA_X1 i_2 (.A(R[0]), .B(L[0]), .CO(n_3), .S(n_2));
   FA_X1 i_3 (.A(R[1]), .B(L[1]), .CI(n_3), .CO(n_4), .S(plus[1]));
   FA_X1 i_4 (.A(R[2]), .B(L[2]), .CI(n_4), .CO(n_5), .S(plus[2]));
   FA_X1 i_5 (.A(R[3]), .B(L[3]), .CI(n_5), .CO(n_6), .S(plus[3]));
   FA_X1 i_6 (.A(R[4]), .B(L[4]), .CI(n_6), .CO(n_7), .S(plus[4]));
   FA_X1 i_7 (.A(R[5]), .B(L[5]), .CI(n_7), .CO(n_8), .S(plus[5]));
   FA_X1 i_8 (.A(R[6]), .B(L[6]), .CI(n_8), .CO(n_9), .S(plus[6]));
   FA_X1 i_9 (.A(R[7]), .B(L[7]), .CI(n_9), .CO(n_10), .S(plus[7]));
   FA_X1 i_10 (.A(R[8]), .B(L[8]), .CI(n_10), .CO(n_11), .S(plus[8]));
   FA_X1 i_11 (.A(R[9]), .B(L[9]), .CI(n_11), .CO(n_12), .S(plus[9]));
   FA_X1 i_12 (.A(R[10]), .B(L[10]), .CI(n_12), .CO(n_13), .S(plus[10]));
   FA_X1 i_13 (.A(R[11]), .B(L[11]), .CI(n_13), .CO(n_14), .S(plus[11]));
   FA_X1 i_14 (.A(R[12]), .B(L[12]), .CI(n_14), .CO(n_15), .S(plus[12]));
   FA_X1 i_15 (.A(R[13]), .B(L[13]), .CI(n_15), .CO(n_16), .S(plus[13]));
   FA_X1 i_16 (.A(R[14]), .B(L[14]), .CI(n_16), .CO(n_17), .S(plus[14]));
   FA_X1 i_17 (.A(L[15]), .B(R[15]), .CI(n_17), .CO(n_18), .S(plus[15]));
   FA_X1 i_18 (.A(n_0), .B(n_1), .CI(n_18), .CO(n_19), .S(plus[16]));
   INV_X1 i_19 (.A(n_19), .ZN(plus[27]));
endmodule

module datapath__0_21(R, L, plus);
   input [26:0]R;
   input [26:0]L;
   output [26:0]plus;

   INV_X1 i_0 (.A(R[15]), .ZN(n_0));
   INV_X1 i_1 (.A(L[26]), .ZN(n_1));
   HA_X1 i_2 (.A(R[0]), .B(L[0]), .CO(n_3), .S(n_2));
   FA_X1 i_3 (.A(R[1]), .B(L[1]), .CI(n_3), .CO(n_4), .S(plus[1]));
   FA_X1 i_4 (.A(R[2]), .B(L[2]), .CI(n_4), .CO(n_5), .S(plus[2]));
   FA_X1 i_5 (.A(R[3]), .B(L[3]), .CI(n_5), .CO(n_6), .S(plus[3]));
   FA_X1 i_6 (.A(R[4]), .B(L[4]), .CI(n_6), .CO(n_7), .S(plus[4]));
   FA_X1 i_7 (.A(R[5]), .B(L[5]), .CI(n_7), .CO(n_8), .S(plus[5]));
   FA_X1 i_8 (.A(R[6]), .B(L[6]), .CI(n_8), .CO(n_9), .S(plus[6]));
   FA_X1 i_9 (.A(R[7]), .B(L[7]), .CI(n_9), .CO(n_10), .S(plus[7]));
   FA_X1 i_10 (.A(R[8]), .B(L[8]), .CI(n_10), .CO(n_11), .S(plus[8]));
   FA_X1 i_11 (.A(R[9]), .B(L[9]), .CI(n_11), .CO(n_12), .S(plus[9]));
   FA_X1 i_12 (.A(R[10]), .B(L[10]), .CI(n_12), .CO(n_13), .S(plus[10]));
   FA_X1 i_13 (.A(R[11]), .B(L[11]), .CI(n_13), .CO(n_14), .S(plus[11]));
   FA_X1 i_14 (.A(R[12]), .B(L[12]), .CI(n_14), .CO(n_15), .S(plus[12]));
   FA_X1 i_15 (.A(R[13]), .B(L[13]), .CI(n_15), .CO(n_16), .S(plus[13]));
   FA_X1 i_16 (.A(R[14]), .B(L[14]), .CI(n_16), .CO(n_17), .S(plus[14]));
   FA_X1 i_17 (.A(L[15]), .B(R[15]), .CI(n_17), .CO(n_18), .S(plus[15]));
   FA_X1 i_18 (.A(n_0), .B(n_1), .CI(n_18), .CO(n_19), .S(plus[16]));
   INV_X1 i_19 (.A(n_19), .ZN(plus[26]));
endmodule

module datapath__0_25(R, L, plus);
   input [25:0]R;
   input [25:0]L;
   output [25:0]plus;

   INV_X1 i_0 (.A(R[15]), .ZN(n_0));
   INV_X1 i_1 (.A(L[25]), .ZN(n_1));
   HA_X1 i_2 (.A(R[0]), .B(L[0]), .CO(n_3), .S(n_2));
   FA_X1 i_3 (.A(R[1]), .B(L[1]), .CI(n_3), .CO(n_4), .S(plus[1]));
   FA_X1 i_4 (.A(R[2]), .B(L[2]), .CI(n_4), .CO(n_5), .S(plus[2]));
   FA_X1 i_5 (.A(R[3]), .B(L[3]), .CI(n_5), .CO(n_6), .S(plus[3]));
   FA_X1 i_6 (.A(R[4]), .B(L[4]), .CI(n_6), .CO(n_7), .S(plus[4]));
   FA_X1 i_7 (.A(R[5]), .B(L[5]), .CI(n_7), .CO(n_8), .S(plus[5]));
   FA_X1 i_8 (.A(R[6]), .B(L[6]), .CI(n_8), .CO(n_9), .S(plus[6]));
   FA_X1 i_9 (.A(R[7]), .B(L[7]), .CI(n_9), .CO(n_10), .S(plus[7]));
   FA_X1 i_10 (.A(R[8]), .B(L[8]), .CI(n_10), .CO(n_11), .S(plus[8]));
   FA_X1 i_11 (.A(R[9]), .B(L[9]), .CI(n_11), .CO(n_12), .S(plus[9]));
   FA_X1 i_12 (.A(R[10]), .B(L[10]), .CI(n_12), .CO(n_13), .S(plus[10]));
   FA_X1 i_13 (.A(R[11]), .B(L[11]), .CI(n_13), .CO(n_14), .S(plus[11]));
   FA_X1 i_14 (.A(R[12]), .B(L[12]), .CI(n_14), .CO(n_15), .S(plus[12]));
   FA_X1 i_15 (.A(R[13]), .B(L[13]), .CI(n_15), .CO(n_16), .S(plus[13]));
   FA_X1 i_16 (.A(R[14]), .B(L[14]), .CI(n_16), .CO(n_17), .S(plus[14]));
   FA_X1 i_17 (.A(L[15]), .B(R[15]), .CI(n_17), .CO(n_18), .S(plus[15]));
   FA_X1 i_18 (.A(n_0), .B(n_1), .CI(n_18), .CO(n_19), .S(plus[16]));
   INV_X1 i_19 (.A(n_19), .ZN(plus[25]));
endmodule

module datapath__0_29(R, L, plus);
   input [24:0]R;
   input [24:0]L;
   output [24:0]plus;

   INV_X1 i_0 (.A(R[15]), .ZN(n_0));
   INV_X1 i_1 (.A(L[24]), .ZN(n_1));
   HA_X1 i_2 (.A(R[0]), .B(L[0]), .CO(n_2), .S(plus[0]));
   FA_X1 i_3 (.A(R[1]), .B(L[1]), .CI(n_2), .CO(n_3), .S(plus[1]));
   FA_X1 i_4 (.A(R[2]), .B(L[2]), .CI(n_3), .CO(n_4), .S(plus[2]));
   FA_X1 i_5 (.A(R[3]), .B(L[3]), .CI(n_4), .CO(n_5), .S(plus[3]));
   FA_X1 i_6 (.A(R[4]), .B(L[4]), .CI(n_5), .CO(n_6), .S(plus[4]));
   FA_X1 i_7 (.A(R[5]), .B(L[5]), .CI(n_6), .CO(n_7), .S(plus[5]));
   FA_X1 i_8 (.A(R[6]), .B(L[6]), .CI(n_7), .CO(n_8), .S(plus[6]));
   FA_X1 i_9 (.A(R[7]), .B(L[7]), .CI(n_8), .CO(n_9), .S(plus[7]));
   FA_X1 i_10 (.A(R[8]), .B(L[8]), .CI(n_9), .CO(n_10), .S(plus[8]));
   FA_X1 i_11 (.A(R[9]), .B(L[9]), .CI(n_10), .CO(n_11), .S(plus[9]));
   FA_X1 i_12 (.A(R[10]), .B(L[10]), .CI(n_11), .CO(n_12), .S(plus[10]));
   FA_X1 i_13 (.A(R[11]), .B(L[11]), .CI(n_12), .CO(n_13), .S(plus[11]));
   FA_X1 i_14 (.A(R[12]), .B(L[12]), .CI(n_13), .CO(n_14), .S(plus[12]));
   FA_X1 i_15 (.A(R[13]), .B(L[13]), .CI(n_14), .CO(n_15), .S(plus[13]));
   FA_X1 i_16 (.A(R[14]), .B(L[14]), .CI(n_15), .CO(n_16), .S(plus[14]));
   FA_X1 i_17 (.A(L[15]), .B(R[15]), .CI(n_16), .CO(n_17), .S(plus[15]));
   FA_X1 i_18 (.A(n_0), .B(n_1), .CI(n_17), .CO(n_18), .S(plus[16]));
   INV_X1 i_19 (.A(n_18), .ZN(plus[24]));
endmodule

module datapath__0_33(R, L, plus);
   input [23:0]R;
   input [23:0]L;
   output [23:0]plus;

   INV_X1 i_0 (.A(R[15]), .ZN(n_0));
   INV_X1 i_1 (.A(L[23]), .ZN(n_1));
   HA_X1 i_2 (.A(R[0]), .B(L[0]), .CO(n_2), .S(plus[0]));
   FA_X1 i_3 (.A(R[1]), .B(L[1]), .CI(n_2), .CO(n_3), .S(plus[1]));
   FA_X1 i_4 (.A(R[2]), .B(L[2]), .CI(n_3), .CO(n_4), .S(plus[2]));
   FA_X1 i_5 (.A(R[3]), .B(L[3]), .CI(n_4), .CO(n_5), .S(plus[3]));
   FA_X1 i_6 (.A(R[4]), .B(L[4]), .CI(n_5), .CO(n_6), .S(plus[4]));
   FA_X1 i_7 (.A(R[5]), .B(L[5]), .CI(n_6), .CO(n_7), .S(plus[5]));
   FA_X1 i_8 (.A(R[6]), .B(L[6]), .CI(n_7), .CO(n_8), .S(plus[6]));
   FA_X1 i_9 (.A(R[7]), .B(L[7]), .CI(n_8), .CO(n_9), .S(plus[7]));
   FA_X1 i_10 (.A(R[8]), .B(L[8]), .CI(n_9), .CO(n_10), .S(plus[8]));
   FA_X1 i_11 (.A(R[9]), .B(L[9]), .CI(n_10), .CO(n_11), .S(plus[9]));
   FA_X1 i_12 (.A(R[10]), .B(L[10]), .CI(n_11), .CO(n_12), .S(plus[10]));
   FA_X1 i_13 (.A(R[11]), .B(L[11]), .CI(n_12), .CO(n_13), .S(plus[11]));
   FA_X1 i_14 (.A(R[12]), .B(L[12]), .CI(n_13), .CO(n_14), .S(plus[12]));
   FA_X1 i_15 (.A(R[13]), .B(L[13]), .CI(n_14), .CO(n_15), .S(plus[13]));
   FA_X1 i_16 (.A(R[14]), .B(L[14]), .CI(n_15), .CO(n_16), .S(plus[14]));
   FA_X1 i_17 (.A(L[15]), .B(R[15]), .CI(n_16), .CO(n_17), .S(plus[15]));
   FA_X1 i_18 (.A(n_0), .B(n_1), .CI(n_17), .CO(n_18), .S(plus[16]));
   INV_X1 i_19 (.A(n_18), .ZN(plus[23]));
endmodule

module datapath__0_37(R, L, plus);
   input [22:0]R;
   input [22:0]L;
   output [22:0]plus;

   INV_X1 i_0 (.A(R[15]), .ZN(n_0));
   INV_X1 i_1 (.A(L[22]), .ZN(n_1));
   HA_X1 i_2 (.A(R[0]), .B(L[0]), .CO(n_2), .S(plus[0]));
   FA_X1 i_3 (.A(R[1]), .B(L[1]), .CI(n_2), .CO(n_3), .S(plus[1]));
   FA_X1 i_4 (.A(R[2]), .B(L[2]), .CI(n_3), .CO(n_4), .S(plus[2]));
   FA_X1 i_5 (.A(R[3]), .B(L[3]), .CI(n_4), .CO(n_5), .S(plus[3]));
   FA_X1 i_6 (.A(R[4]), .B(L[4]), .CI(n_5), .CO(n_6), .S(plus[4]));
   FA_X1 i_7 (.A(R[5]), .B(L[5]), .CI(n_6), .CO(n_7), .S(plus[5]));
   FA_X1 i_8 (.A(R[6]), .B(L[6]), .CI(n_7), .CO(n_8), .S(plus[6]));
   FA_X1 i_9 (.A(R[7]), .B(L[7]), .CI(n_8), .CO(n_9), .S(plus[7]));
   FA_X1 i_10 (.A(R[8]), .B(L[8]), .CI(n_9), .CO(n_10), .S(plus[8]));
   FA_X1 i_11 (.A(R[9]), .B(L[9]), .CI(n_10), .CO(n_11), .S(plus[9]));
   FA_X1 i_12 (.A(R[10]), .B(L[10]), .CI(n_11), .CO(n_12), .S(plus[10]));
   FA_X1 i_13 (.A(R[11]), .B(L[11]), .CI(n_12), .CO(n_13), .S(plus[11]));
   FA_X1 i_14 (.A(R[12]), .B(L[12]), .CI(n_13), .CO(n_14), .S(plus[12]));
   FA_X1 i_15 (.A(R[13]), .B(L[13]), .CI(n_14), .CO(n_15), .S(plus[13]));
   FA_X1 i_16 (.A(R[14]), .B(L[14]), .CI(n_15), .CO(n_16), .S(plus[14]));
   FA_X1 i_17 (.A(L[15]), .B(R[15]), .CI(n_16), .CO(n_17), .S(plus[15]));
   FA_X1 i_18 (.A(n_0), .B(n_1), .CI(n_17), .CO(n_18), .S(plus[16]));
   INV_X1 i_19 (.A(n_18), .ZN(plus[22]));
endmodule

module datapath__0_41(R, L, plus);
   input [21:0]R;
   input [21:0]L;
   output [21:0]plus;

   INV_X1 i_0 (.A(R[15]), .ZN(n_0));
   INV_X1 i_1 (.A(L[21]), .ZN(n_1));
   HA_X1 i_2 (.A(R[0]), .B(L[0]), .CO(n_2), .S(plus[0]));
   FA_X1 i_3 (.A(R[1]), .B(L[1]), .CI(n_2), .CO(n_3), .S(plus[1]));
   FA_X1 i_4 (.A(R[2]), .B(L[2]), .CI(n_3), .CO(n_4), .S(plus[2]));
   FA_X1 i_5 (.A(R[3]), .B(L[3]), .CI(n_4), .CO(n_5), .S(plus[3]));
   FA_X1 i_6 (.A(R[4]), .B(L[4]), .CI(n_5), .CO(n_6), .S(plus[4]));
   FA_X1 i_7 (.A(R[5]), .B(L[5]), .CI(n_6), .CO(n_7), .S(plus[5]));
   FA_X1 i_8 (.A(R[6]), .B(L[6]), .CI(n_7), .CO(n_8), .S(plus[6]));
   FA_X1 i_9 (.A(R[7]), .B(L[7]), .CI(n_8), .CO(n_9), .S(plus[7]));
   FA_X1 i_10 (.A(R[8]), .B(L[8]), .CI(n_9), .CO(n_10), .S(plus[8]));
   FA_X1 i_11 (.A(R[9]), .B(L[9]), .CI(n_10), .CO(n_11), .S(plus[9]));
   FA_X1 i_12 (.A(R[10]), .B(L[10]), .CI(n_11), .CO(n_12), .S(plus[10]));
   FA_X1 i_13 (.A(R[11]), .B(L[11]), .CI(n_12), .CO(n_13), .S(plus[11]));
   FA_X1 i_14 (.A(R[12]), .B(L[12]), .CI(n_13), .CO(n_14), .S(plus[12]));
   FA_X1 i_15 (.A(R[13]), .B(L[13]), .CI(n_14), .CO(n_15), .S(plus[13]));
   FA_X1 i_16 (.A(R[14]), .B(L[14]), .CI(n_15), .CO(n_16), .S(plus[14]));
   FA_X1 i_17 (.A(L[15]), .B(R[15]), .CI(n_16), .CO(n_17), .S(plus[15]));
   FA_X1 i_18 (.A(n_0), .B(n_1), .CI(n_17), .CO(n_18), .S(plus[16]));
   INV_X1 i_19 (.A(n_18), .ZN(plus[21]));
endmodule

module datapath__0_45(R, L, plus);
   input [20:0]R;
   input [20:0]L;
   output [20:0]plus;

   INV_X1 i_0 (.A(R[15]), .ZN(n_0));
   INV_X1 i_1 (.A(L[20]), .ZN(n_1));
   HA_X1 i_2 (.A(R[0]), .B(L[0]), .CO(n_2), .S(plus[0]));
   FA_X1 i_3 (.A(R[1]), .B(L[1]), .CI(n_2), .CO(n_3), .S(plus[1]));
   FA_X1 i_4 (.A(R[2]), .B(L[2]), .CI(n_3), .CO(n_4), .S(plus[2]));
   FA_X1 i_5 (.A(R[3]), .B(L[3]), .CI(n_4), .CO(n_5), .S(plus[3]));
   FA_X1 i_6 (.A(R[4]), .B(L[4]), .CI(n_5), .CO(n_6), .S(plus[4]));
   FA_X1 i_7 (.A(R[5]), .B(L[5]), .CI(n_6), .CO(n_7), .S(plus[5]));
   FA_X1 i_8 (.A(R[6]), .B(L[6]), .CI(n_7), .CO(n_8), .S(plus[6]));
   FA_X1 i_9 (.A(R[7]), .B(L[7]), .CI(n_8), .CO(n_9), .S(plus[7]));
   FA_X1 i_10 (.A(R[8]), .B(L[8]), .CI(n_9), .CO(n_10), .S(plus[8]));
   FA_X1 i_11 (.A(R[9]), .B(L[9]), .CI(n_10), .CO(n_11), .S(plus[9]));
   FA_X1 i_12 (.A(R[10]), .B(L[10]), .CI(n_11), .CO(n_12), .S(plus[10]));
   FA_X1 i_13 (.A(R[11]), .B(L[11]), .CI(n_12), .CO(n_13), .S(plus[11]));
   FA_X1 i_14 (.A(R[12]), .B(L[12]), .CI(n_13), .CO(n_14), .S(plus[12]));
   FA_X1 i_15 (.A(R[13]), .B(L[13]), .CI(n_14), .CO(n_15), .S(plus[13]));
   FA_X1 i_16 (.A(R[14]), .B(L[14]), .CI(n_15), .CO(n_16), .S(plus[14]));
   FA_X1 i_17 (.A(L[15]), .B(R[15]), .CI(n_16), .CO(n_17), .S(plus[15]));
   FA_X1 i_18 (.A(n_0), .B(n_1), .CI(n_17), .CO(n_18), .S(plus[16]));
   INV_X1 i_19 (.A(n_18), .ZN(plus[20]));
endmodule

module datapath__0_49(R, L, plus);
   input [19:0]R;
   input [19:0]L;
   output [19:0]plus;

   INV_X1 i_0 (.A(R[15]), .ZN(n_0));
   INV_X1 i_1 (.A(L[19]), .ZN(n_1));
   HA_X1 i_2 (.A(R[0]), .B(L[0]), .CO(n_2), .S(plus[0]));
   FA_X1 i_3 (.A(R[1]), .B(L[1]), .CI(n_2), .CO(n_3), .S(plus[1]));
   FA_X1 i_4 (.A(R[2]), .B(L[2]), .CI(n_3), .CO(n_4), .S(plus[2]));
   FA_X1 i_5 (.A(R[3]), .B(L[3]), .CI(n_4), .CO(n_5), .S(plus[3]));
   FA_X1 i_6 (.A(R[4]), .B(L[4]), .CI(n_5), .CO(n_6), .S(plus[4]));
   FA_X1 i_7 (.A(R[5]), .B(L[5]), .CI(n_6), .CO(n_7), .S(plus[5]));
   FA_X1 i_8 (.A(R[6]), .B(L[6]), .CI(n_7), .CO(n_8), .S(plus[6]));
   FA_X1 i_9 (.A(R[7]), .B(L[7]), .CI(n_8), .CO(n_9), .S(plus[7]));
   FA_X1 i_10 (.A(R[8]), .B(L[8]), .CI(n_9), .CO(n_10), .S(plus[8]));
   FA_X1 i_11 (.A(R[9]), .B(L[9]), .CI(n_10), .CO(n_11), .S(plus[9]));
   FA_X1 i_12 (.A(R[10]), .B(L[10]), .CI(n_11), .CO(n_12), .S(plus[10]));
   FA_X1 i_13 (.A(R[11]), .B(L[11]), .CI(n_12), .CO(n_13), .S(plus[11]));
   FA_X1 i_14 (.A(R[12]), .B(L[12]), .CI(n_13), .CO(n_14), .S(plus[12]));
   FA_X1 i_15 (.A(R[13]), .B(L[13]), .CI(n_14), .CO(n_15), .S(plus[13]));
   FA_X1 i_16 (.A(R[14]), .B(L[14]), .CI(n_15), .CO(n_16), .S(plus[14]));
   FA_X1 i_17 (.A(L[15]), .B(R[15]), .CI(n_16), .CO(n_17), .S(plus[15]));
   FA_X1 i_18 (.A(n_0), .B(n_1), .CI(n_17), .CO(n_18), .S(plus[16]));
   INV_X1 i_19 (.A(n_18), .ZN(plus[19]));
endmodule

module datapath__0_53(R, L, plus);
   input [18:0]R;
   input [18:0]L;
   output [18:0]plus;

   INV_X1 i_0 (.A(R[15]), .ZN(n_0));
   INV_X1 i_1 (.A(L[18]), .ZN(n_1));
   HA_X1 i_2 (.A(R[0]), .B(L[0]), .CO(n_2), .S(plus[0]));
   FA_X1 i_3 (.A(R[1]), .B(L[1]), .CI(n_2), .CO(n_3), .S(plus[1]));
   FA_X1 i_4 (.A(R[2]), .B(L[2]), .CI(n_3), .CO(n_4), .S(plus[2]));
   FA_X1 i_5 (.A(R[3]), .B(L[3]), .CI(n_4), .CO(n_5), .S(plus[3]));
   FA_X1 i_6 (.A(R[4]), .B(L[4]), .CI(n_5), .CO(n_6), .S(plus[4]));
   FA_X1 i_7 (.A(R[5]), .B(L[5]), .CI(n_6), .CO(n_7), .S(plus[5]));
   FA_X1 i_8 (.A(R[6]), .B(L[6]), .CI(n_7), .CO(n_8), .S(plus[6]));
   FA_X1 i_9 (.A(R[7]), .B(L[7]), .CI(n_8), .CO(n_9), .S(plus[7]));
   FA_X1 i_10 (.A(R[8]), .B(L[8]), .CI(n_9), .CO(n_10), .S(plus[8]));
   FA_X1 i_11 (.A(R[9]), .B(L[9]), .CI(n_10), .CO(n_11), .S(plus[9]));
   FA_X1 i_12 (.A(R[10]), .B(L[10]), .CI(n_11), .CO(n_12), .S(plus[10]));
   FA_X1 i_13 (.A(R[11]), .B(L[11]), .CI(n_12), .CO(n_13), .S(plus[11]));
   FA_X1 i_14 (.A(R[12]), .B(L[12]), .CI(n_13), .CO(n_14), .S(plus[12]));
   FA_X1 i_15 (.A(R[13]), .B(L[13]), .CI(n_14), .CO(n_15), .S(plus[13]));
   FA_X1 i_16 (.A(R[14]), .B(L[14]), .CI(n_15), .CO(n_16), .S(plus[14]));
   FA_X1 i_17 (.A(L[15]), .B(R[15]), .CI(n_16), .CO(n_17), .S(plus[15]));
   FA_X1 i_18 (.A(n_0), .B(n_1), .CI(n_17), .CO(n_18), .S(plus[16]));
   INV_X1 i_19 (.A(n_18), .ZN(plus[18]));
endmodule

module datapath__0_57(R, L, plus);
   input [17:0]R;
   input [17:0]L;
   output [17:0]plus;

   INV_X1 i_0 (.A(R[15]), .ZN(n_0));
   INV_X1 i_1 (.A(L[17]), .ZN(n_1));
   HA_X1 i_2 (.A(R[0]), .B(L[0]), .CO(n_2), .S(plus[0]));
   FA_X1 i_3 (.A(R[1]), .B(L[1]), .CI(n_2), .CO(n_3), .S(plus[1]));
   FA_X1 i_4 (.A(R[2]), .B(L[2]), .CI(n_3), .CO(n_4), .S(plus[2]));
   FA_X1 i_5 (.A(R[3]), .B(L[3]), .CI(n_4), .CO(n_5), .S(plus[3]));
   FA_X1 i_6 (.A(R[4]), .B(L[4]), .CI(n_5), .CO(n_6), .S(plus[4]));
   FA_X1 i_7 (.A(R[5]), .B(L[5]), .CI(n_6), .CO(n_7), .S(plus[5]));
   FA_X1 i_8 (.A(R[6]), .B(L[6]), .CI(n_7), .CO(n_8), .S(plus[6]));
   FA_X1 i_9 (.A(R[7]), .B(L[7]), .CI(n_8), .CO(n_9), .S(plus[7]));
   FA_X1 i_10 (.A(R[8]), .B(L[8]), .CI(n_9), .CO(n_10), .S(plus[8]));
   FA_X1 i_11 (.A(R[9]), .B(L[9]), .CI(n_10), .CO(n_11), .S(plus[9]));
   FA_X1 i_12 (.A(R[10]), .B(L[10]), .CI(n_11), .CO(n_12), .S(plus[10]));
   FA_X1 i_13 (.A(R[11]), .B(L[11]), .CI(n_12), .CO(n_13), .S(plus[11]));
   FA_X1 i_14 (.A(R[12]), .B(L[12]), .CI(n_13), .CO(n_14), .S(plus[12]));
   FA_X1 i_15 (.A(R[13]), .B(L[13]), .CI(n_14), .CO(n_15), .S(plus[13]));
   FA_X1 i_16 (.A(R[14]), .B(L[14]), .CI(n_15), .CO(n_16), .S(plus[14]));
   FA_X1 i_17 (.A(L[15]), .B(R[15]), .CI(n_16), .CO(n_17), .S(plus[15]));
   FA_X1 i_18 (.A(n_0), .B(n_1), .CI(n_17), .CO(n_18), .S(plus[16]));
   INV_X1 i_19 (.A(n_18), .ZN(plus[17]));
endmodule

module datapath__0_60(L, plus, p_0);
   input [16:0]L;
   output [16:0]plus;
   input [16:0]p_0;

   FA_X1 i_117 (.A(p_0[15]), .B(n_2), .CI(n_1), .CO(n_0), .S(plus[15]));
   XNOR2_X1 i_0 (.A(L[1]), .B(p_0[1]), .ZN(n_3));
   INV_X1 i_1 (.A(L[0]), .ZN(n_4));
   NAND2_X1 i_2 (.A1(n_4), .A2(p_0[0]), .ZN(n_5));
   INV_X1 i_3 (.A(n_5), .ZN(n_6));
   INV_X1 i_4 (.A(L[1]), .ZN(n_7));
   AOI22_X1 i_5 (.A1(n_3), .A2(n_6), .B1(n_7), .B2(p_0[1]), .ZN(n_8));
   XOR2_X1 i_6 (.A(p_0[2]), .B(L[2]), .Z(n_9));
   INV_X1 i_7 (.A(p_0[2]), .ZN(n_10));
   OAI22_X1 i_8 (.A1(n_8), .A2(n_9), .B1(n_10), .B2(L[2]), .ZN(n_11));
   XNOR2_X1 i_9 (.A(L[3]), .B(p_0[3]), .ZN(n_12));
   INV_X1 i_10 (.A(L[3]), .ZN(n_13));
   AOI22_X1 i_11 (.A1(n_11), .A2(n_12), .B1(n_13), .B2(p_0[3]), .ZN(n_14));
   XOR2_X1 i_12 (.A(p_0[4]), .B(L[4]), .Z(n_15));
   INV_X1 i_13 (.A(p_0[4]), .ZN(n_16));
   OAI22_X1 i_14 (.A1(n_14), .A2(n_15), .B1(n_16), .B2(L[4]), .ZN(n_17));
   XNOR2_X1 i_15 (.A(L[5]), .B(p_0[5]), .ZN(n_18));
   INV_X1 i_16 (.A(L[5]), .ZN(n_19));
   AOI22_X1 i_17 (.A1(n_17), .A2(n_18), .B1(n_19), .B2(p_0[5]), .ZN(n_20));
   XOR2_X1 i_18 (.A(p_0[6]), .B(L[6]), .Z(n_21));
   INV_X1 i_19 (.A(p_0[6]), .ZN(n_22));
   OAI22_X1 i_20 (.A1(n_20), .A2(n_21), .B1(n_22), .B2(L[6]), .ZN(n_23));
   XNOR2_X1 i_21 (.A(L[7]), .B(p_0[7]), .ZN(n_24));
   INV_X1 i_22 (.A(L[7]), .ZN(n_25));
   AOI22_X1 i_23 (.A1(n_23), .A2(n_24), .B1(n_25), .B2(p_0[7]), .ZN(n_26));
   XOR2_X1 i_24 (.A(p_0[8]), .B(L[8]), .Z(n_27));
   INV_X1 i_25 (.A(p_0[8]), .ZN(n_28));
   OAI22_X1 i_26 (.A1(n_26), .A2(n_27), .B1(n_28), .B2(L[8]), .ZN(n_29));
   XNOR2_X1 i_27 (.A(L[9]), .B(p_0[9]), .ZN(n_30));
   INV_X1 i_28 (.A(L[9]), .ZN(n_31));
   AOI22_X1 i_29 (.A1(n_29), .A2(n_30), .B1(n_31), .B2(p_0[9]), .ZN(n_32));
   XOR2_X1 i_30 (.A(p_0[10]), .B(L[10]), .Z(n_33));
   INV_X1 i_31 (.A(p_0[10]), .ZN(n_34));
   OAI22_X1 i_32 (.A1(n_32), .A2(n_33), .B1(n_34), .B2(L[10]), .ZN(n_35));
   XNOR2_X1 i_33 (.A(L[11]), .B(p_0[11]), .ZN(n_36));
   INV_X1 i_34 (.A(L[11]), .ZN(n_37));
   AOI22_X1 i_35 (.A1(n_35), .A2(n_36), .B1(n_37), .B2(p_0[11]), .ZN(n_38));
   XOR2_X1 i_36 (.A(p_0[12]), .B(L[12]), .Z(n_39));
   INV_X1 i_37 (.A(p_0[12]), .ZN(n_40));
   OAI22_X1 i_38 (.A1(n_38), .A2(n_39), .B1(n_40), .B2(L[12]), .ZN(n_41));
   XNOR2_X1 i_39 (.A(L[13]), .B(p_0[13]), .ZN(n_42));
   INV_X1 i_40 (.A(L[13]), .ZN(n_43));
   AOI22_X1 i_41 (.A1(n_41), .A2(n_42), .B1(n_43), .B2(p_0[13]), .ZN(n_44));
   INV_X1 i_42 (.A(n_44), .ZN(n_45));
   XNOR2_X1 i_43 (.A(L[14]), .B(p_0[14]), .ZN(n_46));
   INV_X1 i_44 (.A(L[14]), .ZN(n_47));
   AOI22_X1 i_45 (.A1(n_45), .A2(n_46), .B1(n_47), .B2(p_0[14]), .ZN(n_1));
   OAI21_X1 i_46 (.A(n_5), .B1(p_0[0]), .B2(n_4), .ZN(plus[0]));
   XOR2_X1 i_47 (.A(n_3), .B(n_5), .Z(plus[1]));
   XNOR2_X1 i_48 (.A(n_8), .B(n_9), .ZN(plus[2]));
   XNOR2_X1 i_49 (.A(n_11), .B(n_12), .ZN(plus[3]));
   XNOR2_X1 i_50 (.A(n_14), .B(n_15), .ZN(plus[4]));
   XNOR2_X1 i_51 (.A(n_17), .B(n_18), .ZN(plus[5]));
   XNOR2_X1 i_52 (.A(n_20), .B(n_21), .ZN(plus[6]));
   XNOR2_X1 i_53 (.A(n_23), .B(n_24), .ZN(plus[7]));
   XNOR2_X1 i_54 (.A(n_26), .B(n_27), .ZN(plus[8]));
   XNOR2_X1 i_55 (.A(n_29), .B(n_30), .ZN(plus[9]));
   XNOR2_X1 i_56 (.A(n_32), .B(n_33), .ZN(plus[10]));
   XNOR2_X1 i_57 (.A(n_35), .B(n_36), .ZN(plus[11]));
   XNOR2_X1 i_58 (.A(n_38), .B(n_39), .ZN(plus[12]));
   XNOR2_X1 i_59 (.A(n_41), .B(n_42), .ZN(plus[13]));
   XOR2_X1 i_60 (.A(n_46), .B(n_44), .Z(plus[14]));
   XNOR2_X1 i_61 (.A(n_0), .B(L[15]), .ZN(n_48));
   XOR2_X1 i_62 (.A(n_48), .B(L[16]), .Z(plus[16]));
   INV_X1 i_63 (.A(L[15]), .ZN(n_2));
endmodule

module fpu_multiplier(mode, clk, rst, enbl, in_a, in_b, out_c, done, err, zero, 
      posv);
   input [1:0]mode;
   input clk;
   input rst;
   input enbl;
   input [63:0]in_a;
   input [63:0]in_b;
   output [63:0]out_c;
   output done;
   output err;
   output zero;
   output posv;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_166;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_180;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_190;
   wire n_0_191;
   wire n_0_192;
   wire n_0_193;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_200;
   wire n_0_201;
   wire n_0_202;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_207;
   wire n_0_208;
   wire n_0_209;
   wire n_0_210;
   wire n_0_211;
   wire n_0_212;
   wire n_0_213;
   wire n_0_214;
   wire n_0_215;
   wire n_0_216;
   wire n_0_217;
   wire n_0_218;
   wire n_0_219;
   wire n_0_220;
   wire n_0_221;
   wire n_0_222;
   wire n_0_223;
   wire n_0_224;
   wire n_0_225;
   wire n_0_226;
   wire n_0_227;
   wire n_0_228;
   wire n_0_229;
   wire n_0_230;
   wire n_0_231;
   wire n_0_232;
   wire n_0_233;
   wire n_0_234;
   wire n_0_235;
   wire n_0_236;
   wire n_0_237;
   wire n_0_238;
   wire n_0_239;
   wire n_0_240;
   wire n_0_241;
   wire n_0_242;
   wire n_0_243;
   wire n_0_244;
   wire n_0_245;
   wire n_0_246;
   wire n_0_247;
   wire n_0_248;
   wire n_0_249;
   wire n_0_250;
   wire n_0_251;
   wire n_0_252;
   wire n_0_253;
   wire n_0_254;
   wire n_0_255;
   wire n_0_256;
   wire n_0_257;
   wire n_0_258;
   wire n_0_259;
   wire n_0_260;
   wire n_0_261;
   wire n_0_262;
   wire error;
   wire n_0_263;
   wire n_0_264;
   wire n_0_4;
   wire n_0_265;
   wire n_0_268;
   wire n_0_267;
   wire n_0_270;
   wire n_0_266;
   wire n_0_1_0;
   wire n_0_269;
   wire n_0_510;
   wire n_0_511;
   wire n_0_512;
   wire n_0_513;
   wire n_0_514;
   wire n_0_515;
   wire n_0_516;
   wire n_0_517;
   wire n_0_518;
   wire n_0_519;
   wire n_0_520;
   wire n_0_521;
   wire n_0_522;
   wire n_0_523;
   wire n_0_524;
   wire n_0_2_0;
   wire n_0_2_1;
   wire n_0_494;
   wire n_0_2_2;
   wire n_0_495;
   wire n_0_2_3;
   wire n_0_496;
   wire n_0_2_4;
   wire n_0_497;
   wire n_0_2_5;
   wire n_0_498;
   wire n_0_2_6;
   wire n_0_499;
   wire n_0_2_7;
   wire n_0_500;
   wire n_0_2_8;
   wire n_0_501;
   wire n_0_2_9;
   wire n_0_502;
   wire n_0_2_10;
   wire n_0_503;
   wire n_0_2_11;
   wire n_0_504;
   wire n_0_2_12;
   wire n_0_505;
   wire n_0_2_13;
   wire n_0_506;
   wire n_0_2_14;
   wire n_0_2_15;
   wire n_0_507;
   wire n_0_2_16;
   wire n_0_508;
   wire n_0_2_17;
   wire n_0_509;
   wire n_0_2_18;
   wire n_0_2_19;
   wire n_0_477;
   wire n_0_2_20;
   wire n_0_478;
   wire n_0_2_21;
   wire n_0_479;
   wire n_0_2_22;
   wire n_0_480;
   wire n_0_2_23;
   wire n_0_481;
   wire n_0_2_24;
   wire n_0_482;
   wire n_0_2_25;
   wire n_0_483;
   wire n_0_2_26;
   wire n_0_484;
   wire n_0_2_27;
   wire n_0_485;
   wire n_0_2_28;
   wire n_0_486;
   wire n_0_2_29;
   wire n_0_487;
   wire n_0_2_30;
   wire n_0_488;
   wire n_0_2_31;
   wire n_0_489;
   wire n_0_2_32;
   wire n_0_490;
   wire n_0_2_33;
   wire n_0_491;
   wire n_0_2_34;
   wire n_0_492;
   wire n_0_2_35;
   wire n_0_493;
   wire n_0_460;
   wire n_0_461;
   wire n_0_462;
   wire n_0_463;
   wire n_0_464;
   wire n_0_465;
   wire n_0_466;
   wire n_0_467;
   wire n_0_468;
   wire n_0_469;
   wire n_0_470;
   wire n_0_471;
   wire n_0_472;
   wire n_0_473;
   wire n_0_474;
   wire n_0_475;
   wire n_0_476;
   wire n_0_443;
   wire n_0_444;
   wire n_0_445;
   wire n_0_446;
   wire n_0_447;
   wire n_0_448;
   wire n_0_449;
   wire n_0_450;
   wire n_0_451;
   wire n_0_452;
   wire n_0_453;
   wire n_0_454;
   wire n_0_455;
   wire n_0_456;
   wire n_0_457;
   wire n_0_458;
   wire n_0_459;
   wire n_0_426;
   wire n_0_427;
   wire n_0_428;
   wire n_0_429;
   wire n_0_430;
   wire n_0_431;
   wire n_0_432;
   wire n_0_433;
   wire n_0_434;
   wire n_0_435;
   wire n_0_436;
   wire n_0_437;
   wire n_0_438;
   wire n_0_439;
   wire n_0_440;
   wire n_0_441;
   wire n_0_442;
   wire n_0_409;
   wire n_0_410;
   wire n_0_411;
   wire n_0_412;
   wire n_0_413;
   wire n_0_414;
   wire n_0_415;
   wire n_0_416;
   wire n_0_417;
   wire n_0_418;
   wire n_0_419;
   wire n_0_420;
   wire n_0_421;
   wire n_0_422;
   wire n_0_423;
   wire n_0_424;
   wire n_0_425;
   wire n_0_391;
   wire n_0_392;
   wire n_0_393;
   wire n_0_394;
   wire n_0_395;
   wire n_0_396;
   wire n_0_397;
   wire n_0_398;
   wire n_0_399;
   wire n_0_400;
   wire n_0_401;
   wire n_0_402;
   wire n_0_403;
   wire n_0_404;
   wire n_0_405;
   wire n_0_406;
   wire n_0_407;
   wire n_0_408;
   wire n_0_373;
   wire n_0_374;
   wire n_0_375;
   wire n_0_376;
   wire n_0_377;
   wire n_0_378;
   wire n_0_379;
   wire n_0_380;
   wire n_0_381;
   wire n_0_382;
   wire n_0_383;
   wire n_0_384;
   wire n_0_385;
   wire n_0_386;
   wire n_0_387;
   wire n_0_388;
   wire n_0_389;
   wire n_0_390;
   wire n_0_355;
   wire n_0_356;
   wire n_0_357;
   wire n_0_358;
   wire n_0_359;
   wire n_0_360;
   wire n_0_361;
   wire n_0_362;
   wire n_0_363;
   wire n_0_364;
   wire n_0_365;
   wire n_0_366;
   wire n_0_367;
   wire n_0_368;
   wire n_0_369;
   wire n_0_370;
   wire n_0_371;
   wire n_0_372;
   wire n_0_337;
   wire n_0_338;
   wire n_0_339;
   wire n_0_340;
   wire n_0_341;
   wire n_0_342;
   wire n_0_343;
   wire n_0_344;
   wire n_0_345;
   wire n_0_346;
   wire n_0_347;
   wire n_0_348;
   wire n_0_349;
   wire n_0_350;
   wire n_0_351;
   wire n_0_352;
   wire n_0_353;
   wire n_0_354;
   wire n_0_319;
   wire n_0_320;
   wire n_0_321;
   wire n_0_322;
   wire n_0_323;
   wire n_0_324;
   wire n_0_325;
   wire n_0_326;
   wire n_0_327;
   wire n_0_328;
   wire n_0_329;
   wire n_0_330;
   wire n_0_331;
   wire n_0_332;
   wire n_0_333;
   wire n_0_334;
   wire n_0_335;
   wire n_0_336;
   wire n_0_301;
   wire n_0_302;
   wire n_0_303;
   wire n_0_304;
   wire n_0_305;
   wire n_0_306;
   wire n_0_307;
   wire n_0_308;
   wire n_0_309;
   wire n_0_310;
   wire n_0_311;
   wire n_0_312;
   wire n_0_313;
   wire n_0_314;
   wire n_0_315;
   wire n_0_316;
   wire n_0_317;
   wire n_0_318;
   wire n_0_283;
   wire n_0_284;
   wire n_0_285;
   wire n_0_286;
   wire n_0_287;
   wire n_0_288;
   wire n_0_289;
   wire n_0_290;
   wire n_0_291;
   wire n_0_292;
   wire n_0_293;
   wire n_0_294;
   wire n_0_295;
   wire n_0_296;
   wire n_0_297;
   wire n_0_298;
   wire n_0_299;
   wire n_0_300;
   wire [31:0]\output ;
   wire n_0_274;
   wire n_0_275;
   wire n_0_276;
   wire n_0_277;
   wire n_0_278;
   wire n_0_279;
   wire n_0_280;
   wire n_0_281;
   wire n_0_2_46;
   wire n_0_2_47;
   wire n_0_2_48;
   wire n_0_2_49;
   wire n_0_2_50;
   wire n_0_2_51;
   wire n_0_2_52;
   wire n_0_2_53;
   wire n_0_282;
   wire n_0_2_36;
   wire n_0_2_37;
   wire n_0_2_38;
   wire n_0_2_39;
   wire n_0_273;
   wire n_0_272;
   wire n_0_2_40;
   wire n_0_2_41;
   wire n_0_2_42;
   wire n_0_2_43;
   wire n_0_2_44;
   wire n_0_2_45;
   wire n_0_271;

   assign out_c[63] = out_c[16];
   assign out_c[62] = out_c[16];
   assign out_c[61] = out_c[16];
   assign out_c[60] = out_c[16];
   assign out_c[59] = out_c[16];
   assign out_c[58] = out_c[16];
   assign out_c[57] = out_c[16];
   assign out_c[56] = out_c[16];
   assign out_c[55] = out_c[16];
   assign out_c[54] = out_c[16];
   assign out_c[53] = out_c[16];
   assign out_c[52] = out_c[16];
   assign out_c[51] = out_c[16];
   assign out_c[50] = out_c[16];
   assign out_c[49] = out_c[16];
   assign out_c[48] = out_c[16];
   assign out_c[47] = out_c[16];
   assign out_c[46] = out_c[16];
   assign out_c[45] = out_c[16];
   assign out_c[44] = out_c[16];
   assign out_c[43] = out_c[16];
   assign out_c[42] = out_c[16];
   assign out_c[41] = out_c[16];
   assign out_c[40] = out_c[16];
   assign out_c[39] = out_c[16];
   assign out_c[38] = out_c[16];
   assign out_c[37] = out_c[16];
   assign out_c[36] = out_c[16];
   assign out_c[35] = out_c[16];
   assign out_c[34] = out_c[16];
   assign out_c[33] = out_c[16];
   assign out_c[32] = out_c[16];
   assign out_c[31] = out_c[16];
   assign out_c[30] = out_c[16];
   assign out_c[29] = out_c[16];
   assign out_c[28] = out_c[16];
   assign out_c[27] = out_c[16];
   assign out_c[26] = out_c[16];
   assign out_c[25] = out_c[16];
   assign out_c[24] = out_c[16];
   assign out_c[23] = out_c[16];
   assign out_c[22] = out_c[16];
   assign out_c[21] = out_c[16];
   assign out_c[20] = out_c[16];
   assign out_c[19] = out_c[16];
   assign out_c[18] = out_c[16];
   assign out_c[17] = out_c[16];

   DFFR_X1 posv_reg (.D(n_0_272), .RN(n_0_267), .CK(n_0_4), .Q(posv), .QN());
   datapath i_0_5 (.R({uc_0, uc_1, uc_2, uc_3, uc_4, uc_5, uc_6, uc_7, uc_8, 
      uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, in_a[15], in_a[14], in_a[13], 
      in_a[12], in_a[11], in_a[10], in_a[9], in_a[8], in_a[7], in_a[6], in_a[5], 
      in_a[4], in_a[3], in_a[2], in_a[1], in_a[0]}), .L({uc_15, uc_16, uc_17, 
      uc_18, uc_19, uc_20, uc_21, uc_22, uc_23, uc_24, uc_25, uc_26, uc_27, 
      uc_28, uc_29, uc_30, n_0_524, n_0_523, n_0_522, n_0_521, n_0_520, n_0_519, 
      n_0_518, n_0_517, n_0_516, n_0_515, n_0_514, n_0_513, n_0_512, n_0_511, 
      n_0_510}), .plus({n_0_16, uc_31, uc_32, uc_33, uc_34, uc_35, uc_36, uc_37, 
      uc_38, uc_39, uc_40, uc_41, uc_42, uc_43, uc_44, n_0_15, n_0_14, n_0_13, 
      n_0_12, n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_3, n_0_2, 
      n_0_1, n_0_0, uc_45}));
   datapath__0_9 i_0_7 (.R({uc_46, uc_47, uc_48, uc_49, uc_50, uc_51, uc_52, 
      uc_53, uc_54, uc_55, uc_56, uc_57, uc_58, uc_59, in_a[15], in_a[14], 
      in_a[13], in_a[12], in_a[11], in_a[10], in_a[9], in_a[8], in_a[7], in_a[6], 
      in_a[5], in_a[4], in_a[3], in_a[2], in_a[1], in_a[0]}), .L({n_0_509, uc_60, 
      uc_61, uc_62, uc_63, uc_64, uc_65, uc_66, uc_67, uc_68, uc_69, uc_70, 
      uc_71, uc_72, uc_73, n_0_508, n_0_507, n_0_506, n_0_505, n_0_504, n_0_503, 
      n_0_502, n_0_501, n_0_500, n_0_499, n_0_498, n_0_497, n_0_496, n_0_495, 
      n_0_494}), .plus({n_0_33, uc_74, uc_75, uc_76, uc_77, uc_78, uc_79, uc_80, 
      uc_81, uc_82, uc_83, uc_84, uc_85, n_0_32, n_0_31, n_0_30, n_0_29, n_0_28, 
      n_0_27, n_0_26, n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, 
      n_0_18, n_0_17, uc_86}));
   datapath__0_13 i_0_9 (.R({uc_87, uc_88, uc_89, uc_90, uc_91, uc_92, uc_93, 
      uc_94, uc_95, uc_96, uc_97, uc_98, uc_99, in_a[15], in_a[14], in_a[13], 
      in_a[12], in_a[11], in_a[10], in_a[9], in_a[8], in_a[7], in_a[6], in_a[5], 
      in_a[4], in_a[3], in_a[2], in_a[1], in_a[0]}), .L({n_0_493, uc_100, uc_101, 
      uc_102, uc_103, uc_104, uc_105, uc_106, uc_107, uc_108, uc_109, uc_110, 
      uc_111, n_0_492, n_0_491, n_0_490, n_0_489, n_0_488, n_0_487, n_0_486, 
      n_0_485, n_0_484, n_0_483, n_0_482, n_0_481, n_0_480, n_0_479, n_0_478, 
      n_0_477}), .plus({n_0_50, uc_112, uc_113, uc_114, uc_115, uc_116, uc_117, 
      uc_118, uc_119, uc_120, uc_121, uc_122, n_0_49, n_0_48, n_0_47, n_0_46, 
      n_0_45, n_0_44, n_0_43, n_0_42, n_0_41, n_0_40, n_0_39, n_0_38, n_0_37, 
      n_0_36, n_0_35, n_0_34, uc_123}));
   datapath__0_17 i_0_11 (.R({uc_124, uc_125, uc_126, uc_127, uc_128, uc_129, 
      uc_130, uc_131, uc_132, uc_133, uc_134, uc_135, in_a[15], in_a[14], 
      in_a[13], in_a[12], in_a[11], in_a[10], in_a[9], in_a[8], in_a[7], in_a[6], 
      in_a[5], in_a[4], in_a[3], in_a[2], in_a[1], in_a[0]}), .L({n_0_476, 
      uc_136, uc_137, uc_138, uc_139, uc_140, uc_141, uc_142, uc_143, uc_144, 
      uc_145, uc_146, n_0_475, n_0_474, n_0_473, n_0_472, n_0_471, n_0_470, 
      n_0_469, n_0_468, n_0_467, n_0_466, n_0_465, n_0_464, n_0_463, n_0_462, 
      n_0_461, n_0_460}), .plus({n_0_67, uc_147, uc_148, uc_149, uc_150, uc_151, 
      uc_152, uc_153, uc_154, uc_155, uc_156, n_0_66, n_0_65, n_0_64, n_0_63, 
      n_0_62, n_0_61, n_0_60, n_0_59, n_0_58, n_0_57, n_0_56, n_0_55, n_0_54, 
      n_0_53, n_0_52, n_0_51, uc_157}));
   datapath__0_21 i_0_13 (.R({uc_158, uc_159, uc_160, uc_161, uc_162, uc_163, 
      uc_164, uc_165, uc_166, uc_167, uc_168, in_a[15], in_a[14], in_a[13], 
      in_a[12], in_a[11], in_a[10], in_a[9], in_a[8], in_a[7], in_a[6], in_a[5], 
      in_a[4], in_a[3], in_a[2], in_a[1], in_a[0]}), .L({n_0_459, uc_169, uc_170, 
      uc_171, uc_172, uc_173, uc_174, uc_175, uc_176, uc_177, uc_178, n_0_458, 
      n_0_457, n_0_456, n_0_455, n_0_454, n_0_453, n_0_452, n_0_451, n_0_450, 
      n_0_449, n_0_448, n_0_447, n_0_446, n_0_445, n_0_444, n_0_443}), .plus({
      n_0_84, uc_179, uc_180, uc_181, uc_182, uc_183, uc_184, uc_185, uc_186, 
      uc_187, n_0_83, n_0_82, n_0_81, n_0_80, n_0_79, n_0_78, n_0_77, n_0_76, 
      n_0_75, n_0_74, n_0_73, n_0_72, n_0_71, n_0_70, n_0_69, n_0_68, uc_188}));
   datapath__0_25 i_0_15 (.R({uc_189, uc_190, uc_191, uc_192, uc_193, uc_194, 
      uc_195, uc_196, uc_197, uc_198, in_a[15], in_a[14], in_a[13], in_a[12], 
      in_a[11], in_a[10], in_a[9], in_a[8], in_a[7], in_a[6], in_a[5], in_a[4], 
      in_a[3], in_a[2], in_a[1], in_a[0]}), .L({n_0_442, uc_199, uc_200, uc_201, 
      uc_202, uc_203, uc_204, uc_205, uc_206, uc_207, n_0_441, n_0_440, n_0_439, 
      n_0_438, n_0_437, n_0_436, n_0_435, n_0_434, n_0_433, n_0_432, n_0_431, 
      n_0_430, n_0_429, n_0_428, n_0_427, n_0_426}), .plus({n_0_101, uc_208, 
      uc_209, uc_210, uc_211, uc_212, uc_213, uc_214, uc_215, n_0_100, n_0_99, 
      n_0_98, n_0_97, n_0_96, n_0_95, n_0_94, n_0_93, n_0_92, n_0_91, n_0_90, 
      n_0_89, n_0_88, n_0_87, n_0_86, n_0_85, uc_216}));
   datapath__0_29 i_0_17 (.R({uc_217, uc_218, uc_219, uc_220, uc_221, uc_222, 
      uc_223, uc_224, uc_225, in_a[15], in_a[14], in_a[13], in_a[12], in_a[11], 
      in_a[10], in_a[9], in_a[8], in_a[7], in_a[6], in_a[5], in_a[4], in_a[3], 
      in_a[2], in_a[1], in_a[0]}), .L({n_0_425, uc_226, uc_227, uc_228, uc_229, 
      uc_230, uc_231, uc_232, uc_233, n_0_424, n_0_423, n_0_422, n_0_421, 
      n_0_420, n_0_419, n_0_418, n_0_417, n_0_416, n_0_415, n_0_414, n_0_413, 
      n_0_412, n_0_411, n_0_410, n_0_409}), .plus({n_0_119, uc_234, uc_235, 
      uc_236, uc_237, uc_238, uc_239, uc_240, n_0_118, n_0_117, n_0_116, n_0_115, 
      n_0_114, n_0_113, n_0_112, n_0_111, n_0_110, n_0_109, n_0_108, n_0_107, 
      n_0_106, n_0_105, n_0_104, n_0_103, n_0_102}));
   datapath__0_33 i_0_19 (.R({uc_241, uc_242, uc_243, uc_244, uc_245, uc_246, 
      uc_247, uc_248, in_a[15], in_a[14], in_a[13], in_a[12], in_a[11], in_a[10], 
      in_a[9], in_a[8], in_a[7], in_a[6], in_a[5], in_a[4], in_a[3], in_a[2], 
      in_a[1], in_a[0]}), .L({n_0_408, uc_249, uc_250, uc_251, uc_252, uc_253, 
      uc_254, uc_255, n_0_407, n_0_406, n_0_405, n_0_404, n_0_403, n_0_402, 
      n_0_401, n_0_400, n_0_399, n_0_398, n_0_397, n_0_396, n_0_395, n_0_394, 
      n_0_393, n_0_392}), .plus({n_0_137, uc_256, uc_257, uc_258, uc_259, uc_260, 
      uc_261, n_0_136, n_0_135, n_0_134, n_0_133, n_0_132, n_0_131, n_0_130, 
      n_0_129, n_0_128, n_0_127, n_0_126, n_0_125, n_0_124, n_0_123, n_0_122, 
      n_0_121, n_0_120}));
   datapath__0_37 i_0_21 (.R({uc_262, uc_263, uc_264, uc_265, uc_266, uc_267, 
      uc_268, in_a[15], in_a[14], in_a[13], in_a[12], in_a[11], in_a[10], 
      in_a[9], in_a[8], in_a[7], in_a[6], in_a[5], in_a[4], in_a[3], in_a[2], 
      in_a[1], in_a[0]}), .L({n_0_390, uc_269, uc_270, uc_271, uc_272, uc_273, 
      uc_274, n_0_389, n_0_388, n_0_387, n_0_386, n_0_385, n_0_384, n_0_383, 
      n_0_382, n_0_381, n_0_380, n_0_379, n_0_378, n_0_377, n_0_376, n_0_375, 
      n_0_374}), .plus({n_0_155, uc_275, uc_276, uc_277, uc_278, uc_279, n_0_154, 
      n_0_153, n_0_152, n_0_151, n_0_150, n_0_149, n_0_148, n_0_147, n_0_146, 
      n_0_145, n_0_144, n_0_143, n_0_142, n_0_141, n_0_140, n_0_139, n_0_138}));
   datapath__0_41 i_0_23 (.R({uc_280, uc_281, uc_282, uc_283, uc_284, uc_285, 
      in_a[15], in_a[14], in_a[13], in_a[12], in_a[11], in_a[10], in_a[9], 
      in_a[8], in_a[7], in_a[6], in_a[5], in_a[4], in_a[3], in_a[2], in_a[1], 
      in_a[0]}), .L({n_0_372, uc_286, uc_287, uc_288, uc_289, uc_290, n_0_371, 
      n_0_370, n_0_369, n_0_368, n_0_367, n_0_366, n_0_365, n_0_364, n_0_363, 
      n_0_362, n_0_361, n_0_360, n_0_359, n_0_358, n_0_357, n_0_356}), .plus({
      n_0_173, uc_291, uc_292, uc_293, uc_294, n_0_172, n_0_171, n_0_170, 
      n_0_169, n_0_168, n_0_167, n_0_166, n_0_165, n_0_164, n_0_163, n_0_162, 
      n_0_161, n_0_160, n_0_159, n_0_158, n_0_157, n_0_156}));
   datapath__0_45 i_0_25 (.R({uc_295, uc_296, uc_297, uc_298, uc_299, in_a[15], 
      in_a[14], in_a[13], in_a[12], in_a[11], in_a[10], in_a[9], in_a[8], 
      in_a[7], in_a[6], in_a[5], in_a[4], in_a[3], in_a[2], in_a[1], in_a[0]}), 
      .L({n_0_354, uc_300, uc_301, uc_302, uc_303, n_0_353, n_0_352, n_0_351, 
      n_0_350, n_0_349, n_0_348, n_0_347, n_0_346, n_0_345, n_0_344, n_0_343, 
      n_0_342, n_0_341, n_0_340, n_0_339, n_0_338}), .plus({n_0_191, uc_304, 
      uc_305, uc_306, n_0_190, n_0_189, n_0_188, n_0_187, n_0_186, n_0_185, 
      n_0_184, n_0_183, n_0_182, n_0_181, n_0_180, n_0_179, n_0_178, n_0_177, 
      n_0_176, n_0_175, n_0_174}));
   datapath__0_49 i_0_27 (.R({uc_307, uc_308, uc_309, uc_310, in_a[15], in_a[14], 
      in_a[13], in_a[12], in_a[11], in_a[10], in_a[9], in_a[8], in_a[7], in_a[6], 
      in_a[5], in_a[4], in_a[3], in_a[2], in_a[1], in_a[0]}), .L({n_0_336, 
      uc_311, uc_312, uc_313, n_0_335, n_0_334, n_0_333, n_0_332, n_0_331, 
      n_0_330, n_0_329, n_0_328, n_0_327, n_0_326, n_0_325, n_0_324, n_0_323, 
      n_0_322, n_0_321, n_0_320}), .plus({n_0_209, uc_314, uc_315, n_0_208, 
      n_0_207, n_0_206, n_0_205, n_0_204, n_0_203, n_0_202, n_0_201, n_0_200, 
      n_0_199, n_0_198, n_0_197, n_0_196, n_0_195, n_0_194, n_0_193, n_0_192}));
   datapath__0_53 i_0_29 (.R({uc_316, uc_317, uc_318, in_a[15], in_a[14], 
      in_a[13], in_a[12], in_a[11], in_a[10], in_a[9], in_a[8], in_a[7], in_a[6], 
      in_a[5], in_a[4], in_a[3], in_a[2], in_a[1], in_a[0]}), .L({n_0_318, 
      uc_319, uc_320, n_0_317, n_0_316, n_0_315, n_0_314, n_0_313, n_0_312, 
      n_0_311, n_0_310, n_0_309, n_0_308, n_0_307, n_0_306, n_0_305, n_0_304, 
      n_0_303, n_0_302}), .plus({n_0_227, uc_321, n_0_226, n_0_225, n_0_224, 
      n_0_223, n_0_222, n_0_221, n_0_220, n_0_219, n_0_218, n_0_217, n_0_216, 
      n_0_215, n_0_214, n_0_213, n_0_212, n_0_211, n_0_210}));
   datapath__0_57 i_0_31 (.R({uc_322, uc_323, in_a[15], in_a[14], in_a[13], 
      in_a[12], in_a[11], in_a[10], in_a[9], in_a[8], in_a[7], in_a[6], in_a[5], 
      in_a[4], in_a[3], in_a[2], in_a[1], in_a[0]}), .L({n_0_300, uc_324, 
      n_0_299, n_0_298, n_0_297, n_0_296, n_0_295, n_0_294, n_0_293, n_0_292, 
      n_0_291, n_0_290, n_0_289, n_0_288, n_0_287, n_0_286, n_0_285, n_0_284}), 
      .plus({n_0_245, n_0_244, n_0_243, n_0_242, n_0_241, n_0_240, n_0_239, 
      n_0_238, n_0_237, n_0_236, n_0_235, n_0_234, n_0_233, n_0_232, n_0_231, 
      n_0_230, n_0_229, n_0_228}));
   datapath__0_60 i_0_33 (.L({\output [31], \output [30], \output [29], 
      \output [28], \output [27], \output [26], \output [25], \output [24], 
      \output [23], \output [22], \output [21], \output [20], \output [19], 
      \output [18], \output [17], \output [16], \output [15]}), .plus({n_0_262, 
      n_0_261, n_0_260, n_0_259, n_0_258, n_0_257, n_0_256, n_0_255, n_0_254, 
      n_0_253, n_0_252, n_0_251, n_0_250, n_0_249, n_0_248, n_0_247, n_0_246}), 
      .p_0({uc_325, in_a[15], in_a[14], in_a[13], in_a[12], in_a[11], in_a[10], 
      in_a[9], in_a[8], in_a[7], in_a[6], in_a[5], in_a[4], in_a[3], in_a[2], 
      in_a[1], in_a[0]}));
   DFFR_X1 zero_reg (.D(n_0_273), .RN(n_0_267), .CK(n_0_4), .Q(zero), .QN());
   DFFRS_X1 err_reg (.D(n_0_271), .RN(n_0_268), .SN(n_0_270), .CK(n_0_4), 
      .Q(err), .QN());
   DFFRS_X1 done_reg (.D(1'b1), .RN(n_0_266), .SN(n_0_264), .CK(n_0_4), .Q(done), 
      .QN());
   DFFR_X1 \out_c_reg[63]  (.D(n_0_282), .RN(n_0_267), .CK(n_0_4), .Q(out_c[16]), 
      .QN());
   DFFR_X1 \out_c_reg[15]  (.D(n_0_281), .RN(n_0_267), .CK(n_0_4), .Q(out_c[15]), 
      .QN());
   DFFR_X1 \out_c_reg[14]  (.D(n_0_280), .RN(n_0_267), .CK(n_0_4), .Q(out_c[14]), 
      .QN());
   DFFR_X1 \out_c_reg[13]  (.D(n_0_279), .RN(n_0_267), .CK(n_0_4), .Q(out_c[13]), 
      .QN());
   DFFR_X1 \out_c_reg[12]  (.D(n_0_278), .RN(n_0_267), .CK(n_0_4), .Q(out_c[12]), 
      .QN());
   DFFR_X1 \out_c_reg[11]  (.D(n_0_277), .RN(n_0_267), .CK(n_0_4), .Q(out_c[11]), 
      .QN());
   DFFR_X1 \out_c_reg[10]  (.D(n_0_276), .RN(n_0_267), .CK(n_0_4), .Q(out_c[10]), 
      .QN());
   DFFR_X1 \out_c_reg[9]  (.D(n_0_275), .RN(n_0_267), .CK(n_0_4), .Q(out_c[9]), 
      .QN());
   DFFR_X1 \out_c_reg[8]  (.D(n_0_274), .RN(n_0_267), .CK(n_0_4), .Q(out_c[8]), 
      .QN());
   DFFR_X1 \out_c_reg[7]  (.D(\output [14]), .RN(n_0_267), .CK(n_0_4), .Q(
      out_c[7]), .QN());
   DFFR_X1 \out_c_reg[6]  (.D(n_0_283), .RN(n_0_267), .CK(n_0_4), .Q(out_c[6]), 
      .QN());
   DFFR_X1 \out_c_reg[5]  (.D(n_0_301), .RN(n_0_267), .CK(n_0_4), .Q(out_c[5]), 
      .QN());
   DFFR_X1 \out_c_reg[4]  (.D(n_0_319), .RN(n_0_267), .CK(n_0_4), .Q(out_c[4]), 
      .QN());
   DFFR_X1 \out_c_reg[3]  (.D(n_0_337), .RN(n_0_267), .CK(n_0_4), .Q(out_c[3]), 
      .QN());
   DFFR_X1 \out_c_reg[2]  (.D(n_0_355), .RN(n_0_267), .CK(n_0_4), .Q(out_c[2]), 
      .QN());
   DFFR_X1 \out_c_reg[1]  (.D(n_0_373), .RN(n_0_267), .CK(n_0_4), .Q(out_c[1]), 
      .QN());
   DFFR_X1 \out_c_reg[0]  (.D(n_0_391), .RN(n_0_267), .CK(n_0_4), .Q(out_c[0]), 
      .QN());
   DFFR_X1 error_reg (.D(n_0_263), .RN(n_0_264), .CK(clk), .Q(error), .QN());
   MUX2_X1 error_reg_enable_mux_0 (.A(error), .B(n_0_271), .S(n_0_265), .Z(
      n_0_263));
   INV_X1 i_0_0_0 (.A(rst), .ZN(n_0_264));
   CLKGATETST_X1 clk_gate_posv_reg (.CK(clk), .E(n_0_269), .SE(1'b0), .GCK(n_0_4));
   NOR2_X1 i_0_1_0 (.A1(n_0_1_0), .A2(error), .ZN(n_0_265));
   AOI21_X1 i_0_1_1 (.A(rst), .B1(n_0_269), .B2(n_0_1_0), .ZN(n_0_268));
   NOR2_X1 i_0_1_2 (.A1(n_0_1_0), .A2(rst), .ZN(n_0_267));
   OR2_X1 i_0_1_3 (.A1(n_0_269), .A2(n_0_266), .ZN(n_0_270));
   OR2_X1 i_0_1_4 (.A1(rst), .A2(enbl), .ZN(n_0_266));
   INV_X1 i_0_1_5 (.A(enbl), .ZN(n_0_1_0));
   INV_X1 i_0_1_6 (.A(error), .ZN(n_0_269));
   AND2_X1 i_0_2_0 (.A1(in_b[0]), .A2(in_a[1]), .ZN(n_0_510));
   AND2_X1 i_0_2_1 (.A1(in_b[0]), .A2(in_a[2]), .ZN(n_0_511));
   AND2_X1 i_0_2_2 (.A1(in_b[0]), .A2(in_a[3]), .ZN(n_0_512));
   AND2_X1 i_0_2_3 (.A1(in_b[0]), .A2(in_a[4]), .ZN(n_0_513));
   AND2_X1 i_0_2_4 (.A1(in_b[0]), .A2(in_a[5]), .ZN(n_0_514));
   AND2_X1 i_0_2_5 (.A1(in_b[0]), .A2(in_a[6]), .ZN(n_0_515));
   AND2_X1 i_0_2_6 (.A1(in_b[0]), .A2(in_a[7]), .ZN(n_0_516));
   AND2_X1 i_0_2_7 (.A1(in_b[0]), .A2(in_a[8]), .ZN(n_0_517));
   AND2_X1 i_0_2_8 (.A1(in_b[0]), .A2(in_a[9]), .ZN(n_0_518));
   AND2_X1 i_0_2_9 (.A1(in_b[0]), .A2(in_a[10]), .ZN(n_0_519));
   AND2_X1 i_0_2_10 (.A1(in_b[0]), .A2(in_a[11]), .ZN(n_0_520));
   AND2_X1 i_0_2_11 (.A1(in_b[0]), .A2(in_a[12]), .ZN(n_0_521));
   AND2_X1 i_0_2_12 (.A1(in_b[0]), .A2(in_a[13]), .ZN(n_0_522));
   AND2_X1 i_0_2_13 (.A1(in_b[0]), .A2(in_a[14]), .ZN(n_0_523));
   AND2_X1 i_0_2_14 (.A1(in_b[0]), .A2(in_a[15]), .ZN(n_0_524));
   INV_X1 i_0_2_15 (.A(in_b[1]), .ZN(n_0_2_0));
   AOI22_X1 i_0_2_16 (.A1(n_0_2_0), .A2(n_0_511), .B1(in_b[1]), .B2(n_0_0), 
      .ZN(n_0_2_1));
   INV_X1 i_0_2_17 (.A(n_0_2_1), .ZN(n_0_494));
   AOI22_X1 i_0_2_18 (.A1(n_0_2_0), .A2(n_0_512), .B1(in_b[1]), .B2(n_0_1), 
      .ZN(n_0_2_2));
   INV_X1 i_0_2_19 (.A(n_0_2_2), .ZN(n_0_495));
   AOI22_X1 i_0_2_20 (.A1(n_0_2_0), .A2(n_0_513), .B1(in_b[1]), .B2(n_0_2), 
      .ZN(n_0_2_3));
   INV_X1 i_0_2_21 (.A(n_0_2_3), .ZN(n_0_496));
   AOI22_X1 i_0_2_22 (.A1(n_0_2_0), .A2(n_0_514), .B1(in_b[1]), .B2(n_0_3), 
      .ZN(n_0_2_4));
   INV_X1 i_0_2_23 (.A(n_0_2_4), .ZN(n_0_497));
   AOI22_X1 i_0_2_24 (.A1(n_0_2_0), .A2(n_0_515), .B1(in_b[1]), .B2(n_0_5), 
      .ZN(n_0_2_5));
   INV_X1 i_0_2_25 (.A(n_0_2_5), .ZN(n_0_498));
   AOI22_X1 i_0_2_26 (.A1(n_0_2_0), .A2(n_0_516), .B1(in_b[1]), .B2(n_0_6), 
      .ZN(n_0_2_6));
   INV_X1 i_0_2_27 (.A(n_0_2_6), .ZN(n_0_499));
   AOI22_X1 i_0_2_28 (.A1(n_0_2_0), .A2(n_0_517), .B1(in_b[1]), .B2(n_0_7), 
      .ZN(n_0_2_7));
   INV_X1 i_0_2_29 (.A(n_0_2_7), .ZN(n_0_500));
   AOI22_X1 i_0_2_30 (.A1(n_0_2_0), .A2(n_0_518), .B1(in_b[1]), .B2(n_0_8), 
      .ZN(n_0_2_8));
   INV_X1 i_0_2_31 (.A(n_0_2_8), .ZN(n_0_501));
   AOI22_X1 i_0_2_32 (.A1(n_0_2_0), .A2(n_0_519), .B1(in_b[1]), .B2(n_0_9), 
      .ZN(n_0_2_9));
   INV_X1 i_0_2_33 (.A(n_0_2_9), .ZN(n_0_502));
   AOI22_X1 i_0_2_34 (.A1(n_0_2_0), .A2(n_0_520), .B1(in_b[1]), .B2(n_0_10), 
      .ZN(n_0_2_10));
   INV_X1 i_0_2_35 (.A(n_0_2_10), .ZN(n_0_503));
   AOI22_X1 i_0_2_36 (.A1(n_0_2_0), .A2(n_0_521), .B1(in_b[1]), .B2(n_0_11), 
      .ZN(n_0_2_11));
   INV_X1 i_0_2_37 (.A(n_0_2_11), .ZN(n_0_504));
   AOI22_X1 i_0_2_38 (.A1(n_0_2_0), .A2(n_0_522), .B1(in_b[1]), .B2(n_0_12), 
      .ZN(n_0_2_12));
   INV_X1 i_0_2_39 (.A(n_0_2_12), .ZN(n_0_505));
   AOI22_X1 i_0_2_40 (.A1(n_0_2_0), .A2(n_0_523), .B1(in_b[1]), .B2(n_0_13), 
      .ZN(n_0_2_13));
   INV_X1 i_0_2_41 (.A(n_0_2_13), .ZN(n_0_506));
   NAND2_X1 i_0_2_42 (.A1(n_0_2_0), .A2(n_0_524), .ZN(n_0_2_14));
   NAND2_X1 i_0_2_43 (.A1(in_b[1]), .A2(n_0_14), .ZN(n_0_2_15));
   NAND2_X1 i_0_2_44 (.A1(n_0_2_14), .A2(n_0_2_15), .ZN(n_0_507));
   NAND2_X1 i_0_2_45 (.A1(in_b[1]), .A2(n_0_15), .ZN(n_0_2_16));
   NAND2_X1 i_0_2_46 (.A1(n_0_2_14), .A2(n_0_2_16), .ZN(n_0_508));
   NAND2_X1 i_0_2_47 (.A1(in_b[1]), .A2(n_0_16), .ZN(n_0_2_17));
   NAND2_X1 i_0_2_48 (.A1(n_0_2_14), .A2(n_0_2_17), .ZN(n_0_509));
   INV_X1 i_0_2_49 (.A(in_b[2]), .ZN(n_0_2_18));
   AOI22_X1 i_0_2_50 (.A1(n_0_2_18), .A2(n_0_495), .B1(in_b[2]), .B2(n_0_17), 
      .ZN(n_0_2_19));
   INV_X1 i_0_2_51 (.A(n_0_2_19), .ZN(n_0_477));
   AOI22_X1 i_0_2_52 (.A1(n_0_2_18), .A2(n_0_496), .B1(in_b[2]), .B2(n_0_18), 
      .ZN(n_0_2_20));
   INV_X1 i_0_2_53 (.A(n_0_2_20), .ZN(n_0_478));
   AOI22_X1 i_0_2_54 (.A1(n_0_2_18), .A2(n_0_497), .B1(in_b[2]), .B2(n_0_19), 
      .ZN(n_0_2_21));
   INV_X1 i_0_2_55 (.A(n_0_2_21), .ZN(n_0_479));
   AOI22_X1 i_0_2_56 (.A1(n_0_2_18), .A2(n_0_498), .B1(in_b[2]), .B2(n_0_20), 
      .ZN(n_0_2_22));
   INV_X1 i_0_2_57 (.A(n_0_2_22), .ZN(n_0_480));
   AOI22_X1 i_0_2_58 (.A1(n_0_2_18), .A2(n_0_499), .B1(in_b[2]), .B2(n_0_21), 
      .ZN(n_0_2_23));
   INV_X1 i_0_2_59 (.A(n_0_2_23), .ZN(n_0_481));
   AOI22_X1 i_0_2_60 (.A1(n_0_2_18), .A2(n_0_500), .B1(in_b[2]), .B2(n_0_22), 
      .ZN(n_0_2_24));
   INV_X1 i_0_2_61 (.A(n_0_2_24), .ZN(n_0_482));
   AOI22_X1 i_0_2_62 (.A1(n_0_2_18), .A2(n_0_501), .B1(in_b[2]), .B2(n_0_23), 
      .ZN(n_0_2_25));
   INV_X1 i_0_2_63 (.A(n_0_2_25), .ZN(n_0_483));
   AOI22_X1 i_0_2_64 (.A1(n_0_2_18), .A2(n_0_502), .B1(in_b[2]), .B2(n_0_24), 
      .ZN(n_0_2_26));
   INV_X1 i_0_2_65 (.A(n_0_2_26), .ZN(n_0_484));
   AOI22_X1 i_0_2_66 (.A1(n_0_2_18), .A2(n_0_503), .B1(in_b[2]), .B2(n_0_25), 
      .ZN(n_0_2_27));
   INV_X1 i_0_2_67 (.A(n_0_2_27), .ZN(n_0_485));
   AOI22_X1 i_0_2_68 (.A1(n_0_2_18), .A2(n_0_504), .B1(in_b[2]), .B2(n_0_26), 
      .ZN(n_0_2_28));
   INV_X1 i_0_2_69 (.A(n_0_2_28), .ZN(n_0_486));
   AOI22_X1 i_0_2_70 (.A1(n_0_2_18), .A2(n_0_505), .B1(in_b[2]), .B2(n_0_27), 
      .ZN(n_0_2_29));
   INV_X1 i_0_2_71 (.A(n_0_2_29), .ZN(n_0_487));
   AOI22_X1 i_0_2_72 (.A1(n_0_2_18), .A2(n_0_506), .B1(in_b[2]), .B2(n_0_28), 
      .ZN(n_0_2_30));
   INV_X1 i_0_2_73 (.A(n_0_2_30), .ZN(n_0_488));
   AOI22_X1 i_0_2_74 (.A1(n_0_2_18), .A2(n_0_507), .B1(in_b[2]), .B2(n_0_29), 
      .ZN(n_0_2_31));
   INV_X1 i_0_2_75 (.A(n_0_2_31), .ZN(n_0_489));
   AOI22_X1 i_0_2_76 (.A1(n_0_2_18), .A2(n_0_508), .B1(in_b[2]), .B2(n_0_30), 
      .ZN(n_0_2_32));
   INV_X1 i_0_2_77 (.A(n_0_2_32), .ZN(n_0_490));
   AOI22_X1 i_0_2_78 (.A1(n_0_2_18), .A2(n_0_509), .B1(in_b[2]), .B2(n_0_31), 
      .ZN(n_0_2_33));
   INV_X1 i_0_2_79 (.A(n_0_2_33), .ZN(n_0_491));
   AOI22_X1 i_0_2_80 (.A1(n_0_2_18), .A2(n_0_509), .B1(in_b[2]), .B2(n_0_32), 
      .ZN(n_0_2_34));
   INV_X1 i_0_2_81 (.A(n_0_2_34), .ZN(n_0_492));
   AOI22_X1 i_0_2_82 (.A1(n_0_2_18), .A2(n_0_509), .B1(in_b[2]), .B2(n_0_33), 
      .ZN(n_0_2_35));
   INV_X1 i_0_2_83 (.A(n_0_2_35), .ZN(n_0_493));
   MUX2_X1 i_0_2_84 (.A(n_0_478), .B(n_0_34), .S(in_b[3]), .Z(n_0_460));
   MUX2_X1 i_0_2_85 (.A(n_0_479), .B(n_0_35), .S(in_b[3]), .Z(n_0_461));
   MUX2_X1 i_0_2_86 (.A(n_0_480), .B(n_0_36), .S(in_b[3]), .Z(n_0_462));
   MUX2_X1 i_0_2_87 (.A(n_0_481), .B(n_0_37), .S(in_b[3]), .Z(n_0_463));
   MUX2_X1 i_0_2_88 (.A(n_0_482), .B(n_0_38), .S(in_b[3]), .Z(n_0_464));
   MUX2_X1 i_0_2_89 (.A(n_0_483), .B(n_0_39), .S(in_b[3]), .Z(n_0_465));
   MUX2_X1 i_0_2_90 (.A(n_0_484), .B(n_0_40), .S(in_b[3]), .Z(n_0_466));
   MUX2_X1 i_0_2_91 (.A(n_0_485), .B(n_0_41), .S(in_b[3]), .Z(n_0_467));
   MUX2_X1 i_0_2_92 (.A(n_0_486), .B(n_0_42), .S(in_b[3]), .Z(n_0_468));
   MUX2_X1 i_0_2_93 (.A(n_0_487), .B(n_0_43), .S(in_b[3]), .Z(n_0_469));
   MUX2_X1 i_0_2_94 (.A(n_0_488), .B(n_0_44), .S(in_b[3]), .Z(n_0_470));
   MUX2_X1 i_0_2_95 (.A(n_0_489), .B(n_0_45), .S(in_b[3]), .Z(n_0_471));
   MUX2_X1 i_0_2_96 (.A(n_0_490), .B(n_0_46), .S(in_b[3]), .Z(n_0_472));
   MUX2_X1 i_0_2_97 (.A(n_0_491), .B(n_0_47), .S(in_b[3]), .Z(n_0_473));
   MUX2_X1 i_0_2_98 (.A(n_0_492), .B(n_0_48), .S(in_b[3]), .Z(n_0_474));
   MUX2_X1 i_0_2_99 (.A(n_0_493), .B(n_0_49), .S(in_b[3]), .Z(n_0_475));
   MUX2_X1 i_0_2_100 (.A(n_0_493), .B(n_0_50), .S(in_b[3]), .Z(n_0_476));
   MUX2_X1 i_0_2_101 (.A(n_0_461), .B(n_0_51), .S(in_b[4]), .Z(n_0_443));
   MUX2_X1 i_0_2_102 (.A(n_0_462), .B(n_0_52), .S(in_b[4]), .Z(n_0_444));
   MUX2_X1 i_0_2_103 (.A(n_0_463), .B(n_0_53), .S(in_b[4]), .Z(n_0_445));
   MUX2_X1 i_0_2_104 (.A(n_0_464), .B(n_0_54), .S(in_b[4]), .Z(n_0_446));
   MUX2_X1 i_0_2_105 (.A(n_0_465), .B(n_0_55), .S(in_b[4]), .Z(n_0_447));
   MUX2_X1 i_0_2_106 (.A(n_0_466), .B(n_0_56), .S(in_b[4]), .Z(n_0_448));
   MUX2_X1 i_0_2_107 (.A(n_0_467), .B(n_0_57), .S(in_b[4]), .Z(n_0_449));
   MUX2_X1 i_0_2_108 (.A(n_0_468), .B(n_0_58), .S(in_b[4]), .Z(n_0_450));
   MUX2_X1 i_0_2_109 (.A(n_0_469), .B(n_0_59), .S(in_b[4]), .Z(n_0_451));
   MUX2_X1 i_0_2_110 (.A(n_0_470), .B(n_0_60), .S(in_b[4]), .Z(n_0_452));
   MUX2_X1 i_0_2_111 (.A(n_0_471), .B(n_0_61), .S(in_b[4]), .Z(n_0_453));
   MUX2_X1 i_0_2_112 (.A(n_0_472), .B(n_0_62), .S(in_b[4]), .Z(n_0_454));
   MUX2_X1 i_0_2_113 (.A(n_0_473), .B(n_0_63), .S(in_b[4]), .Z(n_0_455));
   MUX2_X1 i_0_2_114 (.A(n_0_474), .B(n_0_64), .S(in_b[4]), .Z(n_0_456));
   MUX2_X1 i_0_2_115 (.A(n_0_475), .B(n_0_65), .S(in_b[4]), .Z(n_0_457));
   MUX2_X1 i_0_2_116 (.A(n_0_476), .B(n_0_66), .S(in_b[4]), .Z(n_0_458));
   MUX2_X1 i_0_2_117 (.A(n_0_476), .B(n_0_67), .S(in_b[4]), .Z(n_0_459));
   MUX2_X1 i_0_2_118 (.A(n_0_444), .B(n_0_68), .S(in_b[5]), .Z(n_0_426));
   MUX2_X1 i_0_2_119 (.A(n_0_445), .B(n_0_69), .S(in_b[5]), .Z(n_0_427));
   MUX2_X1 i_0_2_120 (.A(n_0_446), .B(n_0_70), .S(in_b[5]), .Z(n_0_428));
   MUX2_X1 i_0_2_121 (.A(n_0_447), .B(n_0_71), .S(in_b[5]), .Z(n_0_429));
   MUX2_X1 i_0_2_122 (.A(n_0_448), .B(n_0_72), .S(in_b[5]), .Z(n_0_430));
   MUX2_X1 i_0_2_123 (.A(n_0_449), .B(n_0_73), .S(in_b[5]), .Z(n_0_431));
   MUX2_X1 i_0_2_124 (.A(n_0_450), .B(n_0_74), .S(in_b[5]), .Z(n_0_432));
   MUX2_X1 i_0_2_125 (.A(n_0_451), .B(n_0_75), .S(in_b[5]), .Z(n_0_433));
   MUX2_X1 i_0_2_126 (.A(n_0_452), .B(n_0_76), .S(in_b[5]), .Z(n_0_434));
   MUX2_X1 i_0_2_127 (.A(n_0_453), .B(n_0_77), .S(in_b[5]), .Z(n_0_435));
   MUX2_X1 i_0_2_128 (.A(n_0_454), .B(n_0_78), .S(in_b[5]), .Z(n_0_436));
   MUX2_X1 i_0_2_129 (.A(n_0_455), .B(n_0_79), .S(in_b[5]), .Z(n_0_437));
   MUX2_X1 i_0_2_130 (.A(n_0_456), .B(n_0_80), .S(in_b[5]), .Z(n_0_438));
   MUX2_X1 i_0_2_131 (.A(n_0_457), .B(n_0_81), .S(in_b[5]), .Z(n_0_439));
   MUX2_X1 i_0_2_132 (.A(n_0_458), .B(n_0_82), .S(in_b[5]), .Z(n_0_440));
   MUX2_X1 i_0_2_133 (.A(n_0_459), .B(n_0_83), .S(in_b[5]), .Z(n_0_441));
   MUX2_X1 i_0_2_134 (.A(n_0_459), .B(n_0_84), .S(in_b[5]), .Z(n_0_442));
   MUX2_X1 i_0_2_135 (.A(n_0_427), .B(n_0_85), .S(in_b[6]), .Z(n_0_409));
   MUX2_X1 i_0_2_136 (.A(n_0_428), .B(n_0_86), .S(in_b[6]), .Z(n_0_410));
   MUX2_X1 i_0_2_137 (.A(n_0_429), .B(n_0_87), .S(in_b[6]), .Z(n_0_411));
   MUX2_X1 i_0_2_138 (.A(n_0_430), .B(n_0_88), .S(in_b[6]), .Z(n_0_412));
   MUX2_X1 i_0_2_139 (.A(n_0_431), .B(n_0_89), .S(in_b[6]), .Z(n_0_413));
   MUX2_X1 i_0_2_140 (.A(n_0_432), .B(n_0_90), .S(in_b[6]), .Z(n_0_414));
   MUX2_X1 i_0_2_141 (.A(n_0_433), .B(n_0_91), .S(in_b[6]), .Z(n_0_415));
   MUX2_X1 i_0_2_142 (.A(n_0_434), .B(n_0_92), .S(in_b[6]), .Z(n_0_416));
   MUX2_X1 i_0_2_143 (.A(n_0_435), .B(n_0_93), .S(in_b[6]), .Z(n_0_417));
   MUX2_X1 i_0_2_144 (.A(n_0_436), .B(n_0_94), .S(in_b[6]), .Z(n_0_418));
   MUX2_X1 i_0_2_145 (.A(n_0_437), .B(n_0_95), .S(in_b[6]), .Z(n_0_419));
   MUX2_X1 i_0_2_146 (.A(n_0_438), .B(n_0_96), .S(in_b[6]), .Z(n_0_420));
   MUX2_X1 i_0_2_147 (.A(n_0_439), .B(n_0_97), .S(in_b[6]), .Z(n_0_421));
   MUX2_X1 i_0_2_148 (.A(n_0_440), .B(n_0_98), .S(in_b[6]), .Z(n_0_422));
   MUX2_X1 i_0_2_149 (.A(n_0_441), .B(n_0_99), .S(in_b[6]), .Z(n_0_423));
   MUX2_X1 i_0_2_150 (.A(n_0_442), .B(n_0_100), .S(in_b[6]), .Z(n_0_424));
   MUX2_X1 i_0_2_151 (.A(n_0_442), .B(n_0_101), .S(in_b[6]), .Z(n_0_425));
   MUX2_X1 i_0_2_152 (.A(n_0_409), .B(n_0_102), .S(in_b[7]), .Z(n_0_391));
   MUX2_X1 i_0_2_153 (.A(n_0_410), .B(n_0_103), .S(in_b[7]), .Z(n_0_392));
   MUX2_X1 i_0_2_154 (.A(n_0_411), .B(n_0_104), .S(in_b[7]), .Z(n_0_393));
   MUX2_X1 i_0_2_155 (.A(n_0_412), .B(n_0_105), .S(in_b[7]), .Z(n_0_394));
   MUX2_X1 i_0_2_156 (.A(n_0_413), .B(n_0_106), .S(in_b[7]), .Z(n_0_395));
   MUX2_X1 i_0_2_157 (.A(n_0_414), .B(n_0_107), .S(in_b[7]), .Z(n_0_396));
   MUX2_X1 i_0_2_158 (.A(n_0_415), .B(n_0_108), .S(in_b[7]), .Z(n_0_397));
   MUX2_X1 i_0_2_159 (.A(n_0_416), .B(n_0_109), .S(in_b[7]), .Z(n_0_398));
   MUX2_X1 i_0_2_160 (.A(n_0_417), .B(n_0_110), .S(in_b[7]), .Z(n_0_399));
   MUX2_X1 i_0_2_161 (.A(n_0_418), .B(n_0_111), .S(in_b[7]), .Z(n_0_400));
   MUX2_X1 i_0_2_162 (.A(n_0_419), .B(n_0_112), .S(in_b[7]), .Z(n_0_401));
   MUX2_X1 i_0_2_163 (.A(n_0_420), .B(n_0_113), .S(in_b[7]), .Z(n_0_402));
   MUX2_X1 i_0_2_164 (.A(n_0_421), .B(n_0_114), .S(in_b[7]), .Z(n_0_403));
   MUX2_X1 i_0_2_165 (.A(n_0_422), .B(n_0_115), .S(in_b[7]), .Z(n_0_404));
   MUX2_X1 i_0_2_166 (.A(n_0_423), .B(n_0_116), .S(in_b[7]), .Z(n_0_405));
   MUX2_X1 i_0_2_167 (.A(n_0_424), .B(n_0_117), .S(in_b[7]), .Z(n_0_406));
   MUX2_X1 i_0_2_168 (.A(n_0_425), .B(n_0_118), .S(in_b[7]), .Z(n_0_407));
   MUX2_X1 i_0_2_169 (.A(n_0_425), .B(n_0_119), .S(in_b[7]), .Z(n_0_408));
   MUX2_X1 i_0_2_170 (.A(n_0_392), .B(n_0_120), .S(in_b[8]), .Z(n_0_373));
   MUX2_X1 i_0_2_171 (.A(n_0_393), .B(n_0_121), .S(in_b[8]), .Z(n_0_374));
   MUX2_X1 i_0_2_172 (.A(n_0_394), .B(n_0_122), .S(in_b[8]), .Z(n_0_375));
   MUX2_X1 i_0_2_173 (.A(n_0_395), .B(n_0_123), .S(in_b[8]), .Z(n_0_376));
   MUX2_X1 i_0_2_174 (.A(n_0_396), .B(n_0_124), .S(in_b[8]), .Z(n_0_377));
   MUX2_X1 i_0_2_175 (.A(n_0_397), .B(n_0_125), .S(in_b[8]), .Z(n_0_378));
   MUX2_X1 i_0_2_176 (.A(n_0_398), .B(n_0_126), .S(in_b[8]), .Z(n_0_379));
   MUX2_X1 i_0_2_177 (.A(n_0_399), .B(n_0_127), .S(in_b[8]), .Z(n_0_380));
   MUX2_X1 i_0_2_178 (.A(n_0_400), .B(n_0_128), .S(in_b[8]), .Z(n_0_381));
   MUX2_X1 i_0_2_179 (.A(n_0_401), .B(n_0_129), .S(in_b[8]), .Z(n_0_382));
   MUX2_X1 i_0_2_180 (.A(n_0_402), .B(n_0_130), .S(in_b[8]), .Z(n_0_383));
   MUX2_X1 i_0_2_181 (.A(n_0_403), .B(n_0_131), .S(in_b[8]), .Z(n_0_384));
   MUX2_X1 i_0_2_182 (.A(n_0_404), .B(n_0_132), .S(in_b[8]), .Z(n_0_385));
   MUX2_X1 i_0_2_183 (.A(n_0_405), .B(n_0_133), .S(in_b[8]), .Z(n_0_386));
   MUX2_X1 i_0_2_184 (.A(n_0_406), .B(n_0_134), .S(in_b[8]), .Z(n_0_387));
   MUX2_X1 i_0_2_185 (.A(n_0_407), .B(n_0_135), .S(in_b[8]), .Z(n_0_388));
   MUX2_X1 i_0_2_186 (.A(n_0_408), .B(n_0_136), .S(in_b[8]), .Z(n_0_389));
   MUX2_X1 i_0_2_187 (.A(n_0_408), .B(n_0_137), .S(in_b[8]), .Z(n_0_390));
   MUX2_X1 i_0_2_188 (.A(n_0_374), .B(n_0_138), .S(in_b[9]), .Z(n_0_355));
   MUX2_X1 i_0_2_189 (.A(n_0_375), .B(n_0_139), .S(in_b[9]), .Z(n_0_356));
   MUX2_X1 i_0_2_190 (.A(n_0_376), .B(n_0_140), .S(in_b[9]), .Z(n_0_357));
   MUX2_X1 i_0_2_191 (.A(n_0_377), .B(n_0_141), .S(in_b[9]), .Z(n_0_358));
   MUX2_X1 i_0_2_192 (.A(n_0_378), .B(n_0_142), .S(in_b[9]), .Z(n_0_359));
   MUX2_X1 i_0_2_193 (.A(n_0_379), .B(n_0_143), .S(in_b[9]), .Z(n_0_360));
   MUX2_X1 i_0_2_194 (.A(n_0_380), .B(n_0_144), .S(in_b[9]), .Z(n_0_361));
   MUX2_X1 i_0_2_195 (.A(n_0_381), .B(n_0_145), .S(in_b[9]), .Z(n_0_362));
   MUX2_X1 i_0_2_196 (.A(n_0_382), .B(n_0_146), .S(in_b[9]), .Z(n_0_363));
   MUX2_X1 i_0_2_197 (.A(n_0_383), .B(n_0_147), .S(in_b[9]), .Z(n_0_364));
   MUX2_X1 i_0_2_198 (.A(n_0_384), .B(n_0_148), .S(in_b[9]), .Z(n_0_365));
   MUX2_X1 i_0_2_199 (.A(n_0_385), .B(n_0_149), .S(in_b[9]), .Z(n_0_366));
   MUX2_X1 i_0_2_200 (.A(n_0_386), .B(n_0_150), .S(in_b[9]), .Z(n_0_367));
   MUX2_X1 i_0_2_201 (.A(n_0_387), .B(n_0_151), .S(in_b[9]), .Z(n_0_368));
   MUX2_X1 i_0_2_202 (.A(n_0_388), .B(n_0_152), .S(in_b[9]), .Z(n_0_369));
   MUX2_X1 i_0_2_203 (.A(n_0_389), .B(n_0_153), .S(in_b[9]), .Z(n_0_370));
   MUX2_X1 i_0_2_204 (.A(n_0_390), .B(n_0_154), .S(in_b[9]), .Z(n_0_371));
   MUX2_X1 i_0_2_205 (.A(n_0_390), .B(n_0_155), .S(in_b[9]), .Z(n_0_372));
   MUX2_X1 i_0_2_206 (.A(n_0_356), .B(n_0_156), .S(in_b[10]), .Z(n_0_337));
   MUX2_X1 i_0_2_207 (.A(n_0_357), .B(n_0_157), .S(in_b[10]), .Z(n_0_338));
   MUX2_X1 i_0_2_208 (.A(n_0_358), .B(n_0_158), .S(in_b[10]), .Z(n_0_339));
   MUX2_X1 i_0_2_209 (.A(n_0_359), .B(n_0_159), .S(in_b[10]), .Z(n_0_340));
   MUX2_X1 i_0_2_210 (.A(n_0_360), .B(n_0_160), .S(in_b[10]), .Z(n_0_341));
   MUX2_X1 i_0_2_211 (.A(n_0_361), .B(n_0_161), .S(in_b[10]), .Z(n_0_342));
   MUX2_X1 i_0_2_212 (.A(n_0_362), .B(n_0_162), .S(in_b[10]), .Z(n_0_343));
   MUX2_X1 i_0_2_213 (.A(n_0_363), .B(n_0_163), .S(in_b[10]), .Z(n_0_344));
   MUX2_X1 i_0_2_214 (.A(n_0_364), .B(n_0_164), .S(in_b[10]), .Z(n_0_345));
   MUX2_X1 i_0_2_215 (.A(n_0_365), .B(n_0_165), .S(in_b[10]), .Z(n_0_346));
   MUX2_X1 i_0_2_216 (.A(n_0_366), .B(n_0_166), .S(in_b[10]), .Z(n_0_347));
   MUX2_X1 i_0_2_217 (.A(n_0_367), .B(n_0_167), .S(in_b[10]), .Z(n_0_348));
   MUX2_X1 i_0_2_218 (.A(n_0_368), .B(n_0_168), .S(in_b[10]), .Z(n_0_349));
   MUX2_X1 i_0_2_219 (.A(n_0_369), .B(n_0_169), .S(in_b[10]), .Z(n_0_350));
   MUX2_X1 i_0_2_220 (.A(n_0_370), .B(n_0_170), .S(in_b[10]), .Z(n_0_351));
   MUX2_X1 i_0_2_221 (.A(n_0_371), .B(n_0_171), .S(in_b[10]), .Z(n_0_352));
   MUX2_X1 i_0_2_222 (.A(n_0_372), .B(n_0_172), .S(in_b[10]), .Z(n_0_353));
   MUX2_X1 i_0_2_223 (.A(n_0_372), .B(n_0_173), .S(in_b[10]), .Z(n_0_354));
   MUX2_X1 i_0_2_224 (.A(n_0_338), .B(n_0_174), .S(in_b[11]), .Z(n_0_319));
   MUX2_X1 i_0_2_225 (.A(n_0_339), .B(n_0_175), .S(in_b[11]), .Z(n_0_320));
   MUX2_X1 i_0_2_226 (.A(n_0_340), .B(n_0_176), .S(in_b[11]), .Z(n_0_321));
   MUX2_X1 i_0_2_227 (.A(n_0_341), .B(n_0_177), .S(in_b[11]), .Z(n_0_322));
   MUX2_X1 i_0_2_228 (.A(n_0_342), .B(n_0_178), .S(in_b[11]), .Z(n_0_323));
   MUX2_X1 i_0_2_229 (.A(n_0_343), .B(n_0_179), .S(in_b[11]), .Z(n_0_324));
   MUX2_X1 i_0_2_230 (.A(n_0_344), .B(n_0_180), .S(in_b[11]), .Z(n_0_325));
   MUX2_X1 i_0_2_231 (.A(n_0_345), .B(n_0_181), .S(in_b[11]), .Z(n_0_326));
   MUX2_X1 i_0_2_232 (.A(n_0_346), .B(n_0_182), .S(in_b[11]), .Z(n_0_327));
   MUX2_X1 i_0_2_233 (.A(n_0_347), .B(n_0_183), .S(in_b[11]), .Z(n_0_328));
   MUX2_X1 i_0_2_234 (.A(n_0_348), .B(n_0_184), .S(in_b[11]), .Z(n_0_329));
   MUX2_X1 i_0_2_235 (.A(n_0_349), .B(n_0_185), .S(in_b[11]), .Z(n_0_330));
   MUX2_X1 i_0_2_236 (.A(n_0_350), .B(n_0_186), .S(in_b[11]), .Z(n_0_331));
   MUX2_X1 i_0_2_237 (.A(n_0_351), .B(n_0_187), .S(in_b[11]), .Z(n_0_332));
   MUX2_X1 i_0_2_238 (.A(n_0_352), .B(n_0_188), .S(in_b[11]), .Z(n_0_333));
   MUX2_X1 i_0_2_239 (.A(n_0_353), .B(n_0_189), .S(in_b[11]), .Z(n_0_334));
   MUX2_X1 i_0_2_240 (.A(n_0_354), .B(n_0_190), .S(in_b[11]), .Z(n_0_335));
   MUX2_X1 i_0_2_241 (.A(n_0_354), .B(n_0_191), .S(in_b[11]), .Z(n_0_336));
   MUX2_X1 i_0_2_242 (.A(n_0_320), .B(n_0_192), .S(in_b[12]), .Z(n_0_301));
   MUX2_X1 i_0_2_243 (.A(n_0_321), .B(n_0_193), .S(in_b[12]), .Z(n_0_302));
   MUX2_X1 i_0_2_244 (.A(n_0_322), .B(n_0_194), .S(in_b[12]), .Z(n_0_303));
   MUX2_X1 i_0_2_245 (.A(n_0_323), .B(n_0_195), .S(in_b[12]), .Z(n_0_304));
   MUX2_X1 i_0_2_246 (.A(n_0_324), .B(n_0_196), .S(in_b[12]), .Z(n_0_305));
   MUX2_X1 i_0_2_247 (.A(n_0_325), .B(n_0_197), .S(in_b[12]), .Z(n_0_306));
   MUX2_X1 i_0_2_248 (.A(n_0_326), .B(n_0_198), .S(in_b[12]), .Z(n_0_307));
   MUX2_X1 i_0_2_249 (.A(n_0_327), .B(n_0_199), .S(in_b[12]), .Z(n_0_308));
   MUX2_X1 i_0_2_250 (.A(n_0_328), .B(n_0_200), .S(in_b[12]), .Z(n_0_309));
   MUX2_X1 i_0_2_251 (.A(n_0_329), .B(n_0_201), .S(in_b[12]), .Z(n_0_310));
   MUX2_X1 i_0_2_252 (.A(n_0_330), .B(n_0_202), .S(in_b[12]), .Z(n_0_311));
   MUX2_X1 i_0_2_253 (.A(n_0_331), .B(n_0_203), .S(in_b[12]), .Z(n_0_312));
   MUX2_X1 i_0_2_254 (.A(n_0_332), .B(n_0_204), .S(in_b[12]), .Z(n_0_313));
   MUX2_X1 i_0_2_255 (.A(n_0_333), .B(n_0_205), .S(in_b[12]), .Z(n_0_314));
   MUX2_X1 i_0_2_256 (.A(n_0_334), .B(n_0_206), .S(in_b[12]), .Z(n_0_315));
   MUX2_X1 i_0_2_257 (.A(n_0_335), .B(n_0_207), .S(in_b[12]), .Z(n_0_316));
   MUX2_X1 i_0_2_258 (.A(n_0_336), .B(n_0_208), .S(in_b[12]), .Z(n_0_317));
   MUX2_X1 i_0_2_259 (.A(n_0_336), .B(n_0_209), .S(in_b[12]), .Z(n_0_318));
   MUX2_X1 i_0_2_260 (.A(n_0_302), .B(n_0_210), .S(in_b[13]), .Z(n_0_283));
   MUX2_X1 i_0_2_261 (.A(n_0_303), .B(n_0_211), .S(in_b[13]), .Z(n_0_284));
   MUX2_X1 i_0_2_262 (.A(n_0_304), .B(n_0_212), .S(in_b[13]), .Z(n_0_285));
   MUX2_X1 i_0_2_263 (.A(n_0_305), .B(n_0_213), .S(in_b[13]), .Z(n_0_286));
   MUX2_X1 i_0_2_264 (.A(n_0_306), .B(n_0_214), .S(in_b[13]), .Z(n_0_287));
   MUX2_X1 i_0_2_265 (.A(n_0_307), .B(n_0_215), .S(in_b[13]), .Z(n_0_288));
   MUX2_X1 i_0_2_266 (.A(n_0_308), .B(n_0_216), .S(in_b[13]), .Z(n_0_289));
   MUX2_X1 i_0_2_267 (.A(n_0_309), .B(n_0_217), .S(in_b[13]), .Z(n_0_290));
   MUX2_X1 i_0_2_268 (.A(n_0_310), .B(n_0_218), .S(in_b[13]), .Z(n_0_291));
   MUX2_X1 i_0_2_269 (.A(n_0_311), .B(n_0_219), .S(in_b[13]), .Z(n_0_292));
   MUX2_X1 i_0_2_270 (.A(n_0_312), .B(n_0_220), .S(in_b[13]), .Z(n_0_293));
   MUX2_X1 i_0_2_271 (.A(n_0_313), .B(n_0_221), .S(in_b[13]), .Z(n_0_294));
   MUX2_X1 i_0_2_272 (.A(n_0_314), .B(n_0_222), .S(in_b[13]), .Z(n_0_295));
   MUX2_X1 i_0_2_273 (.A(n_0_315), .B(n_0_223), .S(in_b[13]), .Z(n_0_296));
   MUX2_X1 i_0_2_274 (.A(n_0_316), .B(n_0_224), .S(in_b[13]), .Z(n_0_297));
   MUX2_X1 i_0_2_275 (.A(n_0_317), .B(n_0_225), .S(in_b[13]), .Z(n_0_298));
   MUX2_X1 i_0_2_276 (.A(n_0_318), .B(n_0_226), .S(in_b[13]), .Z(n_0_299));
   MUX2_X1 i_0_2_277 (.A(n_0_318), .B(n_0_227), .S(in_b[13]), .Z(n_0_300));
   MUX2_X1 i_0_2_278 (.A(n_0_284), .B(n_0_228), .S(in_b[14]), .Z(\output [14]));
   MUX2_X1 i_0_2_279 (.A(n_0_285), .B(n_0_229), .S(in_b[14]), .Z(\output [15]));
   MUX2_X1 i_0_2_280 (.A(n_0_286), .B(n_0_230), .S(in_b[14]), .Z(\output [16]));
   MUX2_X1 i_0_2_281 (.A(n_0_287), .B(n_0_231), .S(in_b[14]), .Z(\output [17]));
   MUX2_X1 i_0_2_282 (.A(n_0_288), .B(n_0_232), .S(in_b[14]), .Z(\output [18]));
   MUX2_X1 i_0_2_283 (.A(n_0_289), .B(n_0_233), .S(in_b[14]), .Z(\output [19]));
   MUX2_X1 i_0_2_284 (.A(n_0_290), .B(n_0_234), .S(in_b[14]), .Z(\output [20]));
   MUX2_X1 i_0_2_285 (.A(n_0_291), .B(n_0_235), .S(in_b[14]), .Z(\output [21]));
   MUX2_X1 i_0_2_286 (.A(n_0_292), .B(n_0_236), .S(in_b[14]), .Z(\output [22]));
   MUX2_X1 i_0_2_287 (.A(n_0_293), .B(n_0_237), .S(in_b[14]), .Z(\output [23]));
   MUX2_X1 i_0_2_288 (.A(n_0_294), .B(n_0_238), .S(in_b[14]), .Z(\output [24]));
   MUX2_X1 i_0_2_289 (.A(n_0_295), .B(n_0_239), .S(in_b[14]), .Z(\output [25]));
   MUX2_X1 i_0_2_290 (.A(n_0_296), .B(n_0_240), .S(in_b[14]), .Z(\output [26]));
   MUX2_X1 i_0_2_291 (.A(n_0_297), .B(n_0_241), .S(in_b[14]), .Z(\output [27]));
   MUX2_X1 i_0_2_292 (.A(n_0_298), .B(n_0_242), .S(in_b[14]), .Z(\output [28]));
   MUX2_X1 i_0_2_293 (.A(n_0_299), .B(n_0_243), .S(in_b[14]), .Z(\output [29]));
   MUX2_X1 i_0_2_294 (.A(n_0_300), .B(n_0_244), .S(in_b[14]), .Z(\output [30]));
   MUX2_X1 i_0_2_295 (.A(n_0_300), .B(n_0_245), .S(in_b[14]), .Z(\output [31]));
   MUX2_X1 i_0_2_296 (.A(\output [15]), .B(n_0_246), .S(in_b[15]), .Z(n_0_274));
   MUX2_X1 i_0_2_297 (.A(\output [16]), .B(n_0_247), .S(in_b[15]), .Z(n_0_275));
   MUX2_X1 i_0_2_298 (.A(\output [17]), .B(n_0_248), .S(in_b[15]), .Z(n_0_276));
   MUX2_X1 i_0_2_299 (.A(\output [18]), .B(n_0_249), .S(in_b[15]), .Z(n_0_277));
   MUX2_X1 i_0_2_300 (.A(\output [19]), .B(n_0_250), .S(in_b[15]), .Z(n_0_278));
   MUX2_X1 i_0_2_301 (.A(\output [20]), .B(n_0_251), .S(in_b[15]), .Z(n_0_279));
   MUX2_X1 i_0_2_302 (.A(\output [21]), .B(n_0_252), .S(in_b[15]), .Z(n_0_280));
   MUX2_X1 i_0_2_303 (.A(\output [22]), .B(n_0_253), .S(in_b[15]), .Z(n_0_281));
   MUX2_X1 i_0_2_304 (.A(\output [23]), .B(n_0_254), .S(in_b[15]), .Z(n_0_2_46));
   MUX2_X1 i_0_2_305 (.A(\output [24]), .B(n_0_255), .S(in_b[15]), .Z(n_0_2_47));
   MUX2_X1 i_0_2_306 (.A(\output [25]), .B(n_0_256), .S(in_b[15]), .Z(n_0_2_48));
   MUX2_X1 i_0_2_307 (.A(\output [26]), .B(n_0_257), .S(in_b[15]), .Z(n_0_2_49));
   MUX2_X1 i_0_2_308 (.A(\output [27]), .B(n_0_258), .S(in_b[15]), .Z(n_0_2_50));
   MUX2_X1 i_0_2_309 (.A(\output [28]), .B(n_0_259), .S(in_b[15]), .Z(n_0_2_51));
   MUX2_X1 i_0_2_310 (.A(\output [29]), .B(n_0_260), .S(in_b[15]), .Z(n_0_2_52));
   MUX2_X1 i_0_2_311 (.A(\output [30]), .B(n_0_261), .S(in_b[15]), .Z(n_0_2_53));
   MUX2_X1 i_0_2_312 (.A(\output [31]), .B(n_0_262), .S(in_b[15]), .Z(n_0_282));
   NOR4_X1 i_0_2_313 (.A1(n_0_391), .A2(n_0_373), .A3(n_0_355), .A4(n_0_337), 
      .ZN(n_0_2_36));
   NOR4_X1 i_0_2_314 (.A1(n_0_319), .A2(n_0_301), .A3(n_0_283), .A4(\output [14]), 
      .ZN(n_0_2_37));
   NOR4_X1 i_0_2_315 (.A1(n_0_274), .A2(n_0_275), .A3(n_0_276), .A4(n_0_277), 
      .ZN(n_0_2_38));
   NOR4_X1 i_0_2_316 (.A1(n_0_278), .A2(n_0_279), .A3(n_0_280), .A4(n_0_281), 
      .ZN(n_0_2_39));
   AND4_X1 i_0_2_317 (.A1(n_0_2_36), .A2(n_0_2_37), .A3(n_0_2_38), .A4(n_0_2_39), 
      .ZN(n_0_273));
   NOR2_X1 i_0_2_318 (.A1(n_0_274), .A2(n_0_273), .ZN(n_0_272));
   AND4_X1 i_0_2_319 (.A1(n_0_2_48), .A2(n_0_2_49), .A3(n_0_2_47), .A4(n_0_281), 
      .ZN(n_0_2_40));
   AND4_X1 i_0_2_320 (.A1(n_0_2_40), .A2(n_0_2_52), .A3(n_0_2_53), .A4(n_0_2_51), 
      .ZN(n_0_2_41));
   AND4_X1 i_0_2_321 (.A1(n_0_2_41), .A2(n_0_282), .A3(n_0_2_46), .A4(n_0_2_50), 
      .ZN(n_0_2_42));
   OR4_X1 i_0_2_322 (.A1(n_0_2_48), .A2(n_0_2_49), .A3(n_0_2_47), .A4(n_0_281), 
      .ZN(n_0_2_43));
   OR4_X1 i_0_2_323 (.A1(n_0_2_43), .A2(n_0_2_52), .A3(n_0_2_53), .A4(n_0_2_51), 
      .ZN(n_0_2_44));
   NOR4_X1 i_0_2_324 (.A1(n_0_2_44), .A2(n_0_282), .A3(n_0_2_46), .A4(n_0_2_50), 
      .ZN(n_0_2_45));
   NOR2_X1 i_0_2_325 (.A1(n_0_2_42), .A2(n_0_2_45), .ZN(n_0_271));
endmodule
