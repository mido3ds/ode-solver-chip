library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.common.all;
use work.solver_pkg.all;


entity solver_test is
    generic (
        WORD_LENGTH : integer := 32;
        ADDR_LENGTH : integer := 16;
        MAX_LENGTH  : integer := 64
    );

    port (
        --in_state       : in std_logic_vector(1 downto 0); --state signal sent from CPU
        clk            : in std_logic;
        rst            : in std_logic;
       -- interp_done_op : in std_logic_vector(1 downto 0);
        in_data        : inout std_logic_vector(WORD_LENGTH - 1 downto 0);
        adr            : inout std_logic_vector(ADDR_LENGTH - 1 downto 0)
        --interrupt      : out std_logic;
        --error_success  : out std_logic
    );
end entity;

architecture rtl of solver_test is
    signal X_intm_rd,first_time, X_intm_wr : std_logic    := '0';
    signal X_intm_address : std_logic_vector(6 downto 0) := (others => '0');
    signal X_intm_data_in, X_intm_data_out : std_logic_vector(WORD_LENGTH - 1 downto 0) := (others => '0');
    signal fsm_write : std_logic_vector(1 downto 0) := (others => '0');

    signal x_temp,x_temp_3 : std_logic_vector(63 downto 0) := (others => '1');
    signal x_temp_2 : std_logic_vector(63 downto 0) := X"1111111122222222";
    
    signal main_fsm, fsm_out : std_logic_vector(2 downto 0) := (others => '0');
    signal N_counter: std_logic_vector(5 downto 0) := "000101";
    signal N_counter_2: std_logic_vector(5 downto 0) := (others => '0');
    signal mode_sig : std_logic_vector(1 downto 0) := "10";
    signal wares : std_logic_vector(2 downto 0) := "001";
    signal procedure_dumm : std_logic_vector(10 downto 0) := (others => '0');
   
    begin
    X_i : entity work.ram generic map (WORD_LENGTH => WORD_LENGTH, NUM_WORDS => 100, ADR_LENGTH=>7)
        port map(
            clk      => clk,
            rd       => X_intm_rd,
            wr       => X_intm_wr,
            address  => X_intm_address,
            data_in  => X_intm_data_in,
            data_out => X_intm_data_out,
            rst      => rst
        );
    
    main_proc : process(clk, rst)
    begin
        if rst = '0' and rising_edge(clk) then
            --Fill X_i with data..
            case( main_fsm ) is
            
                when "000" =>
                    x_temp_2 <= to_vec(to_int(x_temp_2) + 1234567,64);
                    fsm_write <= "11";
                    main_fsm <= "001";

                when "001" =>
                    write_after_read_reg (
                            data_in => x_temp_2,
                            reg_data_in => X_intm_data_in,
                            reg_adrs => X_intm_address,
                            read_enbl => X_intm_rd,
                            write_enbl => X_intm_wr,
                            fsm => fsm_write
                        );

                    if fsm_write = "00" then 
                        main_fsm <= "010";
                        N_counter_2 <= to_vec(to_int(N_counter_2) + 1,6);
                    end if;

                when "010"=>
                    if N_counter_2 = N_counter then
                        main_fsm <= "011";
                        fsm_out <= "111";
                    else
                        fsm_write <= "11";
                        main_fsm <= "001";
                    end if;

                when "011" =>

                    outing(
                        mode => mode_sig,
                        main_adr => adr,
                        data_bus => in_data,
                        x_ware_data_out => X_intm_data_out,
                        x_ware_address => X_intm_address,
                        read_enbl => X_intm_rd,
                        write_enbl => X_intm_wr,
                        c_ware => wares,
                        fsm => fsm_out,
                        N_X_A_B => N_counter,
                        fsm_read => procedure_dumm(10 downto 9),
                        N_X_A_B_counter => procedure_dumm(8 downto 3),
                        c_ware_vec => procedure_dumm(2 downto 0)
                    );
                    if fsm_out = "000" then
                        main_fsm <= "000";
                    end if;
                when others =>
            
            end case ;
            
        end if;
    end process ;
    
    

end architecture;

