/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sat Apr 25 22:08:49 2020
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 1180132999 */

module datapath(in_b_signal, in_a, p_0);
   input [63:0]in_b_signal;
   input [63:0]in_a;
   output [63:0]p_0;

   HA_X1 i_0 (.A(in_b_signal[0]), .B(in_a[0]), .CO(n_0), .S(p_0[0]));
   FA_X1 i_1 (.A(in_b_signal[1]), .B(in_a[1]), .CI(n_0), .CO(n_1), .S(p_0[1]));
   FA_X1 i_2 (.A(in_b_signal[2]), .B(in_a[2]), .CI(n_1), .CO(n_2), .S(p_0[2]));
   FA_X1 i_3 (.A(in_b_signal[3]), .B(in_a[3]), .CI(n_2), .CO(n_3), .S(p_0[3]));
   FA_X1 i_4 (.A(in_b_signal[4]), .B(in_a[4]), .CI(n_3), .CO(n_4), .S(p_0[4]));
   FA_X1 i_5 (.A(in_b_signal[5]), .B(in_a[5]), .CI(n_4), .CO(n_5), .S(p_0[5]));
   FA_X1 i_6 (.A(in_b_signal[6]), .B(in_a[6]), .CI(n_5), .CO(n_6), .S(p_0[6]));
   FA_X1 i_7 (.A(in_b_signal[7]), .B(in_a[7]), .CI(n_6), .CO(n_7), .S(p_0[7]));
   FA_X1 i_8 (.A(in_b_signal[8]), .B(in_a[8]), .CI(n_7), .CO(n_8), .S(p_0[8]));
   FA_X1 i_9 (.A(in_b_signal[9]), .B(in_a[9]), .CI(n_8), .CO(n_9), .S(p_0[9]));
   FA_X1 i_10 (.A(in_b_signal[10]), .B(in_a[10]), .CI(n_9), .CO(n_10), .S(
      p_0[10]));
   FA_X1 i_11 (.A(in_b_signal[11]), .B(in_a[11]), .CI(n_10), .CO(n_11), .S(
      p_0[11]));
   FA_X1 i_12 (.A(in_b_signal[12]), .B(in_a[12]), .CI(n_11), .CO(n_12), .S(
      p_0[12]));
   FA_X1 i_13 (.A(in_b_signal[13]), .B(in_a[13]), .CI(n_12), .CO(n_13), .S(
      p_0[13]));
   FA_X1 i_14 (.A(in_b_signal[14]), .B(in_a[14]), .CI(n_13), .CO(n_14), .S(
      p_0[14]));
   FA_X1 i_15 (.A(in_b_signal[15]), .B(in_a[15]), .CI(n_14), .CO(n_15), .S(
      p_0[15]));
   FA_X1 i_16 (.A(in_b_signal[16]), .B(in_a[16]), .CI(n_15), .CO(n_16), .S(
      p_0[16]));
   FA_X1 i_17 (.A(in_b_signal[17]), .B(in_a[17]), .CI(n_16), .CO(n_17), .S(
      p_0[17]));
   FA_X1 i_18 (.A(in_b_signal[18]), .B(in_a[18]), .CI(n_17), .CO(n_18), .S(
      p_0[18]));
   FA_X1 i_19 (.A(in_b_signal[19]), .B(in_a[19]), .CI(n_18), .CO(n_19), .S(
      p_0[19]));
   FA_X1 i_20 (.A(in_b_signal[20]), .B(in_a[20]), .CI(n_19), .CO(n_20), .S(
      p_0[20]));
   FA_X1 i_21 (.A(in_b_signal[21]), .B(in_a[21]), .CI(n_20), .CO(n_21), .S(
      p_0[21]));
   FA_X1 i_22 (.A(in_b_signal[22]), .B(in_a[22]), .CI(n_21), .CO(n_22), .S(
      p_0[22]));
   FA_X1 i_23 (.A(in_b_signal[23]), .B(in_a[23]), .CI(n_22), .CO(n_23), .S(
      p_0[23]));
   FA_X1 i_24 (.A(in_b_signal[24]), .B(in_a[24]), .CI(n_23), .CO(n_24), .S(
      p_0[24]));
   FA_X1 i_25 (.A(in_b_signal[25]), .B(in_a[25]), .CI(n_24), .CO(n_25), .S(
      p_0[25]));
   FA_X1 i_26 (.A(in_b_signal[26]), .B(in_a[26]), .CI(n_25), .CO(n_26), .S(
      p_0[26]));
   FA_X1 i_27 (.A(in_b_signal[27]), .B(in_a[27]), .CI(n_26), .CO(n_27), .S(
      p_0[27]));
   FA_X1 i_28 (.A(in_b_signal[28]), .B(in_a[28]), .CI(n_27), .CO(n_28), .S(
      p_0[28]));
   FA_X1 i_29 (.A(in_b_signal[29]), .B(in_a[29]), .CI(n_28), .CO(n_29), .S(
      p_0[29]));
   FA_X1 i_30 (.A(in_b_signal[30]), .B(in_a[30]), .CI(n_29), .CO(n_30), .S(
      p_0[30]));
   FA_X1 i_31 (.A(in_b_signal[31]), .B(in_a[31]), .CI(n_30), .CO(n_31), .S(
      p_0[31]));
   FA_X1 i_32 (.A(in_b_signal[32]), .B(in_a[32]), .CI(n_31), .CO(n_32), .S(
      p_0[32]));
   FA_X1 i_33 (.A(in_b_signal[33]), .B(in_a[33]), .CI(n_32), .CO(n_33), .S(
      p_0[33]));
   FA_X1 i_34 (.A(in_b_signal[34]), .B(in_a[34]), .CI(n_33), .CO(n_34), .S(
      p_0[34]));
   FA_X1 i_35 (.A(in_b_signal[35]), .B(in_a[35]), .CI(n_34), .CO(n_35), .S(
      p_0[35]));
   FA_X1 i_36 (.A(in_b_signal[36]), .B(in_a[36]), .CI(n_35), .CO(n_36), .S(
      p_0[36]));
   FA_X1 i_37 (.A(in_b_signal[37]), .B(in_a[37]), .CI(n_36), .CO(n_37), .S(
      p_0[37]));
   FA_X1 i_38 (.A(in_b_signal[38]), .B(in_a[38]), .CI(n_37), .CO(n_38), .S(
      p_0[38]));
   FA_X1 i_39 (.A(in_b_signal[39]), .B(in_a[39]), .CI(n_38), .CO(n_39), .S(
      p_0[39]));
   FA_X1 i_40 (.A(in_b_signal[40]), .B(in_a[40]), .CI(n_39), .CO(n_40), .S(
      p_0[40]));
   FA_X1 i_41 (.A(in_b_signal[41]), .B(in_a[41]), .CI(n_40), .CO(n_41), .S(
      p_0[41]));
   FA_X1 i_42 (.A(in_b_signal[42]), .B(in_a[42]), .CI(n_41), .CO(n_42), .S(
      p_0[42]));
   FA_X1 i_43 (.A(in_b_signal[43]), .B(in_a[43]), .CI(n_42), .CO(n_43), .S(
      p_0[43]));
   FA_X1 i_44 (.A(in_b_signal[44]), .B(in_a[44]), .CI(n_43), .CO(n_44), .S(
      p_0[44]));
   FA_X1 i_45 (.A(in_b_signal[45]), .B(in_a[45]), .CI(n_44), .CO(n_45), .S(
      p_0[45]));
   FA_X1 i_46 (.A(in_b_signal[46]), .B(in_a[46]), .CI(n_45), .CO(n_46), .S(
      p_0[46]));
   FA_X1 i_47 (.A(in_b_signal[47]), .B(in_a[47]), .CI(n_46), .CO(n_47), .S(
      p_0[47]));
   FA_X1 i_48 (.A(in_b_signal[48]), .B(in_a[48]), .CI(n_47), .CO(n_48), .S(
      p_0[48]));
   FA_X1 i_49 (.A(in_b_signal[49]), .B(in_a[49]), .CI(n_48), .CO(n_49), .S(
      p_0[49]));
   FA_X1 i_50 (.A(in_b_signal[50]), .B(in_a[50]), .CI(n_49), .CO(n_50), .S(
      p_0[50]));
   FA_X1 i_51 (.A(in_b_signal[51]), .B(in_a[51]), .CI(n_50), .CO(n_51), .S(
      p_0[51]));
   FA_X1 i_52 (.A(in_b_signal[52]), .B(in_a[52]), .CI(n_51), .CO(n_52), .S(
      p_0[52]));
   FA_X1 i_53 (.A(in_b_signal[53]), .B(in_a[53]), .CI(n_52), .CO(n_53), .S(
      p_0[53]));
   FA_X1 i_54 (.A(in_b_signal[54]), .B(in_a[54]), .CI(n_53), .CO(n_54), .S(
      p_0[54]));
   FA_X1 i_55 (.A(in_b_signal[55]), .B(in_a[55]), .CI(n_54), .CO(n_55), .S(
      p_0[55]));
   FA_X1 i_56 (.A(in_b_signal[56]), .B(in_a[56]), .CI(n_55), .CO(n_56), .S(
      p_0[56]));
   FA_X1 i_57 (.A(in_b_signal[57]), .B(in_a[57]), .CI(n_56), .CO(n_57), .S(
      p_0[57]));
   FA_X1 i_58 (.A(in_b_signal[58]), .B(in_a[58]), .CI(n_57), .CO(n_58), .S(
      p_0[58]));
   FA_X1 i_59 (.A(in_b_signal[59]), .B(in_a[59]), .CI(n_58), .CO(n_59), .S(
      p_0[59]));
   FA_X1 i_60 (.A(in_b_signal[60]), .B(in_a[60]), .CI(n_59), .CO(n_60), .S(
      p_0[60]));
   FA_X1 i_61 (.A(in_b_signal[61]), .B(in_a[61]), .CI(n_60), .CO(n_61), .S(
      p_0[61]));
   FA_X1 i_62 (.A(in_b_signal[62]), .B(in_a[62]), .CI(n_61), .CO(n_62), .S(
      p_0[62]));
   XNOR2_X1 i_63 (.A(in_b_signal[63]), .B(in_a[63]), .ZN(n_63));
   XNOR2_X1 i_64 (.A(n_63), .B(n_62), .ZN(p_0[63]));
endmodule

module datapath__0_6(plus, in_b);
   output [63:0]plus;
   input [63:0]in_b;

   XOR2_X1 i_0 (.A(in_b[1]), .B(in_b[0]), .Z(plus[1]));
   AND2_X1 i_1 (.A1(n_61), .A2(n_0), .ZN(plus[2]));
   OAI21_X1 i_2 (.A(in_b[2]), .B1(in_b[1]), .B2(in_b[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(in_b[3]), .B(n_61), .Z(plus[3]));
   XOR2_X1 i_4 (.A(in_b[4]), .B(n_60), .Z(plus[4]));
   XOR2_X1 i_5 (.A(in_b[5]), .B(n_59), .Z(plus[5]));
   AND2_X1 i_6 (.A1(n_58), .A2(n_1), .ZN(plus[6]));
   OAI21_X1 i_7 (.A(in_b[6]), .B1(n_59), .B2(in_b[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(in_b[7]), .B(n_58), .Z(plus[7]));
   XOR2_X1 i_9 (.A(in_b[8]), .B(n_57), .Z(plus[8]));
   AND2_X1 i_10 (.A1(n_56), .A2(n_2), .ZN(plus[9]));
   OAI21_X1 i_11 (.A(in_b[9]), .B1(n_57), .B2(in_b[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(in_b[10]), .B(n_56), .Z(plus[10]));
   XNOR2_X1 i_13 (.A(in_b[11]), .B(n_55), .ZN(plus[11]));
   XOR2_X1 i_14 (.A(in_b[12]), .B(n_54), .Z(plus[12]));
   XNOR2_X1 i_15 (.A(in_b[13]), .B(n_53), .ZN(plus[13]));
   XOR2_X1 i_16 (.A(in_b[14]), .B(n_52), .Z(plus[14]));
   AND2_X1 i_17 (.A1(n_51), .A2(n_3), .ZN(plus[15]));
   OAI21_X1 i_18 (.A(in_b[15]), .B1(n_52), .B2(in_b[14]), .ZN(n_3));
   XOR2_X1 i_19 (.A(in_b[16]), .B(n_51), .Z(plus[16]));
   XOR2_X1 i_20 (.A(in_b[17]), .B(n_50), .Z(plus[17]));
   XOR2_X1 i_21 (.A(in_b[18]), .B(n_49), .Z(plus[18]));
   XNOR2_X1 i_22 (.A(in_b[19]), .B(n_48), .ZN(plus[19]));
   XNOR2_X1 i_23 (.A(in_b[20]), .B(n_47), .ZN(plus[20]));
   XNOR2_X1 i_24 (.A(in_b[21]), .B(n_46), .ZN(plus[21]));
   XOR2_X1 i_25 (.A(in_b[22]), .B(n_45), .Z(plus[22]));
   XOR2_X1 i_26 (.A(in_b[23]), .B(n_44), .Z(plus[23]));
   XNOR2_X1 i_27 (.A(in_b[24]), .B(n_43), .ZN(plus[24]));
   XNOR2_X1 i_28 (.A(in_b[25]), .B(n_42), .ZN(plus[25]));
   XNOR2_X1 i_29 (.A(in_b[26]), .B(n_41), .ZN(plus[26]));
   XOR2_X1 i_30 (.A(in_b[27]), .B(n_40), .Z(plus[27]));
   XOR2_X1 i_31 (.A(in_b[28]), .B(n_39), .Z(plus[28]));
   XNOR2_X1 i_32 (.A(in_b[29]), .B(n_38), .ZN(plus[29]));
   XNOR2_X1 i_33 (.A(in_b[30]), .B(n_37), .ZN(plus[30]));
   XNOR2_X1 i_34 (.A(in_b[31]), .B(n_36), .ZN(plus[31]));
   XOR2_X1 i_35 (.A(in_b[32]), .B(n_35), .Z(plus[32]));
   XOR2_X1 i_36 (.A(in_b[33]), .B(n_34), .Z(plus[33]));
   XNOR2_X1 i_37 (.A(in_b[34]), .B(n_33), .ZN(plus[34]));
   XNOR2_X1 i_38 (.A(in_b[35]), .B(n_32), .ZN(plus[35]));
   XNOR2_X1 i_39 (.A(in_b[36]), .B(n_31), .ZN(plus[36]));
   XOR2_X1 i_40 (.A(in_b[37]), .B(n_30), .Z(plus[37]));
   XOR2_X1 i_41 (.A(in_b[38]), .B(n_29), .Z(plus[38]));
   XNOR2_X1 i_42 (.A(in_b[39]), .B(n_28), .ZN(plus[39]));
   XNOR2_X1 i_43 (.A(in_b[40]), .B(n_27), .ZN(plus[40]));
   XOR2_X1 i_44 (.A(in_b[41]), .B(n_26), .Z(plus[41]));
   XNOR2_X1 i_45 (.A(in_b[42]), .B(n_25), .ZN(plus[42]));
   XOR2_X1 i_46 (.A(in_b[43]), .B(n_24), .Z(plus[43]));
   AND2_X1 i_47 (.A1(n_23), .A2(n_4), .ZN(plus[44]));
   OAI21_X1 i_48 (.A(in_b[44]), .B1(n_24), .B2(in_b[43]), .ZN(n_4));
   XOR2_X1 i_49 (.A(in_b[45]), .B(n_23), .Z(plus[45]));
   XOR2_X1 i_50 (.A(in_b[46]), .B(n_22), .Z(plus[46]));
   XOR2_X1 i_51 (.A(in_b[47]), .B(n_21), .Z(plus[47]));
   XOR2_X1 i_52 (.A(in_b[48]), .B(n_20), .Z(plus[48]));
   XNOR2_X1 i_53 (.A(in_b[49]), .B(n_19), .ZN(plus[49]));
   XNOR2_X1 i_54 (.A(in_b[50]), .B(n_18), .ZN(plus[50]));
   XNOR2_X1 i_55 (.A(in_b[51]), .B(n_17), .ZN(plus[51]));
   XOR2_X1 i_56 (.A(in_b[52]), .B(n_16), .Z(plus[52]));
   XNOR2_X1 i_57 (.A(in_b[53]), .B(n_15), .ZN(plus[53]));
   XNOR2_X1 i_58 (.A(in_b[54]), .B(n_14), .ZN(plus[54]));
   XNOR2_X1 i_59 (.A(in_b[55]), .B(n_13), .ZN(plus[55]));
   XOR2_X1 i_60 (.A(in_b[56]), .B(n_12), .Z(plus[56]));
   AND2_X1 i_61 (.A1(n_11), .A2(n_5), .ZN(plus[57]));
   OAI21_X1 i_62 (.A(in_b[57]), .B1(n_12), .B2(in_b[56]), .ZN(n_5));
   XOR2_X1 i_63 (.A(in_b[58]), .B(n_11), .Z(plus[58]));
   XNOR2_X1 i_64 (.A(in_b[59]), .B(n_10), .ZN(plus[59]));
   XNOR2_X1 i_65 (.A(in_b[60]), .B(n_9), .ZN(plus[60]));
   XOR2_X1 i_66 (.A(in_b[61]), .B(n_8), .Z(plus[61]));
   XNOR2_X1 i_67 (.A(in_b[62]), .B(n_7), .ZN(plus[62]));
   XNOR2_X1 i_68 (.A(in_b[63]), .B(n_6), .ZN(plus[63]));
   NOR3_X1 i_69 (.A1(n_8), .A2(in_b[61]), .A3(in_b[62]), .ZN(n_6));
   NOR2_X1 i_70 (.A1(n_8), .A2(in_b[61]), .ZN(n_7));
   NAND2_X1 i_71 (.A1(n_9), .A2(n_72), .ZN(n_8));
   NOR3_X1 i_72 (.A1(n_11), .A2(in_b[58]), .A3(in_b[59]), .ZN(n_9));
   NOR2_X1 i_73 (.A1(n_11), .A2(in_b[58]), .ZN(n_10));
   OR3_X1 i_74 (.A1(n_12), .A2(in_b[56]), .A3(in_b[57]), .ZN(n_11));
   NAND2_X1 i_75 (.A1(n_13), .A2(n_71), .ZN(n_12));
   NOR4_X1 i_76 (.A1(n_16), .A2(in_b[52]), .A3(in_b[53]), .A4(in_b[54]), 
      .ZN(n_13));
   NOR3_X1 i_77 (.A1(n_16), .A2(in_b[52]), .A3(in_b[53]), .ZN(n_14));
   NOR2_X1 i_78 (.A1(n_16), .A2(in_b[52]), .ZN(n_15));
   NAND2_X1 i_79 (.A1(n_17), .A2(n_70), .ZN(n_16));
   NOR4_X1 i_80 (.A1(n_20), .A2(in_b[48]), .A3(in_b[49]), .A4(in_b[50]), 
      .ZN(n_17));
   NOR3_X1 i_81 (.A1(n_20), .A2(in_b[48]), .A3(in_b[49]), .ZN(n_18));
   NOR2_X1 i_82 (.A1(n_20), .A2(in_b[48]), .ZN(n_19));
   OR2_X1 i_83 (.A1(n_21), .A2(in_b[47]), .ZN(n_20));
   OR2_X1 i_84 (.A1(n_22), .A2(in_b[46]), .ZN(n_21));
   OR2_X1 i_85 (.A1(n_23), .A2(in_b[45]), .ZN(n_22));
   OR3_X1 i_86 (.A1(n_24), .A2(in_b[43]), .A3(in_b[44]), .ZN(n_23));
   NAND2_X1 i_87 (.A1(n_25), .A2(n_69), .ZN(n_24));
   NOR2_X1 i_88 (.A1(n_26), .A2(in_b[41]), .ZN(n_25));
   NAND2_X1 i_89 (.A1(n_27), .A2(n_68), .ZN(n_26));
   NOR3_X1 i_90 (.A1(n_29), .A2(in_b[38]), .A3(in_b[39]), .ZN(n_27));
   NOR2_X1 i_91 (.A1(n_29), .A2(in_b[38]), .ZN(n_28));
   OR2_X1 i_92 (.A1(n_30), .A2(in_b[37]), .ZN(n_29));
   NAND2_X1 i_93 (.A1(n_31), .A2(n_67), .ZN(n_30));
   NOR4_X1 i_94 (.A1(n_34), .A2(in_b[33]), .A3(in_b[34]), .A4(in_b[35]), 
      .ZN(n_31));
   NOR3_X1 i_95 (.A1(n_34), .A2(in_b[33]), .A3(in_b[34]), .ZN(n_32));
   NOR2_X1 i_96 (.A1(n_34), .A2(in_b[33]), .ZN(n_33));
   OR2_X1 i_97 (.A1(n_35), .A2(in_b[32]), .ZN(n_34));
   NAND2_X1 i_98 (.A1(n_36), .A2(n_66), .ZN(n_35));
   NOR4_X1 i_99 (.A1(n_39), .A2(in_b[28]), .A3(in_b[29]), .A4(in_b[30]), 
      .ZN(n_36));
   NOR3_X1 i_100 (.A1(n_39), .A2(in_b[28]), .A3(in_b[29]), .ZN(n_37));
   NOR2_X1 i_101 (.A1(n_39), .A2(in_b[28]), .ZN(n_38));
   OR2_X1 i_102 (.A1(n_40), .A2(in_b[27]), .ZN(n_39));
   NAND2_X1 i_103 (.A1(n_41), .A2(n_65), .ZN(n_40));
   NOR4_X1 i_104 (.A1(n_44), .A2(in_b[23]), .A3(in_b[24]), .A4(in_b[25]), 
      .ZN(n_41));
   NOR3_X1 i_105 (.A1(n_44), .A2(in_b[23]), .A3(in_b[24]), .ZN(n_42));
   NOR2_X1 i_106 (.A1(n_44), .A2(in_b[23]), .ZN(n_43));
   OR2_X1 i_107 (.A1(n_45), .A2(in_b[22]), .ZN(n_44));
   NAND2_X1 i_108 (.A1(n_46), .A2(n_64), .ZN(n_45));
   NOR4_X1 i_109 (.A1(n_49), .A2(in_b[18]), .A3(in_b[19]), .A4(in_b[20]), 
      .ZN(n_46));
   NOR3_X1 i_110 (.A1(n_49), .A2(in_b[18]), .A3(in_b[19]), .ZN(n_47));
   NOR2_X1 i_111 (.A1(n_49), .A2(in_b[18]), .ZN(n_48));
   OR2_X1 i_112 (.A1(n_50), .A2(in_b[17]), .ZN(n_49));
   OR2_X1 i_113 (.A1(n_51), .A2(in_b[16]), .ZN(n_50));
   OR3_X1 i_114 (.A1(n_52), .A2(in_b[14]), .A3(in_b[15]), .ZN(n_51));
   NAND2_X1 i_115 (.A1(n_53), .A2(n_63), .ZN(n_52));
   NOR2_X1 i_116 (.A1(n_54), .A2(in_b[12]), .ZN(n_53));
   NAND2_X1 i_117 (.A1(n_55), .A2(n_62), .ZN(n_54));
   NOR2_X1 i_118 (.A1(n_56), .A2(in_b[10]), .ZN(n_55));
   OR3_X1 i_119 (.A1(n_57), .A2(in_b[8]), .A3(in_b[9]), .ZN(n_56));
   OR2_X1 i_120 (.A1(n_58), .A2(in_b[7]), .ZN(n_57));
   OR3_X1 i_121 (.A1(n_59), .A2(in_b[5]), .A3(in_b[6]), .ZN(n_58));
   OR2_X1 i_122 (.A1(n_60), .A2(in_b[4]), .ZN(n_59));
   OR2_X1 i_123 (.A1(n_61), .A2(in_b[3]), .ZN(n_60));
   OR3_X1 i_124 (.A1(in_b[2]), .A2(in_b[1]), .A3(in_b[0]), .ZN(n_61));
   INV_X1 i_125 (.A(in_b[11]), .ZN(n_62));
   INV_X1 i_126 (.A(in_b[13]), .ZN(n_63));
   INV_X1 i_127 (.A(in_b[21]), .ZN(n_64));
   INV_X1 i_128 (.A(in_b[26]), .ZN(n_65));
   INV_X1 i_129 (.A(in_b[31]), .ZN(n_66));
   INV_X1 i_130 (.A(in_b[36]), .ZN(n_67));
   INV_X1 i_131 (.A(in_b[40]), .ZN(n_68));
   INV_X1 i_132 (.A(in_b[42]), .ZN(n_69));
   INV_X1 i_133 (.A(in_b[51]), .ZN(n_70));
   INV_X1 i_134 (.A(in_b[55]), .ZN(n_71));
   INV_X1 i_135 (.A(in_b[60]), .ZN(n_72));
endmodule

module fpu_adder(mode, clk, rst, enbl, add_sub, in_a, in_b, out_c, done, err, 
      zero, posv);
   input [1:0]mode;
   input clk;
   input rst;
   input enbl;
   input add_sub;
   input [63:0]in_a;
   input [63:0]in_b;
   output [63:0]out_c;
   output done;
   output err;
   output zero;
   output posv;

   wire F59;
   wire F58;
   wire F57;
   wire F56;
   wire F55;
   wire F54;
   wire F53;
   wire F52;
   wire F51;
   wire F50;
   wire F49;
   wire F48;
   wire F47;
   wire F46;
   wire F45;
   wire F44;
   wire F43;
   wire F42;
   wire F41;
   wire F40;
   wire F39;
   wire F38;
   wire F37;
   wire F36;
   wire F35;
   wire F34;
   wire F33;
   wire F32;
   wire F31;
   wire F30;
   wire F29;
   wire F28;
   wire F27;
   wire F26;
   wire F25;
   wire F24;
   wire F23;
   wire F22;
   wire F21;
   wire F20;
   wire F19;
   wire F18;
   wire F17;
   wire F16;
   wire F15;
   wire F14;
   wire F13;
   wire F12;
   wire F11;
   wire F10;
   wire F9;
   wire F8;
   wire F7;
   wire F6;
   wire F5;
   wire F4;
   wire F3;
   wire F2;
   wire F1;
   wire F0;
   wire F;

   DLH_X1 \out_c_signal_reg[63]  (.D(n_70), .G(n_71), .Q(n_4));
   DLH_X1 \out_c_signal_reg[62]  (.D(n_69), .G(n_71), .Q(n_5));
   DLH_X1 \out_c_signal_reg[61]  (.D(n_68), .G(n_71), .Q(F59));
   DLH_X1 \out_c_signal_reg[60]  (.D(n_67), .G(n_71), .Q(F58));
   DLH_X1 \out_c_signal_reg[59]  (.D(n_66), .G(n_71), .Q(F57));
   DLH_X1 \out_c_signal_reg[58]  (.D(n_65), .G(n_71), .Q(F56));
   DLH_X1 \out_c_signal_reg[57]  (.D(n_64), .G(n_71), .Q(F55));
   DLH_X1 \out_c_signal_reg[56]  (.D(n_63), .G(n_71), .Q(F54));
   DLH_X1 \out_c_signal_reg[55]  (.D(n_62), .G(n_71), .Q(F53));
   DLH_X1 \out_c_signal_reg[54]  (.D(n_61), .G(n_71), .Q(F52));
   DLH_X1 \out_c_signal_reg[53]  (.D(n_60), .G(n_71), .Q(F51));
   DLH_X1 \out_c_signal_reg[52]  (.D(n_59), .G(n_71), .Q(F50));
   DLH_X1 \out_c_signal_reg[51]  (.D(n_58), .G(n_71), .Q(F49));
   DLH_X1 \out_c_signal_reg[50]  (.D(n_57), .G(n_71), .Q(F48));
   DLH_X1 \out_c_signal_reg[49]  (.D(n_56), .G(n_71), .Q(F47));
   DLH_X1 \out_c_signal_reg[48]  (.D(n_55), .G(n_71), .Q(F46));
   DLH_X1 \out_c_signal_reg[47]  (.D(n_54), .G(n_71), .Q(F45));
   DLH_X1 \out_c_signal_reg[46]  (.D(n_53), .G(n_71), .Q(F44));
   DLH_X1 \out_c_signal_reg[45]  (.D(n_52), .G(n_71), .Q(F43));
   DLH_X1 \out_c_signal_reg[44]  (.D(n_51), .G(n_71), .Q(F42));
   DLH_X1 \out_c_signal_reg[43]  (.D(n_50), .G(n_71), .Q(F41));
   DLH_X1 \out_c_signal_reg[42]  (.D(n_49), .G(n_71), .Q(F40));
   DLH_X1 \out_c_signal_reg[41]  (.D(n_48), .G(n_71), .Q(F39));
   DLH_X1 \out_c_signal_reg[40]  (.D(n_47), .G(n_71), .Q(F38));
   DLH_X1 \out_c_signal_reg[39]  (.D(n_46), .G(n_71), .Q(F37));
   DLH_X1 \out_c_signal_reg[38]  (.D(n_45), .G(n_71), .Q(F36));
   DLH_X1 \out_c_signal_reg[37]  (.D(n_44), .G(n_71), .Q(F35));
   DLH_X1 \out_c_signal_reg[36]  (.D(n_43), .G(n_71), .Q(F34));
   DLH_X1 \out_c_signal_reg[35]  (.D(n_42), .G(n_71), .Q(F33));
   DLH_X1 \out_c_signal_reg[34]  (.D(n_41), .G(n_71), .Q(F32));
   DLH_X1 \out_c_signal_reg[33]  (.D(n_40), .G(n_71), .Q(F31));
   DLH_X1 \out_c_signal_reg[32]  (.D(n_39), .G(n_71), .Q(F30));
   DLH_X1 \out_c_signal_reg[31]  (.D(n_38), .G(n_71), .Q(F29));
   DLH_X1 \out_c_signal_reg[30]  (.D(n_37), .G(n_71), .Q(F28));
   DLH_X1 \out_c_signal_reg[29]  (.D(n_36), .G(n_71), .Q(F27));
   DLH_X1 \out_c_signal_reg[28]  (.D(n_35), .G(n_71), .Q(F26));
   DLH_X1 \out_c_signal_reg[27]  (.D(n_34), .G(n_71), .Q(F25));
   DLH_X1 \out_c_signal_reg[26]  (.D(n_33), .G(n_71), .Q(F24));
   DLH_X1 \out_c_signal_reg[25]  (.D(n_32), .G(n_71), .Q(F23));
   DLH_X1 \out_c_signal_reg[24]  (.D(n_31), .G(n_71), .Q(F22));
   DLH_X1 \out_c_signal_reg[23]  (.D(n_30), .G(n_71), .Q(F21));
   DLH_X1 \out_c_signal_reg[22]  (.D(n_29), .G(n_71), .Q(F20));
   DLH_X1 \out_c_signal_reg[21]  (.D(n_28), .G(n_71), .Q(F19));
   DLH_X1 \out_c_signal_reg[20]  (.D(n_27), .G(n_71), .Q(F18));
   DLH_X1 \out_c_signal_reg[19]  (.D(n_26), .G(n_71), .Q(F17));
   DLH_X1 \out_c_signal_reg[18]  (.D(n_25), .G(n_71), .Q(F16));
   DLH_X1 \out_c_signal_reg[17]  (.D(n_24), .G(n_71), .Q(F15));
   DLH_X1 \out_c_signal_reg[16]  (.D(n_23), .G(n_71), .Q(F14));
   DLH_X1 \out_c_signal_reg[15]  (.D(n_22), .G(n_71), .Q(F13));
   DLH_X1 \out_c_signal_reg[14]  (.D(n_21), .G(n_71), .Q(F12));
   DLH_X1 \out_c_signal_reg[13]  (.D(n_20), .G(n_71), .Q(F11));
   DLH_X1 \out_c_signal_reg[12]  (.D(n_19), .G(n_71), .Q(F10));
   DLH_X1 \out_c_signal_reg[11]  (.D(n_18), .G(n_71), .Q(F9));
   DLH_X1 \out_c_signal_reg[10]  (.D(n_17), .G(n_71), .Q(F8));
   DLH_X1 \out_c_signal_reg[9]  (.D(n_16), .G(n_71), .Q(F7));
   DLH_X1 \out_c_signal_reg[8]  (.D(n_15), .G(n_71), .Q(F6));
   DLH_X1 \out_c_signal_reg[7]  (.D(n_14), .G(n_71), .Q(F5));
   DLH_X1 \out_c_signal_reg[6]  (.D(n_13), .G(n_71), .Q(F4));
   DLH_X1 \out_c_signal_reg[5]  (.D(n_12), .G(n_71), .Q(F3));
   DLH_X1 \out_c_signal_reg[4]  (.D(n_11), .G(n_71), .Q(F2));
   DLH_X1 \out_c_signal_reg[3]  (.D(n_10), .G(n_71), .Q(F1));
   DLH_X1 \out_c_signal_reg[2]  (.D(n_9), .G(n_71), .Q(F0));
   DLH_X1 \out_c_signal_reg[1]  (.D(n_8), .G(n_71), .Q(F));
   DLH_X1 \out_c_signal_reg[0]  (.D(n_7), .G(n_71), .Q(n_6));
   datapath i_7 (.in_b_signal({n_72, n_73, n_74, n_75, n_76, n_77, n_78, n_79, 
      n_80, n_81, n_82, n_83, n_84, n_85, n_86, n_87, n_88, n_89, n_90, n_91, 
      n_92, n_93, n_94, n_95, n_96, n_97, n_98, n_99, n_100, n_101, n_102, n_103, 
      n_104, n_105, n_106, n_107, n_108, n_109, n_110, n_111, n_112, n_113, 
      n_114, n_115, n_116, n_117, n_118, n_119, n_120, n_121, n_122, n_123, 
      n_124, n_125, n_126, n_127, n_128, n_129, n_130, n_131, n_132, n_133, 
      n_134, n_135}), .in_a(in_a), .p_0({n_70, n_69, n_68, n_67, n_66, n_65, 
      n_64, n_63, n_62, n_61, n_60, n_59, n_58, n_57, n_56, n_55, n_54, n_53, 
      n_52, n_51, n_50, n_49, n_48, n_47, n_46, n_45, n_44, n_43, n_42, n_41, 
      n_40, n_39, n_38, n_37, n_36, n_35, n_34, n_33, n_32, n_31, n_30, n_29, 
      n_28, n_27, n_26, n_25, n_24, n_23, n_22, n_21, n_20, n_19, n_18, n_17, 
      n_16, n_15, n_14, n_13, n_12, n_11, n_10, n_9, n_8, n_7}));
   DLH_X1 \in_b_signal_reg[63]  (.D(n_3), .G(n_71), .Q(n_72));
   DLH_X1 \in_b_signal_reg[62]  (.D(n_2), .G(n_71), .Q(n_73));
   DLH_X1 \in_b_signal_reg[61]  (.D(n_1), .G(n_71), .Q(n_74));
   DLH_X1 \in_b_signal_reg[60]  (.D(n_0), .G(n_71), .Q(n_75));
   DLH_X1 \in_b_signal_reg[59]  (.D(n_194), .G(n_71), .Q(n_76));
   DLH_X1 \in_b_signal_reg[58]  (.D(n_193), .G(n_71), .Q(n_77));
   DLH_X1 \in_b_signal_reg[57]  (.D(n_192), .G(n_71), .Q(n_78));
   DLH_X1 \in_b_signal_reg[56]  (.D(n_191), .G(n_71), .Q(n_79));
   DLH_X1 \in_b_signal_reg[55]  (.D(n_190), .G(n_71), .Q(n_80));
   DLH_X1 \in_b_signal_reg[54]  (.D(n_189), .G(n_71), .Q(n_81));
   DLH_X1 \in_b_signal_reg[53]  (.D(n_188), .G(n_71), .Q(n_82));
   DLH_X1 \in_b_signal_reg[52]  (.D(n_187), .G(n_71), .Q(n_83));
   DLH_X1 \in_b_signal_reg[51]  (.D(n_186), .G(n_71), .Q(n_84));
   DLH_X1 \in_b_signal_reg[50]  (.D(n_185), .G(n_71), .Q(n_85));
   DLH_X1 \in_b_signal_reg[49]  (.D(n_184), .G(n_71), .Q(n_86));
   DLH_X1 \in_b_signal_reg[48]  (.D(n_183), .G(n_71), .Q(n_87));
   DLH_X1 \in_b_signal_reg[47]  (.D(n_182), .G(n_71), .Q(n_88));
   DLH_X1 \in_b_signal_reg[46]  (.D(n_181), .G(n_71), .Q(n_89));
   DLH_X1 \in_b_signal_reg[45]  (.D(n_180), .G(n_71), .Q(n_90));
   DLH_X1 \in_b_signal_reg[44]  (.D(n_179), .G(n_71), .Q(n_91));
   DLH_X1 \in_b_signal_reg[43]  (.D(n_178), .G(n_71), .Q(n_92));
   DLH_X1 \in_b_signal_reg[42]  (.D(n_177), .G(n_71), .Q(n_93));
   DLH_X1 \in_b_signal_reg[41]  (.D(n_176), .G(n_71), .Q(n_94));
   DLH_X1 \in_b_signal_reg[40]  (.D(n_175), .G(n_71), .Q(n_95));
   DLH_X1 \in_b_signal_reg[39]  (.D(n_174), .G(n_71), .Q(n_96));
   DLH_X1 \in_b_signal_reg[38]  (.D(n_173), .G(n_71), .Q(n_97));
   DLH_X1 \in_b_signal_reg[37]  (.D(n_172), .G(n_71), .Q(n_98));
   DLH_X1 \in_b_signal_reg[36]  (.D(n_171), .G(n_71), .Q(n_99));
   DLH_X1 \in_b_signal_reg[35]  (.D(n_170), .G(n_71), .Q(n_100));
   DLH_X1 \in_b_signal_reg[34]  (.D(n_169), .G(n_71), .Q(n_101));
   DLH_X1 \in_b_signal_reg[33]  (.D(n_168), .G(n_71), .Q(n_102));
   DLH_X1 \in_b_signal_reg[32]  (.D(n_167), .G(n_71), .Q(n_103));
   DLH_X1 \in_b_signal_reg[31]  (.D(n_166), .G(n_71), .Q(n_104));
   DLH_X1 \in_b_signal_reg[30]  (.D(n_165), .G(n_71), .Q(n_105));
   DLH_X1 \in_b_signal_reg[29]  (.D(n_164), .G(n_71), .Q(n_106));
   DLH_X1 \in_b_signal_reg[28]  (.D(n_163), .G(n_71), .Q(n_107));
   DLH_X1 \in_b_signal_reg[27]  (.D(n_162), .G(n_71), .Q(n_108));
   DLH_X1 \in_b_signal_reg[26]  (.D(n_161), .G(n_71), .Q(n_109));
   DLH_X1 \in_b_signal_reg[25]  (.D(n_160), .G(n_71), .Q(n_110));
   DLH_X1 \in_b_signal_reg[24]  (.D(n_159), .G(n_71), .Q(n_111));
   DLH_X1 \in_b_signal_reg[23]  (.D(n_158), .G(n_71), .Q(n_112));
   DLH_X1 \in_b_signal_reg[22]  (.D(n_157), .G(n_71), .Q(n_113));
   DLH_X1 \in_b_signal_reg[21]  (.D(n_156), .G(n_71), .Q(n_114));
   DLH_X1 \in_b_signal_reg[20]  (.D(n_155), .G(n_71), .Q(n_115));
   DLH_X1 \in_b_signal_reg[19]  (.D(n_154), .G(n_71), .Q(n_116));
   DLH_X1 \in_b_signal_reg[18]  (.D(n_153), .G(n_71), .Q(n_117));
   DLH_X1 \in_b_signal_reg[17]  (.D(n_152), .G(n_71), .Q(n_118));
   DLH_X1 \in_b_signal_reg[16]  (.D(n_151), .G(n_71), .Q(n_119));
   DLH_X1 \in_b_signal_reg[15]  (.D(n_150), .G(n_71), .Q(n_120));
   DLH_X1 \in_b_signal_reg[14]  (.D(n_149), .G(n_71), .Q(n_121));
   DLH_X1 \in_b_signal_reg[13]  (.D(n_148), .G(n_71), .Q(n_122));
   DLH_X1 \in_b_signal_reg[12]  (.D(n_147), .G(n_71), .Q(n_123));
   DLH_X1 \in_b_signal_reg[11]  (.D(n_146), .G(n_71), .Q(n_124));
   DLH_X1 \in_b_signal_reg[10]  (.D(n_145), .G(n_71), .Q(n_125));
   DLH_X1 \in_b_signal_reg[9]  (.D(n_144), .G(n_71), .Q(n_126));
   DLH_X1 \in_b_signal_reg[8]  (.D(n_143), .G(n_71), .Q(n_127));
   DLH_X1 \in_b_signal_reg[7]  (.D(n_142), .G(n_71), .Q(n_128));
   DLH_X1 \in_b_signal_reg[6]  (.D(n_141), .G(n_71), .Q(n_129));
   DLH_X1 \in_b_signal_reg[5]  (.D(n_140), .G(n_71), .Q(n_130));
   DLH_X1 \in_b_signal_reg[4]  (.D(n_139), .G(n_71), .Q(n_131));
   DLH_X1 \in_b_signal_reg[3]  (.D(n_138), .G(n_71), .Q(n_132));
   DLH_X1 \in_b_signal_reg[2]  (.D(n_137), .G(n_71), .Q(n_133));
   DLH_X1 \in_b_signal_reg[1]  (.D(n_136), .G(n_71), .Q(n_134));
   DLH_X1 \in_b_signal_reg[0]  (.D(in_b[0]), .G(n_71), .Q(n_135));
   datapath__0_6 i_9 (.plus({n_3, n_2, n_1, n_0, n_194, n_193, n_192, n_191, 
      n_190, n_189, n_188, n_187, n_186, n_185, n_184, n_183, n_182, n_181, 
      n_180, n_179, n_178, n_177, n_176, n_175, n_174, n_173, n_172, n_171, 
      n_170, n_169, n_168, n_167, n_166, n_165, n_164, n_163, n_162, n_161, 
      n_160, n_159, n_158, n_157, n_156, n_155, n_154, n_153, n_152, n_151, 
      n_150, n_149, n_148, n_147, n_146, n_145, n_144, n_143, n_142, n_141, 
      n_140, n_139, n_138, n_137, n_136, uc_0}), .in_b(in_b));
   INV_X1 i_0_0 (.A(rst), .ZN(n_71));
   AND2_X1 i_0_1 (.A1(n_71), .A2(n_6), .ZN(out_c[0]));
   AND2_X1 i_0_2 (.A1(n_71), .A2(F), .ZN(out_c[1]));
   AND2_X1 i_0_3 (.A1(n_71), .A2(F0), .ZN(out_c[2]));
   AND2_X1 i_0_4 (.A1(n_71), .A2(F1), .ZN(out_c[3]));
   AND2_X1 i_0_5 (.A1(n_71), .A2(F2), .ZN(out_c[4]));
   AND2_X1 i_0_6 (.A1(n_71), .A2(F3), .ZN(out_c[5]));
   AND2_X1 i_0_7 (.A1(n_71), .A2(F4), .ZN(out_c[6]));
   AND2_X1 i_0_8 (.A1(n_71), .A2(F5), .ZN(out_c[7]));
   AND2_X1 i_0_9 (.A1(n_71), .A2(F6), .ZN(out_c[8]));
   AND2_X1 i_0_10 (.A1(n_71), .A2(F7), .ZN(out_c[9]));
   AND2_X1 i_0_11 (.A1(n_71), .A2(F8), .ZN(out_c[10]));
   AND2_X1 i_0_12 (.A1(n_71), .A2(F9), .ZN(out_c[11]));
   AND2_X1 i_0_13 (.A1(n_71), .A2(F10), .ZN(out_c[12]));
   AND2_X1 i_0_14 (.A1(n_71), .A2(F11), .ZN(out_c[13]));
   AND2_X1 i_0_15 (.A1(n_71), .A2(F12), .ZN(out_c[14]));
   AND2_X1 i_0_16 (.A1(n_71), .A2(F13), .ZN(out_c[15]));
   AND2_X1 i_0_17 (.A1(n_71), .A2(F14), .ZN(out_c[16]));
   AND2_X1 i_0_18 (.A1(n_71), .A2(F15), .ZN(out_c[17]));
   AND2_X1 i_0_19 (.A1(n_71), .A2(F16), .ZN(out_c[18]));
   AND2_X1 i_0_20 (.A1(n_71), .A2(F17), .ZN(out_c[19]));
   AND2_X1 i_0_21 (.A1(n_71), .A2(F18), .ZN(out_c[20]));
   AND2_X1 i_0_22 (.A1(n_71), .A2(F19), .ZN(out_c[21]));
   AND2_X1 i_0_23 (.A1(n_71), .A2(F20), .ZN(out_c[22]));
   AND2_X1 i_0_24 (.A1(n_71), .A2(F21), .ZN(out_c[23]));
   AND2_X1 i_0_25 (.A1(n_71), .A2(F22), .ZN(out_c[24]));
   AND2_X1 i_0_26 (.A1(n_71), .A2(F23), .ZN(out_c[25]));
   AND2_X1 i_0_27 (.A1(n_71), .A2(F24), .ZN(out_c[26]));
   AND2_X1 i_0_28 (.A1(n_71), .A2(F25), .ZN(out_c[27]));
   AND2_X1 i_0_29 (.A1(n_71), .A2(F26), .ZN(out_c[28]));
   AND2_X1 i_0_30 (.A1(n_71), .A2(F27), .ZN(out_c[29]));
   AND2_X1 i_0_31 (.A1(n_71), .A2(F28), .ZN(out_c[30]));
   AND2_X1 i_0_32 (.A1(n_71), .A2(F29), .ZN(out_c[31]));
   AND2_X1 i_0_33 (.A1(n_71), .A2(F30), .ZN(out_c[32]));
   AND2_X1 i_0_34 (.A1(n_71), .A2(F31), .ZN(out_c[33]));
   AND2_X1 i_0_35 (.A1(n_71), .A2(F32), .ZN(out_c[34]));
   AND2_X1 i_0_36 (.A1(n_71), .A2(F33), .ZN(out_c[35]));
   AND2_X1 i_0_37 (.A1(n_71), .A2(F34), .ZN(out_c[36]));
   AND2_X1 i_0_38 (.A1(n_71), .A2(F35), .ZN(out_c[37]));
   AND2_X1 i_0_39 (.A1(n_71), .A2(F36), .ZN(out_c[38]));
   AND2_X1 i_0_40 (.A1(n_71), .A2(F37), .ZN(out_c[39]));
   AND2_X1 i_0_41 (.A1(n_71), .A2(F38), .ZN(out_c[40]));
   AND2_X1 i_0_42 (.A1(n_71), .A2(F39), .ZN(out_c[41]));
   AND2_X1 i_0_43 (.A1(n_71), .A2(F40), .ZN(out_c[42]));
   AND2_X1 i_0_44 (.A1(n_71), .A2(F41), .ZN(out_c[43]));
   AND2_X1 i_0_45 (.A1(n_71), .A2(F42), .ZN(out_c[44]));
   AND2_X1 i_0_46 (.A1(n_71), .A2(F43), .ZN(out_c[45]));
   AND2_X1 i_0_47 (.A1(n_71), .A2(F44), .ZN(out_c[46]));
   AND2_X1 i_0_48 (.A1(n_71), .A2(F45), .ZN(out_c[47]));
   AND2_X1 i_0_49 (.A1(n_71), .A2(F46), .ZN(out_c[48]));
   AND2_X1 i_0_50 (.A1(n_71), .A2(F47), .ZN(out_c[49]));
   AND2_X1 i_0_51 (.A1(n_71), .A2(F48), .ZN(out_c[50]));
   AND2_X1 i_0_52 (.A1(n_71), .A2(F49), .ZN(out_c[51]));
   AND2_X1 i_0_53 (.A1(n_71), .A2(F50), .ZN(out_c[52]));
   AND2_X1 i_0_54 (.A1(n_71), .A2(F51), .ZN(out_c[53]));
   AND2_X1 i_0_55 (.A1(n_71), .A2(F52), .ZN(out_c[54]));
   AND2_X1 i_0_56 (.A1(n_71), .A2(F53), .ZN(out_c[55]));
   AND2_X1 i_0_57 (.A1(n_71), .A2(F54), .ZN(out_c[56]));
   AND2_X1 i_0_58 (.A1(n_71), .A2(F55), .ZN(out_c[57]));
   AND2_X1 i_0_59 (.A1(n_71), .A2(F56), .ZN(out_c[58]));
   AND2_X1 i_0_60 (.A1(n_71), .A2(F57), .ZN(out_c[59]));
   AND2_X1 i_0_61 (.A1(n_71), .A2(F58), .ZN(out_c[60]));
   AND2_X1 i_0_62 (.A1(n_71), .A2(F59), .ZN(out_c[61]));
   AND2_X1 i_0_63 (.A1(n_71), .A2(n_5), .ZN(out_c[62]));
   AND2_X1 i_0_64 (.A1(n_71), .A2(n_4), .ZN(out_c[63]));
endmodule

module datapath__0_143(in_b, p_0);
   input [63:0]in_b;
   output [63:0]p_0;

   XOR2_X1 i_0 (.A(in_b[1]), .B(in_b[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_61), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(in_b[2]), .B1(in_b[1]), .B2(in_b[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(in_b[3]), .B(n_61), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(in_b[4]), .B(n_60), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(in_b[5]), .B(n_59), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_58), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(in_b[6]), .B1(n_59), .B2(in_b[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(in_b[7]), .B(n_58), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(in_b[8]), .B(n_57), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_56), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(in_b[9]), .B1(n_57), .B2(in_b[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(in_b[10]), .B(n_56), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(in_b[11]), .B(n_55), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(in_b[12]), .B(n_54), .Z(p_0[12]));
   XNOR2_X1 i_15 (.A(in_b[13]), .B(n_53), .ZN(p_0[13]));
   XOR2_X1 i_16 (.A(in_b[14]), .B(n_52), .Z(p_0[14]));
   AND2_X1 i_17 (.A1(n_51), .A2(n_3), .ZN(p_0[15]));
   OAI21_X1 i_18 (.A(in_b[15]), .B1(n_52), .B2(in_b[14]), .ZN(n_3));
   XOR2_X1 i_19 (.A(in_b[16]), .B(n_51), .Z(p_0[16]));
   XOR2_X1 i_20 (.A(in_b[17]), .B(n_50), .Z(p_0[17]));
   XOR2_X1 i_21 (.A(in_b[18]), .B(n_49), .Z(p_0[18]));
   XNOR2_X1 i_22 (.A(in_b[19]), .B(n_48), .ZN(p_0[19]));
   XNOR2_X1 i_23 (.A(in_b[20]), .B(n_47), .ZN(p_0[20]));
   XNOR2_X1 i_24 (.A(in_b[21]), .B(n_46), .ZN(p_0[21]));
   XOR2_X1 i_25 (.A(in_b[22]), .B(n_45), .Z(p_0[22]));
   XOR2_X1 i_26 (.A(in_b[23]), .B(n_44), .Z(p_0[23]));
   XNOR2_X1 i_27 (.A(in_b[24]), .B(n_43), .ZN(p_0[24]));
   XNOR2_X1 i_28 (.A(in_b[25]), .B(n_42), .ZN(p_0[25]));
   XNOR2_X1 i_29 (.A(in_b[26]), .B(n_41), .ZN(p_0[26]));
   XOR2_X1 i_30 (.A(in_b[27]), .B(n_40), .Z(p_0[27]));
   XOR2_X1 i_31 (.A(in_b[28]), .B(n_39), .Z(p_0[28]));
   XNOR2_X1 i_32 (.A(in_b[29]), .B(n_38), .ZN(p_0[29]));
   XNOR2_X1 i_33 (.A(in_b[30]), .B(n_37), .ZN(p_0[30]));
   XNOR2_X1 i_34 (.A(in_b[31]), .B(n_36), .ZN(p_0[31]));
   XOR2_X1 i_35 (.A(in_b[32]), .B(n_35), .Z(p_0[32]));
   XOR2_X1 i_36 (.A(in_b[33]), .B(n_34), .Z(p_0[33]));
   XNOR2_X1 i_37 (.A(in_b[34]), .B(n_33), .ZN(p_0[34]));
   XNOR2_X1 i_38 (.A(in_b[35]), .B(n_32), .ZN(p_0[35]));
   XNOR2_X1 i_39 (.A(in_b[36]), .B(n_31), .ZN(p_0[36]));
   XOR2_X1 i_40 (.A(in_b[37]), .B(n_30), .Z(p_0[37]));
   XOR2_X1 i_41 (.A(in_b[38]), .B(n_29), .Z(p_0[38]));
   XNOR2_X1 i_42 (.A(in_b[39]), .B(n_28), .ZN(p_0[39]));
   XNOR2_X1 i_43 (.A(in_b[40]), .B(n_27), .ZN(p_0[40]));
   XOR2_X1 i_44 (.A(in_b[41]), .B(n_26), .Z(p_0[41]));
   XNOR2_X1 i_45 (.A(in_b[42]), .B(n_25), .ZN(p_0[42]));
   XOR2_X1 i_46 (.A(in_b[43]), .B(n_24), .Z(p_0[43]));
   AND2_X1 i_47 (.A1(n_23), .A2(n_4), .ZN(p_0[44]));
   OAI21_X1 i_48 (.A(in_b[44]), .B1(n_24), .B2(in_b[43]), .ZN(n_4));
   XOR2_X1 i_49 (.A(in_b[45]), .B(n_23), .Z(p_0[45]));
   XOR2_X1 i_50 (.A(in_b[46]), .B(n_22), .Z(p_0[46]));
   XOR2_X1 i_51 (.A(in_b[47]), .B(n_21), .Z(p_0[47]));
   XOR2_X1 i_52 (.A(in_b[48]), .B(n_20), .Z(p_0[48]));
   XNOR2_X1 i_53 (.A(in_b[49]), .B(n_19), .ZN(p_0[49]));
   XNOR2_X1 i_54 (.A(in_b[50]), .B(n_18), .ZN(p_0[50]));
   XNOR2_X1 i_55 (.A(in_b[51]), .B(n_17), .ZN(p_0[51]));
   XOR2_X1 i_56 (.A(in_b[52]), .B(n_16), .Z(p_0[52]));
   XNOR2_X1 i_57 (.A(in_b[53]), .B(n_15), .ZN(p_0[53]));
   XNOR2_X1 i_58 (.A(in_b[54]), .B(n_14), .ZN(p_0[54]));
   XNOR2_X1 i_59 (.A(in_b[55]), .B(n_13), .ZN(p_0[55]));
   XOR2_X1 i_60 (.A(in_b[56]), .B(n_12), .Z(p_0[56]));
   AND2_X1 i_61 (.A1(n_11), .A2(n_5), .ZN(p_0[57]));
   OAI21_X1 i_62 (.A(in_b[57]), .B1(n_12), .B2(in_b[56]), .ZN(n_5));
   XOR2_X1 i_63 (.A(in_b[58]), .B(n_11), .Z(p_0[58]));
   XNOR2_X1 i_64 (.A(in_b[59]), .B(n_10), .ZN(p_0[59]));
   XNOR2_X1 i_65 (.A(in_b[60]), .B(n_9), .ZN(p_0[60]));
   XOR2_X1 i_66 (.A(in_b[61]), .B(n_8), .Z(p_0[61]));
   XNOR2_X1 i_67 (.A(in_b[62]), .B(n_7), .ZN(p_0[62]));
   XNOR2_X1 i_68 (.A(in_b[63]), .B(n_6), .ZN(p_0[63]));
   NOR3_X1 i_69 (.A1(n_8), .A2(in_b[61]), .A3(in_b[62]), .ZN(n_6));
   NOR2_X1 i_70 (.A1(n_8), .A2(in_b[61]), .ZN(n_7));
   NAND2_X1 i_71 (.A1(n_9), .A2(n_72), .ZN(n_8));
   NOR3_X1 i_72 (.A1(n_11), .A2(in_b[58]), .A3(in_b[59]), .ZN(n_9));
   NOR2_X1 i_73 (.A1(n_11), .A2(in_b[58]), .ZN(n_10));
   OR3_X1 i_74 (.A1(n_12), .A2(in_b[56]), .A3(in_b[57]), .ZN(n_11));
   NAND2_X1 i_75 (.A1(n_13), .A2(n_71), .ZN(n_12));
   NOR4_X1 i_76 (.A1(n_16), .A2(in_b[52]), .A3(in_b[53]), .A4(in_b[54]), 
      .ZN(n_13));
   NOR3_X1 i_77 (.A1(n_16), .A2(in_b[52]), .A3(in_b[53]), .ZN(n_14));
   NOR2_X1 i_78 (.A1(n_16), .A2(in_b[52]), .ZN(n_15));
   NAND2_X1 i_79 (.A1(n_17), .A2(n_70), .ZN(n_16));
   NOR4_X1 i_80 (.A1(n_20), .A2(in_b[48]), .A3(in_b[49]), .A4(in_b[50]), 
      .ZN(n_17));
   NOR3_X1 i_81 (.A1(n_20), .A2(in_b[48]), .A3(in_b[49]), .ZN(n_18));
   NOR2_X1 i_82 (.A1(n_20), .A2(in_b[48]), .ZN(n_19));
   OR2_X1 i_83 (.A1(n_21), .A2(in_b[47]), .ZN(n_20));
   OR2_X1 i_84 (.A1(n_22), .A2(in_b[46]), .ZN(n_21));
   OR2_X1 i_85 (.A1(n_23), .A2(in_b[45]), .ZN(n_22));
   OR3_X1 i_86 (.A1(n_24), .A2(in_b[43]), .A3(in_b[44]), .ZN(n_23));
   NAND2_X1 i_87 (.A1(n_25), .A2(n_69), .ZN(n_24));
   NOR2_X1 i_88 (.A1(n_26), .A2(in_b[41]), .ZN(n_25));
   NAND2_X1 i_89 (.A1(n_27), .A2(n_68), .ZN(n_26));
   NOR3_X1 i_90 (.A1(n_29), .A2(in_b[38]), .A3(in_b[39]), .ZN(n_27));
   NOR2_X1 i_91 (.A1(n_29), .A2(in_b[38]), .ZN(n_28));
   OR2_X1 i_92 (.A1(n_30), .A2(in_b[37]), .ZN(n_29));
   NAND2_X1 i_93 (.A1(n_31), .A2(n_67), .ZN(n_30));
   NOR4_X1 i_94 (.A1(n_34), .A2(in_b[33]), .A3(in_b[34]), .A4(in_b[35]), 
      .ZN(n_31));
   NOR3_X1 i_95 (.A1(n_34), .A2(in_b[33]), .A3(in_b[34]), .ZN(n_32));
   NOR2_X1 i_96 (.A1(n_34), .A2(in_b[33]), .ZN(n_33));
   OR2_X1 i_97 (.A1(n_35), .A2(in_b[32]), .ZN(n_34));
   NAND2_X1 i_98 (.A1(n_36), .A2(n_66), .ZN(n_35));
   NOR4_X1 i_99 (.A1(n_39), .A2(in_b[28]), .A3(in_b[29]), .A4(in_b[30]), 
      .ZN(n_36));
   NOR3_X1 i_100 (.A1(n_39), .A2(in_b[28]), .A3(in_b[29]), .ZN(n_37));
   NOR2_X1 i_101 (.A1(n_39), .A2(in_b[28]), .ZN(n_38));
   OR2_X1 i_102 (.A1(n_40), .A2(in_b[27]), .ZN(n_39));
   NAND2_X1 i_103 (.A1(n_41), .A2(n_65), .ZN(n_40));
   NOR4_X1 i_104 (.A1(n_44), .A2(in_b[23]), .A3(in_b[24]), .A4(in_b[25]), 
      .ZN(n_41));
   NOR3_X1 i_105 (.A1(n_44), .A2(in_b[23]), .A3(in_b[24]), .ZN(n_42));
   NOR2_X1 i_106 (.A1(n_44), .A2(in_b[23]), .ZN(n_43));
   OR2_X1 i_107 (.A1(n_45), .A2(in_b[22]), .ZN(n_44));
   NAND2_X1 i_108 (.A1(n_46), .A2(n_64), .ZN(n_45));
   NOR4_X1 i_109 (.A1(n_49), .A2(in_b[18]), .A3(in_b[19]), .A4(in_b[20]), 
      .ZN(n_46));
   NOR3_X1 i_110 (.A1(n_49), .A2(in_b[18]), .A3(in_b[19]), .ZN(n_47));
   NOR2_X1 i_111 (.A1(n_49), .A2(in_b[18]), .ZN(n_48));
   OR2_X1 i_112 (.A1(n_50), .A2(in_b[17]), .ZN(n_49));
   OR2_X1 i_113 (.A1(n_51), .A2(in_b[16]), .ZN(n_50));
   OR3_X1 i_114 (.A1(n_52), .A2(in_b[14]), .A3(in_b[15]), .ZN(n_51));
   NAND2_X1 i_115 (.A1(n_53), .A2(n_63), .ZN(n_52));
   NOR2_X1 i_116 (.A1(n_54), .A2(in_b[12]), .ZN(n_53));
   NAND2_X1 i_117 (.A1(n_55), .A2(n_62), .ZN(n_54));
   NOR2_X1 i_118 (.A1(n_56), .A2(in_b[10]), .ZN(n_55));
   OR3_X1 i_119 (.A1(n_57), .A2(in_b[8]), .A3(in_b[9]), .ZN(n_56));
   OR2_X1 i_120 (.A1(n_58), .A2(in_b[7]), .ZN(n_57));
   OR3_X1 i_121 (.A1(n_59), .A2(in_b[5]), .A3(in_b[6]), .ZN(n_58));
   OR2_X1 i_122 (.A1(n_60), .A2(in_b[4]), .ZN(n_59));
   OR2_X1 i_123 (.A1(n_61), .A2(in_b[3]), .ZN(n_60));
   OR3_X1 i_124 (.A1(in_b[2]), .A2(in_b[1]), .A3(in_b[0]), .ZN(n_61));
   INV_X1 i_125 (.A(in_b[11]), .ZN(n_62));
   INV_X1 i_126 (.A(in_b[13]), .ZN(n_63));
   INV_X1 i_127 (.A(in_b[21]), .ZN(n_64));
   INV_X1 i_128 (.A(in_b[26]), .ZN(n_65));
   INV_X1 i_129 (.A(in_b[31]), .ZN(n_66));
   INV_X1 i_130 (.A(in_b[36]), .ZN(n_67));
   INV_X1 i_131 (.A(in_b[40]), .ZN(n_68));
   INV_X1 i_132 (.A(in_b[42]), .ZN(n_69));
   INV_X1 i_133 (.A(in_b[51]), .ZN(n_70));
   INV_X1 i_134 (.A(in_b[55]), .ZN(n_71));
   INV_X1 i_135 (.A(in_b[60]), .ZN(n_72));
endmodule

module datapath__0_146(in_a, p_0);
   input [63:0]in_a;
   output [63:0]p_0;

   XOR2_X1 i_0 (.A(in_a[1]), .B(in_a[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_54), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(in_a[2]), .B1(in_a[1]), .B2(in_a[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(in_a[3]), .B(n_54), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(in_a[4]), .B(n_53), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(in_a[5]), .B(n_52), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_51), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(in_a[6]), .B1(n_52), .B2(in_a[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(in_a[7]), .B(n_51), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(in_a[8]), .B(n_50), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_49), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(in_a[9]), .B1(n_50), .B2(in_a[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(in_a[10]), .B(n_49), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(in_a[11]), .B(n_48), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(in_a[12]), .B(n_47), .Z(p_0[12]));
   XNOR2_X1 i_15 (.A(in_a[13]), .B(n_46), .ZN(p_0[13]));
   XOR2_X1 i_16 (.A(in_a[14]), .B(n_45), .Z(p_0[14]));
   AND2_X1 i_17 (.A1(n_44), .A2(n_3), .ZN(p_0[15]));
   OAI21_X1 i_18 (.A(in_a[15]), .B1(n_45), .B2(in_a[14]), .ZN(n_3));
   XOR2_X1 i_19 (.A(in_a[16]), .B(n_44), .Z(p_0[16]));
   XOR2_X1 i_20 (.A(in_a[17]), .B(n_43), .Z(p_0[17]));
   XOR2_X1 i_21 (.A(in_a[18]), .B(n_42), .Z(p_0[18]));
   XOR2_X1 i_22 (.A(in_a[19]), .B(n_41), .Z(p_0[19]));
   XNOR2_X1 i_23 (.A(in_a[20]), .B(n_40), .ZN(p_0[20]));
   XNOR2_X1 i_24 (.A(in_a[21]), .B(n_39), .ZN(p_0[21]));
   XNOR2_X1 i_25 (.A(in_a[22]), .B(n_38), .ZN(p_0[22]));
   XOR2_X1 i_26 (.A(in_a[23]), .B(n_37), .Z(p_0[23]));
   XNOR2_X1 i_27 (.A(in_a[24]), .B(n_36), .ZN(p_0[24]));
   XNOR2_X1 i_28 (.A(in_a[25]), .B(n_35), .ZN(p_0[25]));
   XNOR2_X1 i_29 (.A(in_a[26]), .B(n_34), .ZN(p_0[26]));
   XOR2_X1 i_30 (.A(in_a[27]), .B(n_33), .Z(p_0[27]));
   XOR2_X1 i_31 (.A(in_a[28]), .B(n_32), .Z(p_0[28]));
   XNOR2_X1 i_32 (.A(in_a[29]), .B(n_31), .ZN(p_0[29]));
   XNOR2_X1 i_33 (.A(in_a[30]), .B(n_30), .ZN(p_0[30]));
   XNOR2_X1 i_34 (.A(in_a[31]), .B(n_29), .ZN(p_0[31]));
   XOR2_X1 i_35 (.A(in_a[32]), .B(n_28), .Z(p_0[32]));
   XOR2_X1 i_36 (.A(in_a[33]), .B(n_27), .Z(p_0[33]));
   XNOR2_X1 i_37 (.A(in_a[34]), .B(n_26), .ZN(p_0[34]));
   XNOR2_X1 i_38 (.A(in_a[35]), .B(n_25), .ZN(p_0[35]));
   XOR2_X1 i_39 (.A(in_a[36]), .B(n_24), .Z(p_0[36]));
   XOR2_X1 i_40 (.A(in_a[37]), .B(n_23), .Z(p_0[37]));
   XOR2_X1 i_41 (.A(in_a[38]), .B(n_22), .Z(p_0[38]));
   XNOR2_X1 i_42 (.A(in_a[39]), .B(n_21), .ZN(p_0[39]));
   XNOR2_X1 i_43 (.A(in_a[40]), .B(n_20), .ZN(p_0[40]));
   XNOR2_X1 i_44 (.A(in_a[41]), .B(n_19), .ZN(p_0[41]));
   XOR2_X1 i_45 (.A(in_a[42]), .B(n_18), .Z(p_0[42]));
   XOR2_X1 i_46 (.A(in_a[43]), .B(n_17), .Z(p_0[43]));
   XNOR2_X1 i_47 (.A(in_a[44]), .B(n_16), .ZN(p_0[44]));
   XNOR2_X1 i_48 (.A(in_a[45]), .B(n_15), .ZN(p_0[45]));
   XNOR2_X1 i_49 (.A(in_a[46]), .B(n_14), .ZN(p_0[46]));
   XOR2_X1 i_50 (.A(in_a[47]), .B(n_13), .Z(p_0[47]));
   XOR2_X1 i_51 (.A(in_a[48]), .B(n_12), .Z(p_0[48]));
   XNOR2_X1 i_52 (.A(in_a[49]), .B(n_11), .ZN(p_0[49]));
   XNOR2_X1 i_53 (.A(in_a[50]), .B(n_10), .ZN(p_0[50]));
   XOR2_X1 i_54 (.A(in_a[51]), .B(n_9), .Z(p_0[51]));
   AND2_X1 i_55 (.A1(n_8), .A2(n_4), .ZN(p_0[52]));
   OAI21_X1 i_56 (.A(in_a[52]), .B1(n_9), .B2(in_a[51]), .ZN(n_4));
   XOR2_X1 i_57 (.A(in_a[53]), .B(n_8), .Z(p_0[53]));
   XNOR2_X1 i_58 (.A(in_a[54]), .B(n_7), .ZN(p_0[54]));
   XNOR2_X1 i_59 (.A(in_a[55]), .B(n_6), .ZN(p_0[55]));
   XNOR2_X1 i_60 (.A(in_a[56]), .B(n_5), .ZN(p_0[56]));
   NOR4_X1 i_61 (.A1(n_8), .A2(in_a[53]), .A3(in_a[54]), .A4(in_a[55]), .ZN(n_5));
   NOR3_X1 i_62 (.A1(n_8), .A2(in_a[53]), .A3(in_a[54]), .ZN(n_6));
   NOR2_X1 i_63 (.A1(n_8), .A2(in_a[53]), .ZN(n_7));
   OR3_X1 i_64 (.A1(n_9), .A2(in_a[51]), .A3(in_a[52]), .ZN(n_8));
   NAND2_X1 i_65 (.A1(n_10), .A2(n_63), .ZN(n_9));
   NOR3_X1 i_66 (.A1(n_12), .A2(in_a[48]), .A3(in_a[49]), .ZN(n_10));
   NOR2_X1 i_67 (.A1(n_12), .A2(in_a[48]), .ZN(n_11));
   OR2_X1 i_68 (.A1(n_13), .A2(in_a[47]), .ZN(n_12));
   NAND2_X1 i_69 (.A1(n_14), .A2(n_62), .ZN(n_13));
   NOR4_X1 i_70 (.A1(n_17), .A2(in_a[43]), .A3(in_a[44]), .A4(in_a[45]), 
      .ZN(n_14));
   NOR3_X1 i_71 (.A1(n_17), .A2(in_a[43]), .A3(in_a[44]), .ZN(n_15));
   NOR2_X1 i_72 (.A1(n_17), .A2(in_a[43]), .ZN(n_16));
   OR2_X1 i_73 (.A1(n_18), .A2(in_a[42]), .ZN(n_17));
   NAND2_X1 i_74 (.A1(n_19), .A2(n_61), .ZN(n_18));
   NOR4_X1 i_75 (.A1(n_22), .A2(in_a[38]), .A3(in_a[39]), .A4(in_a[40]), 
      .ZN(n_19));
   NOR3_X1 i_76 (.A1(n_22), .A2(in_a[38]), .A3(in_a[39]), .ZN(n_20));
   NOR2_X1 i_77 (.A1(n_22), .A2(in_a[38]), .ZN(n_21));
   OR2_X1 i_78 (.A1(n_23), .A2(in_a[37]), .ZN(n_22));
   OR2_X1 i_79 (.A1(n_24), .A2(in_a[36]), .ZN(n_23));
   NAND2_X1 i_80 (.A1(n_25), .A2(n_60), .ZN(n_24));
   NOR3_X1 i_81 (.A1(n_27), .A2(in_a[33]), .A3(in_a[34]), .ZN(n_25));
   NOR2_X1 i_82 (.A1(n_27), .A2(in_a[33]), .ZN(n_26));
   OR2_X1 i_83 (.A1(n_28), .A2(in_a[32]), .ZN(n_27));
   NAND2_X1 i_84 (.A1(n_29), .A2(n_59), .ZN(n_28));
   NOR4_X1 i_85 (.A1(n_32), .A2(in_a[28]), .A3(in_a[29]), .A4(in_a[30]), 
      .ZN(n_29));
   NOR3_X1 i_86 (.A1(n_32), .A2(in_a[28]), .A3(in_a[29]), .ZN(n_30));
   NOR2_X1 i_87 (.A1(n_32), .A2(in_a[28]), .ZN(n_31));
   OR2_X1 i_88 (.A1(n_33), .A2(in_a[27]), .ZN(n_32));
   NAND2_X1 i_89 (.A1(n_34), .A2(n_58), .ZN(n_33));
   NOR4_X1 i_90 (.A1(n_37), .A2(in_a[23]), .A3(in_a[24]), .A4(in_a[25]), 
      .ZN(n_34));
   NOR3_X1 i_91 (.A1(n_37), .A2(in_a[23]), .A3(in_a[24]), .ZN(n_35));
   NOR2_X1 i_92 (.A1(n_37), .A2(in_a[23]), .ZN(n_36));
   NAND2_X1 i_93 (.A1(n_38), .A2(n_57), .ZN(n_37));
   NOR4_X1 i_94 (.A1(n_41), .A2(in_a[19]), .A3(in_a[20]), .A4(in_a[21]), 
      .ZN(n_38));
   NOR3_X1 i_95 (.A1(n_41), .A2(in_a[19]), .A3(in_a[20]), .ZN(n_39));
   NOR2_X1 i_96 (.A1(n_41), .A2(in_a[19]), .ZN(n_40));
   OR2_X1 i_97 (.A1(n_42), .A2(in_a[18]), .ZN(n_41));
   OR2_X1 i_98 (.A1(n_43), .A2(in_a[17]), .ZN(n_42));
   OR2_X1 i_99 (.A1(n_44), .A2(in_a[16]), .ZN(n_43));
   OR3_X1 i_100 (.A1(n_45), .A2(in_a[14]), .A3(in_a[15]), .ZN(n_44));
   NAND2_X1 i_101 (.A1(n_46), .A2(n_56), .ZN(n_45));
   NOR2_X1 i_102 (.A1(n_47), .A2(in_a[12]), .ZN(n_46));
   NAND2_X1 i_103 (.A1(n_48), .A2(n_55), .ZN(n_47));
   NOR2_X1 i_104 (.A1(n_49), .A2(in_a[10]), .ZN(n_48));
   OR3_X1 i_105 (.A1(n_50), .A2(in_a[8]), .A3(in_a[9]), .ZN(n_49));
   OR2_X1 i_106 (.A1(n_51), .A2(in_a[7]), .ZN(n_50));
   OR3_X1 i_107 (.A1(n_52), .A2(in_a[5]), .A3(in_a[6]), .ZN(n_51));
   OR2_X1 i_108 (.A1(n_53), .A2(in_a[4]), .ZN(n_52));
   OR2_X1 i_109 (.A1(n_54), .A2(in_a[3]), .ZN(n_53));
   OR3_X1 i_110 (.A1(in_a[2]), .A2(in_a[1]), .A3(in_a[0]), .ZN(n_54));
   INV_X1 i_111 (.A(in_a[11]), .ZN(n_55));
   INV_X1 i_112 (.A(in_a[13]), .ZN(n_56));
   INV_X1 i_113 (.A(in_a[22]), .ZN(n_57));
   INV_X1 i_114 (.A(in_a[26]), .ZN(n_58));
   INV_X1 i_115 (.A(in_a[31]), .ZN(n_59));
   INV_X1 i_116 (.A(in_a[35]), .ZN(n_60));
   INV_X1 i_117 (.A(in_a[41]), .ZN(n_61));
   INV_X1 i_118 (.A(in_a[46]), .ZN(n_62));
   INV_X1 i_119 (.A(in_a[50]), .ZN(n_63));
endmodule

module datapath__0_43(i, p_0);
   input [31:0]i;
   output [31:0]p_0;

   HA_X1 i_0 (.A(i[1]), .B(i[0]), .CO(n_0), .S(p_0[1]));
   HA_X1 i_1 (.A(i[2]), .B(n_0), .CO(n_1), .S(p_0[2]));
   HA_X1 i_2 (.A(i[3]), .B(n_1), .CO(n_2), .S(p_0[3]));
   HA_X1 i_3 (.A(i[4]), .B(n_2), .CO(n_3), .S(p_0[4]));
   HA_X1 i_4 (.A(i[5]), .B(n_3), .CO(n_4), .S(p_0[5]));
   HA_X1 i_5 (.A(i[6]), .B(n_4), .CO(n_5), .S(p_0[6]));
   HA_X1 i_6 (.A(i[7]), .B(n_5), .CO(n_6), .S(p_0[7]));
   HA_X1 i_7 (.A(i[8]), .B(n_6), .CO(n_7), .S(p_0[8]));
   HA_X1 i_8 (.A(i[9]), .B(n_7), .CO(n_8), .S(p_0[9]));
   HA_X1 i_9 (.A(i[10]), .B(n_8), .CO(n_9), .S(p_0[10]));
   HA_X1 i_11 (.A(i[11]), .B(n_9), .CO(n_10), .S(p_0[11]));
   HA_X1 i_12 (.A(i[12]), .B(n_10), .CO(n_11), .S(p_0[12]));
   HA_X1 i_13 (.A(i[13]), .B(n_11), .CO(n_12), .S(p_0[13]));
   HA_X1 i_14 (.A(i[14]), .B(n_12), .CO(n_13), .S(p_0[14]));
   HA_X1 i_15 (.A(i[15]), .B(n_13), .CO(n_14), .S(p_0[15]));
   HA_X1 i_16 (.A(i[16]), .B(n_14), .CO(n_15), .S(p_0[16]));
   HA_X1 i_17 (.A(i[17]), .B(n_15), .CO(n_16), .S(p_0[17]));
   HA_X1 i_18 (.A(i[18]), .B(n_16), .CO(n_17), .S(p_0[18]));
   HA_X1 i_19 (.A(i[19]), .B(n_17), .CO(n_18), .S(p_0[19]));
   HA_X1 i_10 (.A(i[20]), .B(n_18), .CO(n_19), .S(p_0[20]));
   HA_X1 i_20 (.A(i[21]), .B(n_19), .CO(n_20), .S(p_0[21]));
   HA_X1 i_21 (.A(i[22]), .B(n_20), .CO(n_21), .S(p_0[22]));
   HA_X1 i_22 (.A(i[23]), .B(n_21), .CO(n_22), .S(p_0[23]));
   HA_X1 i_23 (.A(i[24]), .B(n_22), .CO(n_23), .S(p_0[24]));
   HA_X1 i_24 (.A(i[25]), .B(n_23), .CO(n_24), .S(p_0[25]));
   HA_X1 i_25 (.A(i[26]), .B(n_24), .CO(n_25), .S(p_0[26]));
   HA_X1 i_26 (.A(i[27]), .B(n_25), .CO(n_26), .S(p_0[27]));
   HA_X1 i_27 (.A(i[28]), .B(n_26), .CO(n_27), .S(p_0[28]));
   HA_X1 i_28 (.A(i[29]), .B(n_27), .CO(n_28), .S(p_0[29]));
   HA_X1 i_29 (.A(i[30]), .B(n_28), .CO(n_29), .S(p_0[30]));
   XOR2_X1 i_30 (.A(i[31]), .B(n_29), .Z(p_0[31]));
   INV_X1 i_31 (.A(i[0]), .ZN(p_0[0]));
endmodule

module datapath__0_162(plus, quotient);
   output [63:0]plus;
   input [63:0]quotient;

   XOR2_X1 i_0 (.A(quotient[1]), .B(quotient[0]), .Z(plus[1]));
   AND2_X1 i_1 (.A1(n_61), .A2(n_0), .ZN(plus[2]));
   OAI21_X1 i_2 (.A(quotient[2]), .B1(quotient[1]), .B2(quotient[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(quotient[3]), .B(n_61), .Z(plus[3]));
   XOR2_X1 i_4 (.A(quotient[4]), .B(n_60), .Z(plus[4]));
   XOR2_X1 i_5 (.A(quotient[5]), .B(n_59), .Z(plus[5]));
   AND2_X1 i_6 (.A1(n_58), .A2(n_1), .ZN(plus[6]));
   OAI21_X1 i_7 (.A(quotient[6]), .B1(n_59), .B2(quotient[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(quotient[7]), .B(n_58), .Z(plus[7]));
   XOR2_X1 i_9 (.A(quotient[8]), .B(n_57), .Z(plus[8]));
   AND2_X1 i_10 (.A1(n_56), .A2(n_2), .ZN(plus[9]));
   OAI21_X1 i_11 (.A(quotient[9]), .B1(n_57), .B2(quotient[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(quotient[10]), .B(n_56), .Z(plus[10]));
   XNOR2_X1 i_13 (.A(quotient[11]), .B(n_55), .ZN(plus[11]));
   XOR2_X1 i_14 (.A(quotient[12]), .B(n_54), .Z(plus[12]));
   XNOR2_X1 i_15 (.A(quotient[13]), .B(n_53), .ZN(plus[13]));
   XOR2_X1 i_16 (.A(quotient[14]), .B(n_52), .Z(plus[14]));
   AND2_X1 i_17 (.A1(n_51), .A2(n_3), .ZN(plus[15]));
   OAI21_X1 i_18 (.A(quotient[15]), .B1(n_52), .B2(quotient[14]), .ZN(n_3));
   XOR2_X1 i_19 (.A(quotient[16]), .B(n_51), .Z(plus[16]));
   XOR2_X1 i_20 (.A(quotient[17]), .B(n_50), .Z(plus[17]));
   XOR2_X1 i_21 (.A(quotient[18]), .B(n_49), .Z(plus[18]));
   XNOR2_X1 i_22 (.A(quotient[19]), .B(n_48), .ZN(plus[19]));
   XNOR2_X1 i_23 (.A(quotient[20]), .B(n_47), .ZN(plus[20]));
   XNOR2_X1 i_24 (.A(quotient[21]), .B(n_46), .ZN(plus[21]));
   XOR2_X1 i_25 (.A(quotient[22]), .B(n_45), .Z(plus[22]));
   XOR2_X1 i_26 (.A(quotient[23]), .B(n_44), .Z(plus[23]));
   XNOR2_X1 i_27 (.A(quotient[24]), .B(n_43), .ZN(plus[24]));
   XNOR2_X1 i_28 (.A(quotient[25]), .B(n_42), .ZN(plus[25]));
   XNOR2_X1 i_29 (.A(quotient[26]), .B(n_41), .ZN(plus[26]));
   XOR2_X1 i_30 (.A(quotient[27]), .B(n_40), .Z(plus[27]));
   XOR2_X1 i_31 (.A(quotient[28]), .B(n_39), .Z(plus[28]));
   XNOR2_X1 i_32 (.A(quotient[29]), .B(n_38), .ZN(plus[29]));
   XNOR2_X1 i_33 (.A(quotient[30]), .B(n_37), .ZN(plus[30]));
   XNOR2_X1 i_34 (.A(quotient[31]), .B(n_36), .ZN(plus[31]));
   XOR2_X1 i_35 (.A(quotient[32]), .B(n_35), .Z(plus[32]));
   XOR2_X1 i_36 (.A(quotient[33]), .B(n_34), .Z(plus[33]));
   XNOR2_X1 i_37 (.A(quotient[34]), .B(n_33), .ZN(plus[34]));
   XNOR2_X1 i_38 (.A(quotient[35]), .B(n_32), .ZN(plus[35]));
   XNOR2_X1 i_39 (.A(quotient[36]), .B(n_31), .ZN(plus[36]));
   XOR2_X1 i_40 (.A(quotient[37]), .B(n_30), .Z(plus[37]));
   XOR2_X1 i_41 (.A(quotient[38]), .B(n_29), .Z(plus[38]));
   XNOR2_X1 i_42 (.A(quotient[39]), .B(n_28), .ZN(plus[39]));
   XNOR2_X1 i_43 (.A(quotient[40]), .B(n_27), .ZN(plus[40]));
   XOR2_X1 i_44 (.A(quotient[41]), .B(n_26), .Z(plus[41]));
   XNOR2_X1 i_45 (.A(quotient[42]), .B(n_25), .ZN(plus[42]));
   XOR2_X1 i_46 (.A(quotient[43]), .B(n_24), .Z(plus[43]));
   AND2_X1 i_47 (.A1(n_23), .A2(n_4), .ZN(plus[44]));
   OAI21_X1 i_48 (.A(quotient[44]), .B1(n_24), .B2(quotient[43]), .ZN(n_4));
   XOR2_X1 i_49 (.A(quotient[45]), .B(n_23), .Z(plus[45]));
   XOR2_X1 i_50 (.A(quotient[46]), .B(n_22), .Z(plus[46]));
   XOR2_X1 i_51 (.A(quotient[47]), .B(n_21), .Z(plus[47]));
   XOR2_X1 i_52 (.A(quotient[48]), .B(n_20), .Z(plus[48]));
   XNOR2_X1 i_53 (.A(quotient[49]), .B(n_19), .ZN(plus[49]));
   XNOR2_X1 i_54 (.A(quotient[50]), .B(n_18), .ZN(plus[50]));
   XNOR2_X1 i_55 (.A(quotient[51]), .B(n_17), .ZN(plus[51]));
   XOR2_X1 i_56 (.A(quotient[52]), .B(n_16), .Z(plus[52]));
   XNOR2_X1 i_57 (.A(quotient[53]), .B(n_15), .ZN(plus[53]));
   XNOR2_X1 i_58 (.A(quotient[54]), .B(n_14), .ZN(plus[54]));
   XNOR2_X1 i_59 (.A(quotient[55]), .B(n_13), .ZN(plus[55]));
   XOR2_X1 i_60 (.A(quotient[56]), .B(n_12), .Z(plus[56]));
   AND2_X1 i_61 (.A1(n_11), .A2(n_5), .ZN(plus[57]));
   OAI21_X1 i_62 (.A(quotient[57]), .B1(n_12), .B2(quotient[56]), .ZN(n_5));
   XOR2_X1 i_63 (.A(quotient[58]), .B(n_11), .Z(plus[58]));
   XNOR2_X1 i_64 (.A(quotient[59]), .B(n_10), .ZN(plus[59]));
   XNOR2_X1 i_65 (.A(quotient[60]), .B(n_9), .ZN(plus[60]));
   XOR2_X1 i_66 (.A(quotient[61]), .B(n_8), .Z(plus[61]));
   XNOR2_X1 i_67 (.A(quotient[62]), .B(n_7), .ZN(plus[62]));
   XNOR2_X1 i_68 (.A(quotient[63]), .B(n_6), .ZN(plus[63]));
   NOR3_X1 i_69 (.A1(n_8), .A2(quotient[61]), .A3(quotient[62]), .ZN(n_6));
   NOR2_X1 i_70 (.A1(n_8), .A2(quotient[61]), .ZN(n_7));
   NAND2_X1 i_71 (.A1(n_9), .A2(n_72), .ZN(n_8));
   NOR3_X1 i_72 (.A1(n_11), .A2(quotient[58]), .A3(quotient[59]), .ZN(n_9));
   NOR2_X1 i_73 (.A1(n_11), .A2(quotient[58]), .ZN(n_10));
   OR3_X1 i_74 (.A1(n_12), .A2(quotient[56]), .A3(quotient[57]), .ZN(n_11));
   NAND2_X1 i_75 (.A1(n_13), .A2(n_71), .ZN(n_12));
   NOR4_X1 i_76 (.A1(n_16), .A2(quotient[52]), .A3(quotient[53]), .A4(
      quotient[54]), .ZN(n_13));
   NOR3_X1 i_77 (.A1(n_16), .A2(quotient[52]), .A3(quotient[53]), .ZN(n_14));
   NOR2_X1 i_78 (.A1(n_16), .A2(quotient[52]), .ZN(n_15));
   NAND2_X1 i_79 (.A1(n_17), .A2(n_70), .ZN(n_16));
   NOR4_X1 i_80 (.A1(n_20), .A2(quotient[48]), .A3(quotient[49]), .A4(
      quotient[50]), .ZN(n_17));
   NOR3_X1 i_81 (.A1(n_20), .A2(quotient[48]), .A3(quotient[49]), .ZN(n_18));
   NOR2_X1 i_82 (.A1(n_20), .A2(quotient[48]), .ZN(n_19));
   OR2_X1 i_83 (.A1(n_21), .A2(quotient[47]), .ZN(n_20));
   OR2_X1 i_84 (.A1(n_22), .A2(quotient[46]), .ZN(n_21));
   OR2_X1 i_85 (.A1(n_23), .A2(quotient[45]), .ZN(n_22));
   OR3_X1 i_86 (.A1(n_24), .A2(quotient[43]), .A3(quotient[44]), .ZN(n_23));
   NAND2_X1 i_87 (.A1(n_25), .A2(n_69), .ZN(n_24));
   NOR2_X1 i_88 (.A1(n_26), .A2(quotient[41]), .ZN(n_25));
   NAND2_X1 i_89 (.A1(n_27), .A2(n_68), .ZN(n_26));
   NOR3_X1 i_90 (.A1(n_29), .A2(quotient[38]), .A3(quotient[39]), .ZN(n_27));
   NOR2_X1 i_91 (.A1(n_29), .A2(quotient[38]), .ZN(n_28));
   OR2_X1 i_92 (.A1(n_30), .A2(quotient[37]), .ZN(n_29));
   NAND2_X1 i_93 (.A1(n_31), .A2(n_67), .ZN(n_30));
   NOR4_X1 i_94 (.A1(n_34), .A2(quotient[33]), .A3(quotient[34]), .A4(
      quotient[35]), .ZN(n_31));
   NOR3_X1 i_95 (.A1(n_34), .A2(quotient[33]), .A3(quotient[34]), .ZN(n_32));
   NOR2_X1 i_96 (.A1(n_34), .A2(quotient[33]), .ZN(n_33));
   OR2_X1 i_97 (.A1(n_35), .A2(quotient[32]), .ZN(n_34));
   NAND2_X1 i_98 (.A1(n_36), .A2(n_66), .ZN(n_35));
   NOR4_X1 i_99 (.A1(n_39), .A2(quotient[28]), .A3(quotient[29]), .A4(
      quotient[30]), .ZN(n_36));
   NOR3_X1 i_100 (.A1(n_39), .A2(quotient[28]), .A3(quotient[29]), .ZN(n_37));
   NOR2_X1 i_101 (.A1(n_39), .A2(quotient[28]), .ZN(n_38));
   OR2_X1 i_102 (.A1(n_40), .A2(quotient[27]), .ZN(n_39));
   NAND2_X1 i_103 (.A1(n_41), .A2(n_65), .ZN(n_40));
   NOR4_X1 i_104 (.A1(n_44), .A2(quotient[23]), .A3(quotient[24]), .A4(
      quotient[25]), .ZN(n_41));
   NOR3_X1 i_105 (.A1(n_44), .A2(quotient[23]), .A3(quotient[24]), .ZN(n_42));
   NOR2_X1 i_106 (.A1(n_44), .A2(quotient[23]), .ZN(n_43));
   OR2_X1 i_107 (.A1(n_45), .A2(quotient[22]), .ZN(n_44));
   NAND2_X1 i_108 (.A1(n_46), .A2(n_64), .ZN(n_45));
   NOR4_X1 i_109 (.A1(n_49), .A2(quotient[18]), .A3(quotient[19]), .A4(
      quotient[20]), .ZN(n_46));
   NOR3_X1 i_110 (.A1(n_49), .A2(quotient[18]), .A3(quotient[19]), .ZN(n_47));
   NOR2_X1 i_111 (.A1(n_49), .A2(quotient[18]), .ZN(n_48));
   OR2_X1 i_112 (.A1(n_50), .A2(quotient[17]), .ZN(n_49));
   OR2_X1 i_113 (.A1(n_51), .A2(quotient[16]), .ZN(n_50));
   OR3_X1 i_114 (.A1(n_52), .A2(quotient[14]), .A3(quotient[15]), .ZN(n_51));
   NAND2_X1 i_115 (.A1(n_53), .A2(n_63), .ZN(n_52));
   NOR2_X1 i_116 (.A1(n_54), .A2(quotient[12]), .ZN(n_53));
   NAND2_X1 i_117 (.A1(n_55), .A2(n_62), .ZN(n_54));
   NOR2_X1 i_118 (.A1(n_56), .A2(quotient[10]), .ZN(n_55));
   OR3_X1 i_119 (.A1(n_57), .A2(quotient[8]), .A3(quotient[9]), .ZN(n_56));
   OR2_X1 i_120 (.A1(n_58), .A2(quotient[7]), .ZN(n_57));
   OR3_X1 i_121 (.A1(n_59), .A2(quotient[5]), .A3(quotient[6]), .ZN(n_58));
   OR2_X1 i_122 (.A1(n_60), .A2(quotient[4]), .ZN(n_59));
   OR2_X1 i_123 (.A1(n_61), .A2(quotient[3]), .ZN(n_60));
   OR3_X1 i_124 (.A1(quotient[2]), .A2(quotient[1]), .A3(quotient[0]), .ZN(n_61));
   INV_X1 i_125 (.A(quotient[11]), .ZN(n_62));
   INV_X1 i_126 (.A(quotient[13]), .ZN(n_63));
   INV_X1 i_127 (.A(quotient[21]), .ZN(n_64));
   INV_X1 i_128 (.A(quotient[26]), .ZN(n_65));
   INV_X1 i_129 (.A(quotient[31]), .ZN(n_66));
   INV_X1 i_130 (.A(quotient[36]), .ZN(n_67));
   INV_X1 i_131 (.A(quotient[40]), .ZN(n_68));
   INV_X1 i_132 (.A(quotient[42]), .ZN(n_69));
   INV_X1 i_133 (.A(quotient[51]), .ZN(n_70));
   INV_X1 i_134 (.A(quotient[55]), .ZN(n_71));
   INV_X1 i_135 (.A(quotient[60]), .ZN(n_72));
endmodule

module datapath__0_153(p_0, i);
   output [31:0]p_0;
   input [31:0]i;

   XNOR2_X1 i_0 (.A(i[4]), .B(i[3]), .ZN(p_0[4]));
   XOR2_X1 i_1 (.A(i[5]), .B(n_28), .Z(p_0[5]));
   AND2_X1 i_2 (.A1(n_27), .A2(n_0), .ZN(p_0[6]));
   OAI21_X1 i_3 (.A(i[6]), .B1(i[5]), .B2(n_28), .ZN(n_0));
   XOR2_X1 i_4 (.A(i[7]), .B(n_27), .Z(p_0[7]));
   XNOR2_X1 i_5 (.A(i[8]), .B(n_26), .ZN(p_0[8]));
   XNOR2_X1 i_6 (.A(i[9]), .B(n_25), .ZN(p_0[9]));
   XOR2_X1 i_7 (.A(i[10]), .B(n_24), .Z(p_0[10]));
   XOR2_X1 i_8 (.A(i[11]), .B(n_23), .Z(p_0[11]));
   XNOR2_X1 i_9 (.A(i[12]), .B(n_22), .ZN(p_0[12]));
   XNOR2_X1 i_10 (.A(i[13]), .B(n_21), .ZN(p_0[13]));
   XNOR2_X1 i_11 (.A(i[14]), .B(n_20), .ZN(p_0[14]));
   XOR2_X1 i_12 (.A(i[15]), .B(n_19), .Z(p_0[15]));
   XOR2_X1 i_13 (.A(i[16]), .B(n_18), .Z(p_0[16]));
   AND2_X1 i_14 (.A1(n_17), .A2(n_1), .ZN(p_0[17]));
   OAI21_X1 i_15 (.A(i[17]), .B1(n_18), .B2(i[16]), .ZN(n_1));
   XOR2_X1 i_16 (.A(i[18]), .B(n_17), .Z(p_0[18]));
   XNOR2_X1 i_17 (.A(i[19]), .B(n_16), .ZN(p_0[19]));
   XOR2_X1 i_18 (.A(i[20]), .B(n_15), .Z(p_0[20]));
   XOR2_X1 i_19 (.A(i[21]), .B(n_14), .Z(p_0[21]));
   XOR2_X1 i_20 (.A(i[22]), .B(n_13), .Z(p_0[22]));
   XNOR2_X1 i_21 (.A(i[23]), .B(n_12), .ZN(p_0[23]));
   XNOR2_X1 i_22 (.A(i[24]), .B(n_11), .ZN(p_0[24]));
   XNOR2_X1 i_23 (.A(i[25]), .B(n_10), .ZN(p_0[25]));
   XNOR2_X1 i_24 (.A(i[26]), .B(n_8), .ZN(p_0[26]));
   AND2_X1 i_25 (.A1(n_6), .A2(n_2), .ZN(p_0[27]));
   OAI21_X1 i_26 (.A(i[27]), .B1(n_7), .B2(i[26]), .ZN(n_2));
   XOR2_X1 i_27 (.A(i[28]), .B(n_6), .Z(p_0[28]));
   XNOR2_X1 i_28 (.A(i[29]), .B(n_5), .ZN(p_0[29]));
   XNOR2_X1 i_29 (.A(i[30]), .B(n_4), .ZN(p_0[30]));
   XNOR2_X1 i_30 (.A(i[31]), .B(n_3), .ZN(p_0[31]));
   NOR4_X1 i_31 (.A1(n_6), .A2(i[28]), .A3(i[29]), .A4(i[30]), .ZN(n_3));
   NOR3_X1 i_32 (.A1(n_6), .A2(i[28]), .A3(i[29]), .ZN(n_4));
   NOR2_X1 i_33 (.A1(n_6), .A2(i[28]), .ZN(n_5));
   OR3_X1 i_34 (.A1(n_7), .A2(i[26]), .A3(i[27]), .ZN(n_6));
   INV_X1 i_35 (.A(n_8), .ZN(n_7));
   NOR2_X1 i_36 (.A1(n_9), .A2(i[25]), .ZN(n_8));
   INV_X1 i_37 (.A(n_10), .ZN(n_9));
   NOR4_X1 i_38 (.A1(n_13), .A2(i[22]), .A3(i[23]), .A4(i[24]), .ZN(n_10));
   NOR3_X1 i_39 (.A1(n_13), .A2(i[22]), .A3(i[23]), .ZN(n_11));
   NOR2_X1 i_40 (.A1(n_13), .A2(i[22]), .ZN(n_12));
   OR2_X1 i_41 (.A1(n_14), .A2(i[21]), .ZN(n_13));
   OR2_X1 i_42 (.A1(n_15), .A2(i[20]), .ZN(n_14));
   NAND2_X1 i_43 (.A1(n_16), .A2(n_31), .ZN(n_15));
   NOR2_X1 i_44 (.A1(n_17), .A2(i[18]), .ZN(n_16));
   OR3_X1 i_45 (.A1(n_18), .A2(i[16]), .A3(i[17]), .ZN(n_17));
   OR2_X1 i_46 (.A1(n_19), .A2(i[15]), .ZN(n_18));
   NAND2_X1 i_47 (.A1(n_20), .A2(n_30), .ZN(n_19));
   NOR4_X1 i_48 (.A1(n_23), .A2(i[11]), .A3(i[12]), .A4(i[13]), .ZN(n_20));
   NOR3_X1 i_49 (.A1(n_23), .A2(i[11]), .A3(i[12]), .ZN(n_21));
   NOR2_X1 i_50 (.A1(n_23), .A2(i[11]), .ZN(n_22));
   OR2_X1 i_51 (.A1(n_24), .A2(i[10]), .ZN(n_23));
   NAND2_X1 i_52 (.A1(n_25), .A2(n_29), .ZN(n_24));
   NOR3_X1 i_53 (.A1(n_27), .A2(i[7]), .A3(i[8]), .ZN(n_25));
   NOR2_X1 i_54 (.A1(n_27), .A2(i[7]), .ZN(n_26));
   OR3_X1 i_55 (.A1(i[6]), .A2(i[5]), .A3(n_28), .ZN(n_27));
   AND2_X1 i_56 (.A1(i[4]), .A2(i[3]), .ZN(n_28));
   INV_X1 i_57 (.A(i[1]), .ZN(p_0[1]));
   INV_X1 i_58 (.A(i[2]), .ZN(p_0[2]));
   INV_X1 i_59 (.A(i[9]), .ZN(n_29));
   INV_X1 i_60 (.A(i[14]), .ZN(n_30));
   INV_X1 i_61 (.A(i[19]), .ZN(n_31));
endmodule

module datapath__0_158(p_0, p_1);
   input [31:0]p_0;
   output [31:0]p_1;

   XNOR2_X1 i_0 (.A(p_0[1]), .B(p_0[0]), .ZN(p_1[1]));
   OR2_X1 i_1 (.A1(p_0[1]), .A2(p_0[0]), .ZN(n_0));
   XNOR2_X1 i_2 (.A(p_0[2]), .B(n_0), .ZN(p_1[2]));
   OR2_X1 i_3 (.A1(p_0[2]), .A2(n_0), .ZN(n_1));
   XNOR2_X1 i_4 (.A(p_0[3]), .B(n_1), .ZN(p_1[3]));
   OR2_X1 i_5 (.A1(p_0[3]), .A2(n_1), .ZN(n_2));
   XNOR2_X1 i_6 (.A(p_0[4]), .B(n_2), .ZN(p_1[4]));
   OR2_X1 i_7 (.A1(p_0[4]), .A2(n_2), .ZN(n_3));
   XNOR2_X1 i_8 (.A(p_0[5]), .B(n_3), .ZN(p_1[5]));
   OR2_X1 i_9 (.A1(p_0[5]), .A2(n_3), .ZN(n_4));
   XNOR2_X1 i_10 (.A(p_0[6]), .B(n_4), .ZN(p_1[6]));
   OR2_X1 i_11 (.A1(p_0[6]), .A2(n_4), .ZN(n_5));
   XNOR2_X1 i_12 (.A(p_0[7]), .B(n_5), .ZN(p_1[7]));
   OR2_X1 i_13 (.A1(p_0[7]), .A2(n_5), .ZN(n_6));
   XNOR2_X1 i_14 (.A(p_0[8]), .B(n_6), .ZN(p_1[8]));
   OR2_X1 i_15 (.A1(p_0[8]), .A2(n_6), .ZN(n_7));
   XNOR2_X1 i_16 (.A(p_0[9]), .B(n_7), .ZN(p_1[9]));
   OR2_X1 i_17 (.A1(p_0[9]), .A2(n_7), .ZN(n_8));
   XNOR2_X1 i_18 (.A(p_0[10]), .B(n_8), .ZN(p_1[10]));
   OR2_X1 i_19 (.A1(p_0[10]), .A2(n_8), .ZN(n_9));
   XNOR2_X1 i_20 (.A(p_0[11]), .B(n_9), .ZN(p_1[11]));
   OR2_X1 i_21 (.A1(p_0[11]), .A2(n_9), .ZN(n_10));
   XNOR2_X1 i_22 (.A(p_0[12]), .B(n_10), .ZN(p_1[12]));
   OR2_X1 i_23 (.A1(p_0[12]), .A2(n_10), .ZN(n_11));
   XNOR2_X1 i_24 (.A(p_0[13]), .B(n_11), .ZN(p_1[13]));
   OR2_X1 i_25 (.A1(p_0[13]), .A2(n_11), .ZN(n_12));
   XNOR2_X1 i_26 (.A(p_0[14]), .B(n_12), .ZN(p_1[14]));
   OR2_X1 i_27 (.A1(p_0[14]), .A2(n_12), .ZN(n_13));
   XNOR2_X1 i_28 (.A(p_0[15]), .B(n_13), .ZN(p_1[15]));
   OR2_X1 i_29 (.A1(p_0[15]), .A2(n_13), .ZN(n_14));
   XNOR2_X1 i_30 (.A(p_0[16]), .B(n_14), .ZN(p_1[16]));
   OR2_X1 i_31 (.A1(p_0[16]), .A2(n_14), .ZN(n_15));
   XNOR2_X1 i_32 (.A(p_0[17]), .B(n_15), .ZN(p_1[17]));
   OR2_X1 i_33 (.A1(p_0[17]), .A2(n_15), .ZN(n_16));
   XNOR2_X1 i_34 (.A(p_0[18]), .B(n_16), .ZN(p_1[18]));
   OR2_X1 i_35 (.A1(p_0[18]), .A2(n_16), .ZN(n_17));
   XNOR2_X1 i_36 (.A(p_0[19]), .B(n_17), .ZN(p_1[19]));
   OR2_X1 i_37 (.A1(p_0[19]), .A2(n_17), .ZN(n_18));
   XNOR2_X1 i_38 (.A(p_0[20]), .B(n_18), .ZN(p_1[20]));
   OR2_X1 i_39 (.A1(p_0[20]), .A2(n_18), .ZN(n_19));
   XNOR2_X1 i_40 (.A(p_0[21]), .B(n_19), .ZN(p_1[21]));
   OR2_X1 i_41 (.A1(p_0[21]), .A2(n_19), .ZN(n_20));
   XNOR2_X1 i_42 (.A(p_0[22]), .B(n_20), .ZN(p_1[22]));
   OR2_X1 i_43 (.A1(p_0[22]), .A2(n_20), .ZN(n_21));
   XNOR2_X1 i_44 (.A(p_0[23]), .B(n_21), .ZN(p_1[23]));
   OR2_X1 i_45 (.A1(p_0[23]), .A2(n_21), .ZN(n_22));
   XNOR2_X1 i_46 (.A(p_0[24]), .B(n_22), .ZN(p_1[24]));
   OR2_X1 i_47 (.A1(p_0[24]), .A2(n_22), .ZN(n_23));
   XNOR2_X1 i_48 (.A(p_0[25]), .B(n_23), .ZN(p_1[25]));
   OR2_X1 i_49 (.A1(p_0[25]), .A2(n_23), .ZN(n_24));
   XNOR2_X1 i_50 (.A(p_0[26]), .B(n_24), .ZN(p_1[26]));
   OR2_X1 i_51 (.A1(p_0[26]), .A2(n_24), .ZN(n_25));
   XNOR2_X1 i_52 (.A(p_0[27]), .B(n_25), .ZN(p_1[27]));
   OR2_X1 i_53 (.A1(p_0[27]), .A2(n_25), .ZN(n_26));
   XNOR2_X1 i_54 (.A(p_0[28]), .B(n_26), .ZN(p_1[28]));
   OR2_X1 i_55 (.A1(p_0[28]), .A2(n_26), .ZN(n_27));
   XNOR2_X1 i_56 (.A(p_0[29]), .B(n_27), .ZN(p_1[29]));
   OR2_X1 i_57 (.A1(p_0[29]), .A2(n_27), .ZN(n_28));
   XNOR2_X1 i_58 (.A(p_0[30]), .B(n_28), .ZN(p_1[30]));
   OR2_X1 i_59 (.A1(p_0[30]), .A2(n_28), .ZN(n_29));
   XNOR2_X1 i_60 (.A(p_0[31]), .B(n_29), .ZN(p_1[31]));
endmodule

module fpu_divider(mode, clk, rst, enbl, in_a, in_b, out_c, done, err, zero, 
      posv);
   input [1:0]mode;
   input clk;
   input rst;
   input enbl;
   input [63:0]in_a;
   input [63:0]in_b;
   output [63:0]out_c;
   output done;
   output err;
   output zero;
   output posv;

   wire [63:0]sub;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire [31:0]i;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire [1:0]state;
   wire n_0_217;
   wire [63:0]z;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_166;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_180;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_190;
   wire n_0_191;
   wire n_0_192;
   wire n_0_193;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_200;
   wire n_0_201;
   wire n_0_202;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_207;
   wire n_0_208;
   wire n_0_209;
   wire n_0_210;
   wire n_0_211;
   wire n_0_212;
   wire n_0_213;
   wire n_0_214;
   wire n_0_215;
   wire n_0_216;
   wire n_0_218;
   wire n_0_219;
   wire n_0_220;
   wire n_0_221;
   wire n_0_222;
   wire n_0_223;
   wire n_0_224;
   wire n_0_225;
   wire posv_sig;
   wire zero_sig;
   wire ovfl_sig;
   wire div_by_zero_sig;
   wire [63:0]out_sig;
   wire done_sig;
   wire n_0_226;
   wire n_0_227;
   wire n_0_228;
   wire n_0_229;
   wire n_0_230;
   wire n_0_366;
   wire n_0_367;
   wire n_0_368;
   wire n_0_369;
   wire n_0_370;
   wire n_0_371;
   wire n_0_372;
   wire n_0_373;
   wire n_0_374;
   wire n_0_375;
   wire n_0_376;
   wire n_0_377;
   wire n_0_378;
   wire n_0_379;
   wire n_0_380;
   wire n_0_381;
   wire n_0_382;
   wire n_0_383;
   wire n_0_384;
   wire n_0_385;
   wire n_0_386;
   wire n_0_387;
   wire n_0_388;
   wire n_0_389;
   wire n_0_390;
   wire [63:0]quotient;
   wire n_0_393;
   wire n_0_394;
   wire n_0_395;
   wire n_0_396;
   wire n_0_397;
   wire n_0_398;
   wire n_0_399;
   wire n_0_400;
   wire n_0_401;
   wire n_0_402;
   wire n_0_403;
   wire n_0_404;
   wire n_0_405;
   wire n_0_406;
   wire n_0_407;
   wire n_0_408;
   wire n_0_409;
   wire n_0_410;
   wire n_0_411;
   wire n_0_412;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_231;
   wire n_0_2_0;
   wire n_0_298;
   wire n_0_2_1;
   wire n_0_2_2;
   wire n_0_2_3;
   wire n_0_2_4;
   wire n_0_2_5;
   wire n_0_2_6;
   wire n_0_2_7;
   wire n_0_2_8;
   wire n_0_2_9;
   wire n_0_2_10;
   wire n_0_2_11;
   wire n_0_2_12;
   wire n_0_2_13;
   wire n_0_2_14;
   wire n_0_2_15;
   wire n_0_2_16;
   wire n_0_2_17;
   wire n_0_2_18;
   wire n_0_232;
   wire n_0_2_19;
   wire n_0_233;
   wire n_0_2_20;
   wire n_0_2_21;
   wire n_0_234;
   wire n_0_2_22;
   wire n_0_235;
   wire n_0_2_23;
   wire n_0_236;
   wire n_0_2_24;
   wire n_0_237;
   wire n_0_2_25;
   wire n_0_238;
   wire n_0_2_26;
   wire n_0_239;
   wire n_0_2_27;
   wire n_0_2_28;
   wire n_0_2_29;
   wire n_0_240;
   wire n_0_241;
   wire n_0_242;
   wire n_0_243;
   wire n_0_244;
   wire n_0_245;
   wire n_0_246;
   wire n_0_247;
   wire n_0_2_30;
   wire n_0_2_31;
   wire n_0_2_32;
   wire n_0_248;
   wire n_0_249;
   wire n_0_250;
   wire n_0_251;
   wire n_0_252;
   wire n_0_253;
   wire n_0_254;
   wire n_0_255;
   wire n_0_2_33;
   wire n_0_2_34;
   wire n_0_256;
   wire n_0_257;
   wire n_0_258;
   wire n_0_259;
   wire n_0_260;
   wire n_0_261;
   wire n_0_262;
   wire n_0_263;
   wire n_0_2_35;
   wire n_0_264;
   wire n_0_265;
   wire n_0_266;
   wire n_0_267;
   wire n_0_268;
   wire n_0_269;
   wire n_0_270;
   wire n_0_271;
   wire n_0_2_36;
   wire n_0_272;
   wire n_0_273;
   wire n_0_274;
   wire n_0_275;
   wire n_0_276;
   wire n_0_277;
   wire n_0_278;
   wire n_0_279;
   wire n_0_2_37;
   wire n_0_280;
   wire n_0_281;
   wire n_0_282;
   wire n_0_283;
   wire n_0_284;
   wire n_0_285;
   wire n_0_286;
   wire n_0_287;
   wire n_0_2_38;
   wire n_0_288;
   wire n_0_289;
   wire n_0_290;
   wire n_0_291;
   wire n_0_292;
   wire n_0_293;
   wire n_0_294;
   wire n_0_295;
   wire n_0_2_39;
   wire n_0_2_40;
   wire [63:0]b;
   wire n_0_2_41;
   wire n_0_2_42;
   wire n_0_2_43;
   wire n_0_2_44;
   wire n_0_2_45;
   wire n_0_2_46;
   wire n_0_2_47;
   wire n_0_2_48;
   wire n_0_2_49;
   wire n_0_2_50;
   wire n_0_2_51;
   wire n_0_2_52;
   wire n_0_2_53;
   wire n_0_2_54;
   wire n_0_2_55;
   wire n_0_2_56;
   wire n_0_2_57;
   wire n_0_2_58;
   wire n_0_2_59;
   wire n_0_2_60;
   wire n_0_2_61;
   wire n_0_2_62;
   wire n_0_2_63;
   wire n_0_2_64;
   wire n_0_2_65;
   wire n_0_2_66;
   wire n_0_2_67;
   wire n_0_2_68;
   wire n_0_2_69;
   wire n_0_2_70;
   wire n_0_2_71;
   wire n_0_2_72;
   wire n_0_2_73;
   wire n_0_2_74;
   wire n_0_2_75;
   wire n_0_2_76;
   wire n_0_2_77;
   wire n_0_2_78;
   wire n_0_2_79;
   wire n_0_2_80;
   wire n_0_2_81;
   wire n_0_2_82;
   wire n_0_2_83;
   wire n_0_2_84;
   wire n_0_2_85;
   wire n_0_2_86;
   wire n_0_2_87;
   wire n_0_2_88;
   wire n_0_2_89;
   wire n_0_2_90;
   wire n_0_2_91;
   wire n_0_2_92;
   wire n_0_2_93;
   wire n_0_2_94;
   wire n_0_2_95;
   wire n_0_2_96;
   wire n_0_2_97;
   wire n_0_2_98;
   wire n_0_2_99;
   wire n_0_2_100;
   wire n_0_2_101;
   wire n_0_2_102;
   wire n_0_2_103;
   wire n_0_2_104;
   wire n_0_2_105;
   wire n_0_2_106;
   wire n_0_2_107;
   wire n_0_2_108;
   wire n_0_2_109;
   wire n_0_2_110;
   wire n_0_2_111;
   wire n_0_2_112;
   wire n_0_2_113;
   wire n_0_2_114;
   wire n_0_2_115;
   wire n_0_2_116;
   wire n_0_2_117;
   wire n_0_2_118;
   wire n_0_2_119;
   wire n_0_2_120;
   wire n_0_2_121;
   wire n_0_2_122;
   wire n_0_2_123;
   wire n_0_2_124;
   wire n_0_2_125;
   wire n_0_2_126;
   wire n_0_2_127;
   wire n_0_2_128;
   wire n_0_2_129;
   wire n_0_2_130;
   wire n_0_2_131;
   wire n_0_2_132;
   wire n_0_2_133;
   wire n_0_2_134;
   wire n_0_2_135;
   wire n_0_2_136;
   wire n_0_2_137;
   wire n_0_2_138;
   wire n_0_2_139;
   wire n_0_2_140;
   wire n_0_2_141;
   wire n_0_2_142;
   wire n_0_2_143;
   wire n_0_2_144;
   wire n_0_2_145;
   wire n_0_2_146;
   wire n_0_2_147;
   wire n_0_2_148;
   wire n_0_2_149;
   wire n_0_2_150;
   wire n_0_2_151;
   wire n_0_2_152;
   wire n_0_2_153;
   wire n_0_2_154;
   wire n_0_2_155;
   wire n_0_2_156;
   wire n_0_2_157;
   wire n_0_2_158;
   wire n_0_2_159;
   wire n_0_2_160;
   wire n_0_2_161;
   wire n_0_2_162;
   wire n_0_2_163;
   wire n_0_2_164;
   wire n_0_2_165;
   wire n_0_2_166;
   wire n_0_2_167;
   wire n_0_2_168;
   wire n_0_2_169;
   wire n_0_2_170;
   wire n_0_2_171;
   wire n_0_2_172;
   wire n_0_2_173;
   wire n_0_2_174;
   wire n_0_2_175;
   wire n_0_2_176;
   wire n_0_2_177;
   wire n_0_2_178;
   wire n_0_2_179;
   wire n_0_2_180;
   wire n_0_2_181;
   wire n_0_2_182;
   wire n_0_2_183;
   wire n_0_2_184;
   wire n_0_2_185;
   wire n_0_2_186;
   wire n_0_2_187;
   wire n_0_2_188;
   wire n_0_2_189;
   wire n_0_2_190;
   wire n_0_2_191;
   wire n_0_2_192;
   wire n_0_2_193;
   wire n_0_2_194;
   wire n_0_2_195;
   wire n_0_2_196;
   wire n_0_2_197;
   wire n_0_2_198;
   wire n_0_2_199;
   wire n_0_2_200;
   wire n_0_2_201;
   wire n_0_2_202;
   wire n_0_2_203;
   wire n_0_2_204;
   wire n_0_2_205;
   wire n_0_2_206;
   wire n_0_2_207;
   wire n_0_2_208;
   wire n_0_2_209;
   wire n_0_2_210;
   wire n_0_2_211;
   wire n_0_2_212;
   wire n_0_2_213;
   wire n_0_2_214;
   wire n_0_2_215;
   wire n_0_2_216;
   wire n_0_2_217;
   wire n_0_2_218;
   wire n_0_2_219;
   wire n_0_2_220;
   wire n_0_2_221;
   wire n_0_2_222;
   wire n_0_2_223;
   wire n_0_2_224;
   wire n_0_2_225;
   wire n_0_2_226;
   wire n_0_2_227;
   wire n_0_2_228;
   wire n_0_2_229;
   wire n_0_296;
   wire n_0_2_230;
   wire n_0_2_231;
   wire n_0_2_232;
   wire n_0_2_233;
   wire n_0_2_234;
   wire n_0_2_235;
   wire n_0_2_236;
   wire n_0_2_237;
   wire n_0_2_238;
   wire n_0_2_239;
   wire n_0_2_240;
   wire n_0_2_241;
   wire n_0_2_242;
   wire n_0_2_243;
   wire n_0_2_244;
   wire n_0_2_245;
   wire n_0_2_246;
   wire n_0_2_247;
   wire n_0_2_248;
   wire n_0_2_249;
   wire n_0_2_250;
   wire n_0_2_251;
   wire n_0_2_252;
   wire n_0_2_253;
   wire n_0_2_254;
   wire n_0_2_255;
   wire n_0_2_256;
   wire n_0_2_257;
   wire n_0_2_258;
   wire n_0_2_259;
   wire n_0_2_260;
   wire n_0_2_261;
   wire n_0_2_262;
   wire n_0_2_263;
   wire n_0_2_264;
   wire n_0_2_265;
   wire n_0_2_266;
   wire n_0_2_267;
   wire n_0_2_268;
   wire n_0_2_269;
   wire n_0_2_270;
   wire n_0_2_271;
   wire n_0_2_272;
   wire n_0_2_273;
   wire n_0_2_274;
   wire n_0_2_275;
   wire n_0_2_276;
   wire n_0_2_277;
   wire n_0_2_278;
   wire n_0_2_279;
   wire n_0_2_280;
   wire n_0_2_281;
   wire n_0_2_282;
   wire n_0_2_283;
   wire n_0_2_284;
   wire n_0_2_285;
   wire n_0_2_286;
   wire n_0_2_287;
   wire n_0_2_288;
   wire n_0_2_289;
   wire n_0_2_290;
   wire n_0_2_291;
   wire n_0_2_292;
   wire n_0_2_293;
   wire n_0_2_294;
   wire n_0_2_295;
   wire n_0_2_296;
   wire n_0_2_297;
   wire n_0_2_298;
   wire n_0_2_299;
   wire n_0_2_300;
   wire n_0_2_301;
   wire n_0_2_302;
   wire n_0_2_303;
   wire n_0_2_304;
   wire n_0_2_305;
   wire n_0_2_306;
   wire n_0_2_307;
   wire n_0_2_308;
   wire n_0_2_309;
   wire n_0_2_310;
   wire n_0_2_311;
   wire n_0_2_312;
   wire n_0_2_313;
   wire n_0_2_314;
   wire n_0_2_315;
   wire n_0_2_316;
   wire n_0_2_317;
   wire n_0_2_318;
   wire n_0_2_319;
   wire n_0_2_320;
   wire n_0_2_321;
   wire n_0_2_322;
   wire n_0_2_323;
   wire n_0_2_324;
   wire n_0_2_325;
   wire n_0_2_326;
   wire n_0_2_327;
   wire n_0_2_328;
   wire n_0_2_329;
   wire n_0_2_330;
   wire n_0_2_331;
   wire n_0_2_332;
   wire n_0_2_333;
   wire n_0_2_334;
   wire n_0_2_335;
   wire n_0_2_336;
   wire n_0_2_337;
   wire n_0_2_338;
   wire n_0_2_339;
   wire n_0_2_340;
   wire n_0_2_341;
   wire n_0_2_342;
   wire n_0_2_343;
   wire n_0_2_344;
   wire n_0_2_345;
   wire n_0_2_346;
   wire n_0_2_347;
   wire [63:0]z_next_reg;
   wire n_0_2_348;
   wire n_0_2_349;
   wire n_0_2_350;
   wire n_0_2_351;
   wire n_0_2_352;
   wire n_0_2_353;
   wire n_0_2_354;
   wire n_0_2_355;
   wire n_0_2_356;
   wire n_0_2_357;
   wire n_0_2_358;
   wire n_0_2_359;
   wire n_0_2_360;
   wire n_0_2_361;
   wire n_0_2_362;
   wire n_0_2_363;
   wire n_0_2_364;
   wire n_0_2_365;
   wire n_0_2_366;
   wire n_0_2_367;
   wire n_0_2_368;
   wire n_0_2_369;
   wire n_0_2_370;
   wire n_0_2_371;
   wire n_0_2_372;
   wire n_0_2_373;
   wire n_0_2_374;
   wire n_0_2_375;
   wire n_0_2_376;
   wire n_0_2_377;
   wire n_0_2_378;
   wire n_0_2_379;
   wire n_0_2_380;
   wire n_0_2_381;
   wire n_0_2_382;
   wire n_0_2_383;
   wire n_0_2_384;
   wire n_0_2_385;
   wire n_0_2_386;
   wire n_0_2_387;
   wire n_0_2_388;
   wire n_0_2_389;
   wire n_0_2_390;
   wire n_0_2_391;
   wire n_0_2_392;
   wire n_0_2_393;
   wire n_0_2_394;
   wire n_0_2_395;
   wire n_0_2_396;
   wire n_0_2_397;
   wire n_0_2_398;
   wire n_0_2_399;
   wire n_0_2_400;
   wire n_0_2_401;
   wire n_0_2_402;
   wire n_0_2_403;
   wire n_0_2_404;
   wire n_0_2_405;
   wire n_0_2_406;
   wire n_0_2_407;
   wire n_0_2_408;
   wire n_0_2_409;
   wire n_0_2_410;
   wire n_0_297;
   wire n_0_2_411;
   wire [31:0]i_next_reg;
   wire n_0_2_412;
   wire n_0_2_413;
   wire n_0_2_414;
   wire n_0_2_415;
   wire n_0_2_416;
   wire n_0_2_417;
   wire n_0_2_418;
   wire n_0_2_419;
   wire n_0_2_420;
   wire n_0_2_421;
   wire n_0_2_422;
   wire n_0_2_423;
   wire n_0_2_424;
   wire n_0_2_425;
   wire n_0_2_426;
   wire n_0_2_427;
   wire n_0_2_428;
   wire n_0_2_429;
   wire n_0_2_430;
   wire n_0_2_431;
   wire n_0_2_432;
   wire n_0_2_433;
   wire n_0_2_434;
   wire n_0_2_435;
   wire n_0_2_436;
   wire n_0_2_437;
   wire n_0_2_438;
   wire n_0_2_439;
   wire n_0_2_440;
   wire n_0_2_441;
   wire n_0_2_442;
   wire n_0_2_443;
   wire n_0_2_444;
   wire n_0_2_445;
   wire n_0_2_446;
   wire n_0_2_447;
   wire n_0_2_448;
   wire n_0_2_449;
   wire n_0_2_450;
   wire n_0_2_451;
   wire n_0_2_452;
   wire n_0_2_453;
   wire n_0_2_454;
   wire n_0_2_455;
   wire n_0_2_456;
   wire n_0_2_457;
   wire n_0_299;
   wire n_0_2_458;
   wire n_0_2_459;
   wire n_0_2_460;
   wire n_0_2_461;
   wire n_0_2_462;
   wire n_0_300;
   wire n_0_2_463;
   wire n_0_301;
   wire n_0_2_464;
   wire n_0_302;
   wire n_0_2_465;
   wire n_0_303;
   wire n_0_2_466;
   wire n_0_304;
   wire n_0_2_467;
   wire n_0_305;
   wire n_0_2_468;
   wire n_0_306;
   wire n_0_2_469;
   wire n_0_307;
   wire n_0_2_470;
   wire n_0_308;
   wire n_0_2_471;
   wire n_0_309;
   wire n_0_2_472;
   wire n_0_310;
   wire n_0_2_473;
   wire n_0_311;
   wire n_0_2_474;
   wire n_0_312;
   wire n_0_2_475;
   wire n_0_313;
   wire n_0_2_476;
   wire n_0_314;
   wire n_0_2_477;
   wire n_0_315;
   wire n_0_2_478;
   wire n_0_316;
   wire n_0_2_479;
   wire n_0_317;
   wire n_0_2_480;
   wire n_0_318;
   wire n_0_2_481;
   wire n_0_319;
   wire n_0_2_482;
   wire n_0_320;
   wire n_0_2_483;
   wire n_0_321;
   wire n_0_2_484;
   wire n_0_322;
   wire n_0_2_485;
   wire n_0_323;
   wire n_0_2_486;
   wire n_0_324;
   wire n_0_2_487;
   wire n_0_325;
   wire n_0_2_488;
   wire n_0_326;
   wire n_0_2_489;
   wire n_0_327;
   wire n_0_2_490;
   wire n_0_328;
   wire n_0_2_491;
   wire n_0_329;
   wire n_0_2_492;
   wire n_0_330;
   wire n_0_2_493;
   wire n_0_331;
   wire n_0_2_494;
   wire n_0_332;
   wire n_0_2_495;
   wire n_0_333;
   wire n_0_2_496;
   wire n_0_334;
   wire n_0_2_497;
   wire n_0_335;
   wire n_0_2_498;
   wire n_0_336;
   wire n_0_2_499;
   wire n_0_337;
   wire n_0_2_500;
   wire n_0_338;
   wire n_0_2_501;
   wire n_0_339;
   wire n_0_2_502;
   wire n_0_340;
   wire n_0_2_503;
   wire n_0_341;
   wire n_0_2_504;
   wire n_0_342;
   wire n_0_2_505;
   wire n_0_343;
   wire n_0_2_506;
   wire n_0_344;
   wire n_0_2_507;
   wire n_0_345;
   wire n_0_2_508;
   wire n_0_346;
   wire n_0_2_509;
   wire n_0_347;
   wire n_0_2_510;
   wire n_0_348;
   wire n_0_2_511;
   wire n_0_349;
   wire n_0_2_512;
   wire n_0_350;
   wire n_0_2_513;
   wire n_0_351;
   wire n_0_2_514;
   wire n_0_352;
   wire n_0_2_515;
   wire n_0_353;
   wire n_0_2_516;
   wire n_0_354;
   wire n_0_2_517;
   wire n_0_355;
   wire n_0_2_518;
   wire n_0_356;
   wire n_0_2_519;
   wire n_0_357;
   wire n_0_2_520;
   wire n_0_358;
   wire n_0_2_521;
   wire n_0_359;
   wire n_0_2_522;
   wire n_0_360;
   wire n_0_2_523;
   wire n_0_361;
   wire n_0_2_524;
   wire n_0_362;
   wire n_0_2_525;
   wire n_0_2_526;
   wire n_0_2_527;
   wire n_0_2_528;
   wire n_0_2_529;
   wire n_0_2_530;
   wire n_0_2_531;
   wire n_0_2_532;
   wire n_0_2_533;
   wire n_0_2_534;
   wire n_0_2_535;
   wire n_0_2_536;
   wire n_0_2_537;
   wire n_0_2_538;
   wire n_0_2_539;
   wire n_0_2_540;
   wire n_0_2_541;
   wire n_0_2_542;
   wire n_0_2_543;
   wire n_0_2_544;
   wire n_0_2_545;
   wire n_0_2_546;
   wire n_0_2_547;
   wire n_0_363;
   wire n_0_2_548;
   wire n_0_2_549;
   wire n_0_2_550;
   wire n_0_364;
   wire n_0_2_551;
   wire n_0_2_552;
   wire n_0_2_553;
   wire n_0_2_554;
   wire n_0_2_555;
   wire n_0_2_556;
   wire n_0_2_557;
   wire n_0_2_558;
   wire n_0_2_559;
   wire n_0_2_560;
   wire n_0_2_561;
   wire n_0_2_562;
   wire n_0_2_563;
   wire n_0_2_564;
   wire n_0_2_565;
   wire n_0_2_566;
   wire n_0_2_567;
   wire n_0_2_568;
   wire n_0_2_569;
   wire n_0_2_570;
   wire n_0_2_571;
   wire n_0_2_572;
   wire n_0_2_573;
   wire n_0_2_574;
   wire n_0_2_575;
   wire n_0_2_576;
   wire n_0_2_577;
   wire n_0_365;
   wire n_0_2_578;
   wire n_0_391;
   wire n_0_2_579;
   wire n_0_392;
   wire n_0_2_580;
   wire n_0_2_581;
   wire n_0_2_582;
   wire [1:0]state_next_reg;

   fpu_adder subtractor (.mode(), .clk(), .rst(rst), .enbl(), .add_sub(), 
      .in_a(z), .in_b({b[63], b[62], b[61], b[60], b[59], b[58], b[57], b[56], 
      b[55], b[54], b[53], b[52], b[51], b[50], b[49], b[48], b[47], b[46], 
      b[45], b[44], b[43], b[42], b[41], b[40], b[39], b[38], b[37], b[36], 
      b[35], b[34], b[33], b[32], b[31], b[30], b[29], b[28], b[27], b[26], 
      b[25], b[24], b[23], b[22], b[21], b[20], b[19], b[18], b[17], b[16], 
      b[15], b[14], b[13], b[12], b[11], b[10], b[9], b[8], b[7], b[6], b[5], 
      b[4], b[3], b[2], b[1], in_b[0]}), .out_c(sub), .done(), .err(), .zero(), 
      .posv());
   datapath__0_143 i_0_0 (.in_b(in_b), .p_0({n_0_73, n_0_72, n_0_71, n_0_70, 
      n_0_69, n_0_68, n_0_67, n_0_66, n_0_65, n_0_64, n_0_63, n_0_62, n_0_61, 
      n_0_60, n_0_59, n_0_58, n_0_57, n_0_56, n_0_55, n_0_54, n_0_53, n_0_52, 
      n_0_51, n_0_50, n_0_49, n_0_48, n_0_47, n_0_46, n_0_45, n_0_44, n_0_43, 
      n_0_42, n_0_41, n_0_40, n_0_39, n_0_38, n_0_37, n_0_36, n_0_35, n_0_34, 
      n_0_33, n_0_32, n_0_31, n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, 
      n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, n_0_17, n_0_16, 
      n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, uc_0}));
   datapath__0_146 i_0_3 (.in_a({uc_1, uc_2, uc_3, uc_4, uc_5, uc_6, uc_7, 
      in_a[56], in_a[55], in_a[54], in_a[53], in_a[52], in_a[51], in_a[50], 
      in_a[49], in_a[48], in_a[47], in_a[46], in_a[45], in_a[44], in_a[43], 
      in_a[42], in_a[41], in_a[40], in_a[39], in_a[38], in_a[37], in_a[36], 
      in_a[35], in_a[34], in_a[33], in_a[32], in_a[31], in_a[30], in_a[29], 
      in_a[28], in_a[27], in_a[26], in_a[25], in_a[24], in_a[23], in_a[22], 
      in_a[21], in_a[20], in_a[19], in_a[18], in_a[17], in_a[16], in_a[15], 
      in_a[14], in_a[13], in_a[12], in_a[11], in_a[10], in_a[9], in_a[8], 
      in_a[7], in_a[6], in_a[5], in_a[4], in_a[3], in_a[2], in_a[1], in_a[0]}), 
      .p_0({uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, n_0_129, n_0_128, 
      n_0_127, n_0_126, n_0_125, n_0_124, n_0_123, n_0_122, n_0_121, n_0_120, 
      n_0_119, n_0_118, n_0_117, n_0_116, n_0_115, n_0_114, n_0_113, n_0_112, 
      n_0_111, n_0_110, n_0_109, n_0_108, n_0_107, n_0_106, n_0_105, n_0_104, 
      n_0_103, n_0_102, n_0_101, n_0_100, n_0_99, n_0_98, n_0_97, n_0_96, n_0_95, 
      n_0_94, n_0_93, n_0_92, n_0_91, n_0_90, n_0_89, n_0_88, n_0_87, n_0_86, 
      n_0_85, n_0_84, n_0_83, n_0_82, n_0_81, n_0_80, n_0_79, n_0_78, n_0_77, 
      n_0_76, n_0_75, n_0_74, uc_15}));
   DFFR_X1 \i_reg[31]  (.D(i_next_reg[31]), .RN(n_0_231), .CK(clk), .Q(i[31]), 
      .QN());
   DFFR_X1 \i_reg[30]  (.D(i_next_reg[30]), .RN(n_0_231), .CK(clk), .Q(i[30]), 
      .QN());
   DFFR_X1 \i_reg[29]  (.D(i_next_reg[29]), .RN(n_0_231), .CK(clk), .Q(i[29]), 
      .QN());
   DFFR_X1 \i_reg[28]  (.D(i_next_reg[28]), .RN(n_0_231), .CK(clk), .Q(i[28]), 
      .QN());
   DFFR_X1 \i_reg[27]  (.D(i_next_reg[27]), .RN(n_0_231), .CK(clk), .Q(i[27]), 
      .QN());
   DFFR_X1 \i_reg[26]  (.D(i_next_reg[26]), .RN(n_0_231), .CK(clk), .Q(i[26]), 
      .QN());
   DFFR_X1 \i_reg[25]  (.D(i_next_reg[25]), .RN(n_0_231), .CK(clk), .Q(i[25]), 
      .QN());
   DFFR_X1 \i_reg[24]  (.D(i_next_reg[24]), .RN(n_0_231), .CK(clk), .Q(i[24]), 
      .QN());
   DFFR_X1 \i_reg[23]  (.D(i_next_reg[23]), .RN(n_0_231), .CK(clk), .Q(i[23]), 
      .QN());
   DFFR_X1 \i_reg[22]  (.D(i_next_reg[22]), .RN(n_0_231), .CK(clk), .Q(i[22]), 
      .QN());
   DFFR_X1 \i_reg[21]  (.D(i_next_reg[21]), .RN(n_0_231), .CK(clk), .Q(i[21]), 
      .QN());
   DFFR_X1 \i_reg[20]  (.D(i_next_reg[20]), .RN(n_0_231), .CK(clk), .Q(i[20]), 
      .QN());
   DFFR_X1 \i_reg[19]  (.D(i_next_reg[19]), .RN(n_0_231), .CK(clk), .Q(i[19]), 
      .QN());
   DFFR_X1 \i_reg[18]  (.D(i_next_reg[18]), .RN(n_0_231), .CK(clk), .Q(i[18]), 
      .QN());
   DFFR_X1 \i_reg[17]  (.D(i_next_reg[17]), .RN(n_0_231), .CK(clk), .Q(i[17]), 
      .QN());
   DFFR_X1 \i_reg[16]  (.D(i_next_reg[16]), .RN(n_0_231), .CK(clk), .Q(i[16]), 
      .QN());
   DFFR_X1 \i_reg[15]  (.D(i_next_reg[15]), .RN(n_0_231), .CK(clk), .Q(i[15]), 
      .QN());
   DFFR_X1 \i_reg[14]  (.D(i_next_reg[14]), .RN(n_0_231), .CK(clk), .Q(i[14]), 
      .QN());
   DFFR_X1 \i_reg[13]  (.D(i_next_reg[13]), .RN(n_0_231), .CK(clk), .Q(i[13]), 
      .QN());
   DFFR_X1 \i_reg[12]  (.D(i_next_reg[12]), .RN(n_0_231), .CK(clk), .Q(i[12]), 
      .QN());
   DFFR_X1 \i_reg[11]  (.D(i_next_reg[11]), .RN(n_0_231), .CK(clk), .Q(i[11]), 
      .QN());
   DFFR_X1 \i_reg[10]  (.D(i_next_reg[10]), .RN(n_0_231), .CK(clk), .Q(i[10]), 
      .QN());
   DFFR_X1 \i_reg[9]  (.D(i_next_reg[9]), .RN(n_0_231), .CK(clk), .Q(i[9]), 
      .QN());
   DFFR_X1 \i_reg[8]  (.D(i_next_reg[8]), .RN(n_0_231), .CK(clk), .Q(i[8]), 
      .QN());
   DFFR_X1 \i_reg[7]  (.D(i_next_reg[7]), .RN(n_0_231), .CK(clk), .Q(i[7]), 
      .QN());
   DFFR_X1 \i_reg[6]  (.D(i_next_reg[6]), .RN(n_0_231), .CK(clk), .Q(i[6]), 
      .QN());
   DFFR_X1 \i_reg[5]  (.D(i_next_reg[5]), .RN(n_0_231), .CK(clk), .Q(i[5]), 
      .QN());
   DFFR_X1 \i_reg[4]  (.D(i_next_reg[4]), .RN(n_0_231), .CK(clk), .Q(i[4]), 
      .QN());
   DFFR_X1 \i_reg[3]  (.D(i_next_reg[3]), .RN(n_0_231), .CK(clk), .Q(i[3]), 
      .QN());
   DFFR_X1 \i_reg[2]  (.D(i_next_reg[2]), .RN(n_0_231), .CK(clk), .Q(i[2]), 
      .QN());
   DFFR_X1 \i_reg[1]  (.D(i_next_reg[1]), .RN(n_0_231), .CK(clk), .Q(i[1]), 
      .QN());
   DFFR_X1 \i_reg[0]  (.D(i_next_reg[0]), .RN(n_0_231), .CK(clk), .Q(i[0]), 
      .QN());
   datapath__0_43 i_0_7 (.i(i), .p_0({n_0_161, n_0_160, n_0_159, n_0_158, 
      n_0_157, n_0_156, n_0_155, n_0_154, n_0_153, n_0_152, n_0_151, n_0_150, 
      n_0_149, n_0_148, n_0_147, n_0_146, n_0_145, n_0_144, n_0_143, n_0_142, 
      n_0_141, n_0_140, n_0_139, n_0_138, n_0_137, n_0_136, n_0_135, n_0_134, 
      n_0_133, n_0_132, n_0_131, n_0_130}));
   DFFR_X1 \state_reg[1]  (.D(state[0]), .RN(n_0_231), .CK(clk), .Q(state[1]), 
      .QN());
   DFFR_X1 \state_reg[0]  (.D(state_next_reg[0]), .RN(n_0_231), .CK(clk), 
      .Q(state[0]), .QN());
   CLKGATETST_X1 clk_gate_z_reg (.CK(clk), .E(n_0_297), .SE(1'b0), .GCK(n_0_217));
   DFFR_X1 \z_reg[63]  (.D(z_next_reg[63]), .RN(n_0_231), .CK(n_0_217), .Q(z[63]), 
      .QN());
   DFFR_X1 \z_reg[62]  (.D(z_next_reg[62]), .RN(n_0_231), .CK(n_0_217), .Q(z[62]), 
      .QN());
   DFFR_X1 \z_reg[61]  (.D(z_next_reg[61]), .RN(n_0_231), .CK(n_0_217), .Q(z[61]), 
      .QN());
   DFFR_X1 \z_reg[60]  (.D(z_next_reg[60]), .RN(n_0_231), .CK(n_0_217), .Q(z[60]), 
      .QN());
   DFFR_X1 \z_reg[59]  (.D(z_next_reg[59]), .RN(n_0_231), .CK(n_0_217), .Q(z[59]), 
      .QN());
   DFFR_X1 \z_reg[58]  (.D(z_next_reg[58]), .RN(n_0_231), .CK(n_0_217), .Q(z[58]), 
      .QN());
   DFFR_X1 \z_reg[57]  (.D(z_next_reg[57]), .RN(n_0_231), .CK(n_0_217), .Q(z[57]), 
      .QN());
   DFFR_X1 \z_reg[56]  (.D(z_next_reg[56]), .RN(n_0_231), .CK(n_0_217), .Q(z[56]), 
      .QN());
   DFFR_X1 \z_reg[55]  (.D(z_next_reg[55]), .RN(n_0_231), .CK(n_0_217), .Q(z[55]), 
      .QN());
   DFFR_X1 \z_reg[54]  (.D(z_next_reg[54]), .RN(n_0_231), .CK(n_0_217), .Q(z[54]), 
      .QN());
   DFFR_X1 \z_reg[53]  (.D(z_next_reg[53]), .RN(n_0_231), .CK(n_0_217), .Q(z[53]), 
      .QN());
   DFFR_X1 \z_reg[52]  (.D(z_next_reg[52]), .RN(n_0_231), .CK(n_0_217), .Q(z[52]), 
      .QN());
   DFFR_X1 \z_reg[51]  (.D(z_next_reg[51]), .RN(n_0_231), .CK(n_0_217), .Q(z[51]), 
      .QN());
   DFFR_X1 \z_reg[50]  (.D(z_next_reg[50]), .RN(n_0_231), .CK(n_0_217), .Q(z[50]), 
      .QN());
   DFFR_X1 \z_reg[49]  (.D(z_next_reg[49]), .RN(n_0_231), .CK(n_0_217), .Q(z[49]), 
      .QN());
   DFFR_X1 \z_reg[48]  (.D(z_next_reg[48]), .RN(n_0_231), .CK(n_0_217), .Q(z[48]), 
      .QN());
   DFFR_X1 \z_reg[47]  (.D(z_next_reg[47]), .RN(n_0_231), .CK(n_0_217), .Q(z[47]), 
      .QN());
   DFFR_X1 \z_reg[46]  (.D(z_next_reg[46]), .RN(n_0_231), .CK(n_0_217), .Q(z[46]), 
      .QN());
   DFFR_X1 \z_reg[45]  (.D(z_next_reg[45]), .RN(n_0_231), .CK(n_0_217), .Q(z[45]), 
      .QN());
   DFFR_X1 \z_reg[44]  (.D(z_next_reg[44]), .RN(n_0_231), .CK(n_0_217), .Q(z[44]), 
      .QN());
   DFFR_X1 \z_reg[43]  (.D(z_next_reg[43]), .RN(n_0_231), .CK(n_0_217), .Q(z[43]), 
      .QN());
   DFFR_X1 \z_reg[42]  (.D(z_next_reg[42]), .RN(n_0_231), .CK(n_0_217), .Q(z[42]), 
      .QN());
   DFFR_X1 \z_reg[41]  (.D(z_next_reg[41]), .RN(n_0_231), .CK(n_0_217), .Q(z[41]), 
      .QN());
   DFFR_X1 \z_reg[40]  (.D(z_next_reg[40]), .RN(n_0_231), .CK(n_0_217), .Q(z[40]), 
      .QN());
   DFFR_X1 \z_reg[39]  (.D(z_next_reg[39]), .RN(n_0_231), .CK(n_0_217), .Q(z[39]), 
      .QN());
   DFFR_X1 \z_reg[38]  (.D(z_next_reg[38]), .RN(n_0_231), .CK(n_0_217), .Q(z[38]), 
      .QN());
   DFFR_X1 \z_reg[37]  (.D(z_next_reg[37]), .RN(n_0_231), .CK(n_0_217), .Q(z[37]), 
      .QN());
   DFFR_X1 \z_reg[36]  (.D(z_next_reg[36]), .RN(n_0_231), .CK(n_0_217), .Q(z[36]), 
      .QN());
   DFFR_X1 \z_reg[35]  (.D(z_next_reg[35]), .RN(n_0_231), .CK(n_0_217), .Q(z[35]), 
      .QN());
   DFFR_X1 \z_reg[34]  (.D(z_next_reg[34]), .RN(n_0_231), .CK(n_0_217), .Q(z[34]), 
      .QN());
   DFFR_X1 \z_reg[33]  (.D(z_next_reg[33]), .RN(n_0_231), .CK(n_0_217), .Q(z[33]), 
      .QN());
   DFFR_X1 \z_reg[32]  (.D(z_next_reg[32]), .RN(n_0_231), .CK(n_0_217), .Q(z[32]), 
      .QN());
   DFFR_X1 \z_reg[31]  (.D(z_next_reg[31]), .RN(n_0_231), .CK(n_0_217), .Q(z[31]), 
      .QN());
   DFFR_X1 \z_reg[30]  (.D(z_next_reg[30]), .RN(n_0_231), .CK(n_0_217), .Q(z[30]), 
      .QN());
   DFFR_X1 \z_reg[29]  (.D(z_next_reg[29]), .RN(n_0_231), .CK(n_0_217), .Q(z[29]), 
      .QN());
   DFFR_X1 \z_reg[28]  (.D(z_next_reg[28]), .RN(n_0_231), .CK(n_0_217), .Q(z[28]), 
      .QN());
   DFFR_X1 \z_reg[27]  (.D(z_next_reg[27]), .RN(n_0_231), .CK(n_0_217), .Q(z[27]), 
      .QN());
   DFFR_X1 \z_reg[26]  (.D(z_next_reg[26]), .RN(n_0_231), .CK(n_0_217), .Q(z[26]), 
      .QN());
   DFFR_X1 \z_reg[25]  (.D(z_next_reg[25]), .RN(n_0_231), .CK(n_0_217), .Q(z[25]), 
      .QN());
   DFFR_X1 \z_reg[24]  (.D(z_next_reg[24]), .RN(n_0_231), .CK(n_0_217), .Q(z[24]), 
      .QN());
   DFFR_X1 \z_reg[23]  (.D(z_next_reg[23]), .RN(n_0_231), .CK(n_0_217), .Q(z[23]), 
      .QN());
   DFFR_X1 \z_reg[22]  (.D(z_next_reg[22]), .RN(n_0_231), .CK(n_0_217), .Q(z[22]), 
      .QN());
   DFFR_X1 \z_reg[21]  (.D(z_next_reg[21]), .RN(n_0_231), .CK(n_0_217), .Q(z[21]), 
      .QN());
   DFFR_X1 \z_reg[20]  (.D(z_next_reg[20]), .RN(n_0_231), .CK(n_0_217), .Q(z[20]), 
      .QN());
   DFFR_X1 \z_reg[19]  (.D(z_next_reg[19]), .RN(n_0_231), .CK(n_0_217), .Q(z[19]), 
      .QN());
   DFFR_X1 \z_reg[18]  (.D(z_next_reg[18]), .RN(n_0_231), .CK(n_0_217), .Q(z[18]), 
      .QN());
   DFFR_X1 \z_reg[17]  (.D(z_next_reg[17]), .RN(n_0_231), .CK(n_0_217), .Q(z[17]), 
      .QN());
   DFFR_X1 \z_reg[16]  (.D(z_next_reg[16]), .RN(n_0_231), .CK(n_0_217), .Q(z[16]), 
      .QN());
   DFFR_X1 \z_reg[15]  (.D(z_next_reg[15]), .RN(n_0_231), .CK(n_0_217), .Q(z[15]), 
      .QN());
   DFFR_X1 \z_reg[14]  (.D(z_next_reg[14]), .RN(n_0_231), .CK(n_0_217), .Q(z[14]), 
      .QN());
   DFFR_X1 \z_reg[13]  (.D(z_next_reg[13]), .RN(n_0_231), .CK(n_0_217), .Q(z[13]), 
      .QN());
   DFFR_X1 \z_reg[12]  (.D(z_next_reg[12]), .RN(n_0_231), .CK(n_0_217), .Q(z[12]), 
      .QN());
   DFFR_X1 \z_reg[11]  (.D(z_next_reg[11]), .RN(n_0_231), .CK(n_0_217), .Q(z[11]), 
      .QN());
   DFFR_X1 \z_reg[10]  (.D(z_next_reg[10]), .RN(n_0_231), .CK(n_0_217), .Q(z[10]), 
      .QN());
   DFFR_X1 \z_reg[9]  (.D(z_next_reg[9]), .RN(n_0_231), .CK(n_0_217), .Q(z[9]), 
      .QN());
   DFFR_X1 \z_reg[8]  (.D(z_next_reg[8]), .RN(n_0_231), .CK(n_0_217), .Q(z[8]), 
      .QN());
   DFFR_X1 \z_reg[7]  (.D(z_next_reg[7]), .RN(n_0_231), .CK(n_0_217), .Q(z[7]), 
      .QN());
   DFFR_X1 \z_reg[6]  (.D(z_next_reg[6]), .RN(n_0_231), .CK(n_0_217), .Q(z[6]), 
      .QN());
   DFFR_X1 \z_reg[5]  (.D(z_next_reg[5]), .RN(n_0_231), .CK(n_0_217), .Q(z[5]), 
      .QN());
   DFFR_X1 \z_reg[4]  (.D(z_next_reg[4]), .RN(n_0_231), .CK(n_0_217), .Q(z[4]), 
      .QN());
   DFFR_X1 \z_reg[3]  (.D(z_next_reg[3]), .RN(n_0_231), .CK(n_0_217), .Q(z[3]), 
      .QN());
   DFFR_X1 \z_reg[2]  (.D(z_next_reg[2]), .RN(n_0_231), .CK(n_0_217), .Q(z[2]), 
      .QN());
   DFFR_X1 \z_reg[1]  (.D(z_next_reg[1]), .RN(n_0_231), .CK(n_0_217), .Q(z[1]), 
      .QN());
   DFFR_X1 \z_reg[0]  (.D(z_next_reg[0]), .RN(n_0_231), .CK(n_0_217), .Q(z[0]), 
      .QN());
   datapath__0_162 i_0_22 (.plus({n_0_225, n_0_224, n_0_223, n_0_222, n_0_221, 
      n_0_220, n_0_219, n_0_218, n_0_216, n_0_215, n_0_214, n_0_213, n_0_212, 
      n_0_211, n_0_210, n_0_209, n_0_208, n_0_207, n_0_206, n_0_205, n_0_204, 
      n_0_203, n_0_202, n_0_201, n_0_200, n_0_199, n_0_198, n_0_197, n_0_196, 
      n_0_195, n_0_194, n_0_193, n_0_192, n_0_191, n_0_190, n_0_189, n_0_188, 
      n_0_187, n_0_186, n_0_185, n_0_184, n_0_183, n_0_182, n_0_181, n_0_180, 
      n_0_179, n_0_178, n_0_177, n_0_176, n_0_175, n_0_174, n_0_173, n_0_172, 
      n_0_171, n_0_170, n_0_169, n_0_168, n_0_167, n_0_166, n_0_165, n_0_164, 
      n_0_163, n_0_162, uc_16}), .quotient(quotient));
   DLH_X1 posv_sig_reg (.D(n_0_392), .G(n_0_391), .Q(posv_sig));
   DLH_X1 zero_sig_reg (.D(n_0_365), .G(n_0_391), .Q(zero_sig));
   DLH_X1 ovfl_sig_reg (.D(n_0_364), .G(n_0_391), .Q(ovfl_sig));
   DLH_X1 div_by_zero_sig_reg (.D(n_0_363), .G(n_0_391), .Q(div_by_zero_sig));
   DLH_X1 \out_sig_reg[63]  (.D(n_0_362), .G(n_0_391), .Q(out_sig[63]));
   DLH_X1 \out_sig_reg[62]  (.D(n_0_361), .G(n_0_391), .Q(out_sig[62]));
   DLH_X1 \out_sig_reg[61]  (.D(n_0_360), .G(n_0_391), .Q(out_sig[61]));
   DLH_X1 \out_sig_reg[60]  (.D(n_0_359), .G(n_0_391), .Q(out_sig[60]));
   DLH_X1 \out_sig_reg[59]  (.D(n_0_358), .G(n_0_391), .Q(out_sig[59]));
   DLH_X1 \out_sig_reg[58]  (.D(n_0_357), .G(n_0_391), .Q(out_sig[58]));
   DLH_X1 \out_sig_reg[57]  (.D(n_0_356), .G(n_0_391), .Q(out_sig[57]));
   DLH_X1 \out_sig_reg[56]  (.D(n_0_355), .G(n_0_391), .Q(out_sig[56]));
   DLH_X1 \out_sig_reg[55]  (.D(n_0_354), .G(n_0_391), .Q(out_sig[55]));
   DLH_X1 \out_sig_reg[54]  (.D(n_0_353), .G(n_0_391), .Q(out_sig[54]));
   DLH_X1 \out_sig_reg[53]  (.D(n_0_352), .G(n_0_391), .Q(out_sig[53]));
   DLH_X1 \out_sig_reg[52]  (.D(n_0_351), .G(n_0_391), .Q(out_sig[52]));
   DLH_X1 \out_sig_reg[51]  (.D(n_0_350), .G(n_0_391), .Q(out_sig[51]));
   DLH_X1 \out_sig_reg[50]  (.D(n_0_349), .G(n_0_391), .Q(out_sig[50]));
   DLH_X1 \out_sig_reg[49]  (.D(n_0_348), .G(n_0_391), .Q(out_sig[49]));
   DLH_X1 \out_sig_reg[48]  (.D(n_0_347), .G(n_0_391), .Q(out_sig[48]));
   DLH_X1 \out_sig_reg[47]  (.D(n_0_346), .G(n_0_391), .Q(out_sig[47]));
   DLH_X1 \out_sig_reg[46]  (.D(n_0_345), .G(n_0_391), .Q(out_sig[46]));
   DLH_X1 \out_sig_reg[45]  (.D(n_0_344), .G(n_0_391), .Q(out_sig[45]));
   DLH_X1 \out_sig_reg[44]  (.D(n_0_343), .G(n_0_391), .Q(out_sig[44]));
   DLH_X1 \out_sig_reg[43]  (.D(n_0_342), .G(n_0_391), .Q(out_sig[43]));
   DLH_X1 \out_sig_reg[42]  (.D(n_0_341), .G(n_0_391), .Q(out_sig[42]));
   DLH_X1 \out_sig_reg[41]  (.D(n_0_340), .G(n_0_391), .Q(out_sig[41]));
   DLH_X1 \out_sig_reg[40]  (.D(n_0_339), .G(n_0_391), .Q(out_sig[40]));
   DLH_X1 \out_sig_reg[39]  (.D(n_0_338), .G(n_0_391), .Q(out_sig[39]));
   DLH_X1 \out_sig_reg[38]  (.D(n_0_337), .G(n_0_391), .Q(out_sig[38]));
   DLH_X1 \out_sig_reg[37]  (.D(n_0_336), .G(n_0_391), .Q(out_sig[37]));
   DLH_X1 \out_sig_reg[36]  (.D(n_0_335), .G(n_0_391), .Q(out_sig[36]));
   DLH_X1 \out_sig_reg[35]  (.D(n_0_334), .G(n_0_391), .Q(out_sig[35]));
   DLH_X1 \out_sig_reg[34]  (.D(n_0_333), .G(n_0_391), .Q(out_sig[34]));
   DLH_X1 \out_sig_reg[33]  (.D(n_0_332), .G(n_0_391), .Q(out_sig[33]));
   DLH_X1 \out_sig_reg[32]  (.D(n_0_331), .G(n_0_391), .Q(out_sig[32]));
   DLH_X1 \out_sig_reg[31]  (.D(n_0_330), .G(n_0_391), .Q(out_sig[31]));
   DLH_X1 \out_sig_reg[30]  (.D(n_0_329), .G(n_0_391), .Q(out_sig[30]));
   DLH_X1 \out_sig_reg[29]  (.D(n_0_328), .G(n_0_391), .Q(out_sig[29]));
   DLH_X1 \out_sig_reg[28]  (.D(n_0_327), .G(n_0_391), .Q(out_sig[28]));
   DLH_X1 \out_sig_reg[27]  (.D(n_0_326), .G(n_0_391), .Q(out_sig[27]));
   DLH_X1 \out_sig_reg[26]  (.D(n_0_325), .G(n_0_391), .Q(out_sig[26]));
   DLH_X1 \out_sig_reg[25]  (.D(n_0_324), .G(n_0_391), .Q(out_sig[25]));
   DLH_X1 \out_sig_reg[24]  (.D(n_0_323), .G(n_0_391), .Q(out_sig[24]));
   DLH_X1 \out_sig_reg[23]  (.D(n_0_322), .G(n_0_391), .Q(out_sig[23]));
   DLH_X1 \out_sig_reg[22]  (.D(n_0_321), .G(n_0_391), .Q(out_sig[22]));
   DLH_X1 \out_sig_reg[21]  (.D(n_0_320), .G(n_0_391), .Q(out_sig[21]));
   DLH_X1 \out_sig_reg[20]  (.D(n_0_319), .G(n_0_391), .Q(out_sig[20]));
   DLH_X1 \out_sig_reg[19]  (.D(n_0_318), .G(n_0_391), .Q(out_sig[19]));
   DLH_X1 \out_sig_reg[18]  (.D(n_0_317), .G(n_0_391), .Q(out_sig[18]));
   DLH_X1 \out_sig_reg[17]  (.D(n_0_316), .G(n_0_391), .Q(out_sig[17]));
   DLH_X1 \out_sig_reg[16]  (.D(n_0_315), .G(n_0_391), .Q(out_sig[16]));
   DLH_X1 \out_sig_reg[15]  (.D(n_0_314), .G(n_0_391), .Q(out_sig[15]));
   DLH_X1 \out_sig_reg[14]  (.D(n_0_313), .G(n_0_391), .Q(out_sig[14]));
   DLH_X1 \out_sig_reg[13]  (.D(n_0_312), .G(n_0_391), .Q(out_sig[13]));
   DLH_X1 \out_sig_reg[12]  (.D(n_0_311), .G(n_0_391), .Q(out_sig[12]));
   DLH_X1 \out_sig_reg[11]  (.D(n_0_310), .G(n_0_391), .Q(out_sig[11]));
   DLH_X1 \out_sig_reg[10]  (.D(n_0_309), .G(n_0_391), .Q(out_sig[10]));
   DLH_X1 \out_sig_reg[9]  (.D(n_0_308), .G(n_0_391), .Q(out_sig[9]));
   DLH_X1 \out_sig_reg[8]  (.D(n_0_307), .G(n_0_391), .Q(out_sig[8]));
   DLH_X1 \out_sig_reg[7]  (.D(n_0_306), .G(n_0_391), .Q(out_sig[7]));
   DLH_X1 \out_sig_reg[6]  (.D(n_0_305), .G(n_0_391), .Q(out_sig[6]));
   DLH_X1 \out_sig_reg[5]  (.D(n_0_304), .G(n_0_391), .Q(out_sig[5]));
   DLH_X1 \out_sig_reg[4]  (.D(n_0_303), .G(n_0_391), .Q(out_sig[4]));
   DLH_X1 \out_sig_reg[3]  (.D(n_0_302), .G(n_0_391), .Q(out_sig[3]));
   DLH_X1 \out_sig_reg[2]  (.D(n_0_301), .G(n_0_391), .Q(out_sig[2]));
   DLH_X1 \out_sig_reg[1]  (.D(n_0_300), .G(n_0_391), .Q(out_sig[1]));
   DLH_X1 \out_sig_reg[0]  (.D(n_0_299), .G(n_0_391), .Q(out_sig[0]));
   DLH_X1 done_sig_reg (.D(n_0_298), .G(n_0_391), .Q(done_sig));
   datapath__0_153 i_0_41 (.p_0({n_0_390, n_0_389, n_0_388, n_0_387, n_0_386, 
      n_0_385, n_0_384, n_0_383, n_0_382, n_0_381, n_0_380, n_0_379, n_0_378, 
      n_0_377, n_0_376, n_0_375, n_0_374, n_0_373, n_0_372, n_0_371, n_0_370, 
      n_0_369, n_0_368, n_0_367, n_0_366, n_0_230, n_0_229, n_0_228, uc_17, 
      n_0_227, n_0_226, uc_18}), .i({i[31], i[30], i[29], i[28], i[27], i[26], 
      i[25], i[24], i[23], i[22], i[21], i[20], i[19], i[18], i[17], i[16], 
      i[15], i[14], i[13], i[12], i[11], i[10], i[9], i[8], i[7], i[6], i[5], 
      i[4], i[3], i[2], i[1], uc_19}));
   DLH_X1 \quotient_reg[63]  (.D(n_0_296), .G(n_0_295), .Q(quotient[63]));
   DLH_X1 \quotient_reg[62]  (.D(n_0_296), .G(n_0_294), .Q(quotient[62]));
   DLH_X1 \quotient_reg[61]  (.D(n_0_296), .G(n_0_293), .Q(quotient[61]));
   DLH_X1 \quotient_reg[60]  (.D(n_0_296), .G(n_0_292), .Q(quotient[60]));
   DLH_X1 \quotient_reg[59]  (.D(n_0_296), .G(n_0_291), .Q(quotient[59]));
   DLH_X1 \quotient_reg[58]  (.D(n_0_296), .G(n_0_290), .Q(quotient[58]));
   DLH_X1 \quotient_reg[57]  (.D(n_0_296), .G(n_0_289), .Q(quotient[57]));
   DLH_X1 \quotient_reg[56]  (.D(n_0_296), .G(n_0_288), .Q(quotient[56]));
   DLH_X1 \quotient_reg[55]  (.D(n_0_296), .G(n_0_287), .Q(quotient[55]));
   DLH_X1 \quotient_reg[54]  (.D(n_0_296), .G(n_0_286), .Q(quotient[54]));
   DLH_X1 \quotient_reg[53]  (.D(n_0_296), .G(n_0_285), .Q(quotient[53]));
   DLH_X1 \quotient_reg[52]  (.D(n_0_296), .G(n_0_284), .Q(quotient[52]));
   DLH_X1 \quotient_reg[51]  (.D(n_0_296), .G(n_0_283), .Q(quotient[51]));
   DLH_X1 \quotient_reg[50]  (.D(n_0_296), .G(n_0_282), .Q(quotient[50]));
   DLH_X1 \quotient_reg[49]  (.D(n_0_296), .G(n_0_281), .Q(quotient[49]));
   DLH_X1 \quotient_reg[48]  (.D(n_0_296), .G(n_0_280), .Q(quotient[48]));
   DLH_X1 \quotient_reg[47]  (.D(n_0_296), .G(n_0_279), .Q(quotient[47]));
   DLH_X1 \quotient_reg[46]  (.D(n_0_296), .G(n_0_278), .Q(quotient[46]));
   DLH_X1 \quotient_reg[45]  (.D(n_0_296), .G(n_0_277), .Q(quotient[45]));
   DLH_X1 \quotient_reg[44]  (.D(n_0_296), .G(n_0_276), .Q(quotient[44]));
   DLH_X1 \quotient_reg[43]  (.D(n_0_296), .G(n_0_275), .Q(quotient[43]));
   DLH_X1 \quotient_reg[42]  (.D(n_0_296), .G(n_0_274), .Q(quotient[42]));
   DLH_X1 \quotient_reg[41]  (.D(n_0_296), .G(n_0_273), .Q(quotient[41]));
   DLH_X1 \quotient_reg[40]  (.D(n_0_296), .G(n_0_272), .Q(quotient[40]));
   DLH_X1 \quotient_reg[39]  (.D(n_0_296), .G(n_0_271), .Q(quotient[39]));
   DLH_X1 \quotient_reg[38]  (.D(n_0_296), .G(n_0_270), .Q(quotient[38]));
   DLH_X1 \quotient_reg[37]  (.D(n_0_296), .G(n_0_269), .Q(quotient[37]));
   DLH_X1 \quotient_reg[36]  (.D(n_0_296), .G(n_0_268), .Q(quotient[36]));
   DLH_X1 \quotient_reg[35]  (.D(n_0_296), .G(n_0_267), .Q(quotient[35]));
   DLH_X1 \quotient_reg[34]  (.D(n_0_296), .G(n_0_266), .Q(quotient[34]));
   DLH_X1 \quotient_reg[33]  (.D(n_0_296), .G(n_0_265), .Q(quotient[33]));
   DLH_X1 \quotient_reg[32]  (.D(n_0_296), .G(n_0_264), .Q(quotient[32]));
   DLH_X1 \quotient_reg[31]  (.D(n_0_296), .G(n_0_263), .Q(quotient[31]));
   DLH_X1 \quotient_reg[30]  (.D(n_0_296), .G(n_0_262), .Q(quotient[30]));
   DLH_X1 \quotient_reg[29]  (.D(n_0_296), .G(n_0_261), .Q(quotient[29]));
   DLH_X1 \quotient_reg[28]  (.D(n_0_296), .G(n_0_260), .Q(quotient[28]));
   DLH_X1 \quotient_reg[27]  (.D(n_0_296), .G(n_0_259), .Q(quotient[27]));
   DLH_X1 \quotient_reg[26]  (.D(n_0_296), .G(n_0_258), .Q(quotient[26]));
   DLH_X1 \quotient_reg[25]  (.D(n_0_296), .G(n_0_257), .Q(quotient[25]));
   DLH_X1 \quotient_reg[24]  (.D(n_0_296), .G(n_0_256), .Q(quotient[24]));
   DLH_X1 \quotient_reg[23]  (.D(n_0_296), .G(n_0_255), .Q(quotient[23]));
   DLH_X1 \quotient_reg[22]  (.D(n_0_296), .G(n_0_254), .Q(quotient[22]));
   DLH_X1 \quotient_reg[21]  (.D(n_0_296), .G(n_0_253), .Q(quotient[21]));
   DLH_X1 \quotient_reg[20]  (.D(n_0_296), .G(n_0_252), .Q(quotient[20]));
   DLH_X1 \quotient_reg[19]  (.D(n_0_296), .G(n_0_251), .Q(quotient[19]));
   DLH_X1 \quotient_reg[18]  (.D(n_0_296), .G(n_0_250), .Q(quotient[18]));
   DLH_X1 \quotient_reg[17]  (.D(n_0_296), .G(n_0_249), .Q(quotient[17]));
   DLH_X1 \quotient_reg[16]  (.D(n_0_296), .G(n_0_248), .Q(quotient[16]));
   DLH_X1 \quotient_reg[15]  (.D(n_0_296), .G(n_0_247), .Q(quotient[15]));
   DLH_X1 \quotient_reg[14]  (.D(n_0_296), .G(n_0_246), .Q(quotient[14]));
   DLH_X1 \quotient_reg[13]  (.D(n_0_296), .G(n_0_245), .Q(quotient[13]));
   DLH_X1 \quotient_reg[12]  (.D(n_0_296), .G(n_0_244), .Q(quotient[12]));
   DLH_X1 \quotient_reg[11]  (.D(n_0_296), .G(n_0_243), .Q(quotient[11]));
   DLH_X1 \quotient_reg[10]  (.D(n_0_296), .G(n_0_242), .Q(quotient[10]));
   DLH_X1 \quotient_reg[9]  (.D(n_0_296), .G(n_0_241), .Q(quotient[9]));
   DLH_X1 \quotient_reg[8]  (.D(n_0_296), .G(n_0_240), .Q(quotient[8]));
   DLH_X1 \quotient_reg[7]  (.D(n_0_296), .G(n_0_239), .Q(quotient[7]));
   DLH_X1 \quotient_reg[6]  (.D(n_0_296), .G(n_0_238), .Q(quotient[6]));
   DLH_X1 \quotient_reg[5]  (.D(n_0_296), .G(n_0_237), .Q(quotient[5]));
   DLH_X1 \quotient_reg[4]  (.D(n_0_296), .G(n_0_236), .Q(quotient[4]));
   DLH_X1 \quotient_reg[3]  (.D(n_0_296), .G(n_0_235), .Q(quotient[3]));
   DLH_X1 \quotient_reg[2]  (.D(n_0_296), .G(n_0_234), .Q(quotient[2]));
   DLH_X1 \quotient_reg[1]  (.D(n_0_296), .G(n_0_233), .Q(quotient[1]));
   DLH_X1 \quotient_reg[0]  (.D(n_0_296), .G(n_0_232), .Q(quotient[0]));
   datapath__0_158 i_0_45 (.p_0({n_0_390, n_0_389, n_0_388, n_0_387, n_0_386, 
      n_0_385, n_0_384, n_0_383, n_0_382, n_0_381, n_0_380, n_0_379, n_0_378, 
      n_0_377, n_0_376, n_0_375, n_0_374, n_0_373, n_0_372, n_0_371, n_0_370, 
      n_0_369, n_0_368, n_0_367, n_0_366, n_0_230, n_0_229, n_0_228, i[3], 
      n_0_227, n_0_226, n_0_130}), .p_1({n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, 
      n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, n_0_0, n_0_412, n_0_411, n_0_410, 
      n_0_409, n_0_408, n_0_407, n_0_406, n_0_405, n_0_404, n_0_403, n_0_402, 
      n_0_401, n_0_400, n_0_399, n_0_398, n_0_397, n_0_396, n_0_395, n_0_394, 
      n_0_393, uc_20}));
   INV_X1 i_0_1_0 (.A(rst), .ZN(n_0_231));
   NOR2_X1 i_0_2_0 (.A1(state[0]), .A2(state[1]), .ZN(n_0_2_0));
   INV_X1 i_0_2_1 (.A(n_0_2_0), .ZN(n_0_298));
   NOR4_X1 i_0_2_2 (.A1(n_0_4), .A2(n_0_3), .A3(n_0_2), .A4(n_0_1), .ZN(n_0_2_1));
   NOR4_X1 i_0_2_3 (.A1(n_0_8), .A2(n_0_7), .A3(n_0_6), .A4(n_0_5), .ZN(n_0_2_2));
   NOR4_X1 i_0_2_4 (.A1(n_0_0), .A2(n_0_412), .A3(n_0_411), .A4(n_0_410), 
      .ZN(n_0_2_3));
   NOR2_X1 i_0_2_5 (.A1(n_0_10), .A2(n_0_9), .ZN(n_0_2_4));
   AND4_X1 i_0_2_6 (.A1(n_0_2_1), .A2(n_0_2_2), .A3(n_0_2_3), .A4(n_0_2_4), 
      .ZN(n_0_2_5));
   NOR4_X1 i_0_2_7 (.A1(n_0_405), .A2(n_0_404), .A3(n_0_403), .A4(n_0_402), 
      .ZN(n_0_2_6));
   NOR4_X1 i_0_2_8 (.A1(n_0_409), .A2(n_0_408), .A3(n_0_407), .A4(n_0_406), 
      .ZN(n_0_2_7));
   NOR4_X1 i_0_2_9 (.A1(n_0_401), .A2(n_0_400), .A3(n_0_399), .A4(n_0_398), 
      .ZN(n_0_2_8));
   AND4_X1 i_0_2_10 (.A1(n_0_2_5), .A2(n_0_2_6), .A3(n_0_2_7), .A4(n_0_2_8), 
      .ZN(n_0_2_9));
   INV_X1 i_0_2_11 (.A(n_0_396), .ZN(n_0_2_10));
   NAND2_X1 i_0_2_12 (.A1(n_0_2_9), .A2(n_0_2_10), .ZN(n_0_2_11));
   NOR2_X1 i_0_2_13 (.A1(n_0_2_11), .A2(n_0_395), .ZN(n_0_2_12));
   INV_X1 i_0_2_14 (.A(n_0_397), .ZN(n_0_2_13));
   NAND2_X1 i_0_2_15 (.A1(n_0_2_12), .A2(n_0_2_13), .ZN(n_0_2_14));
   INV_X1 i_0_2_16 (.A(state[1]), .ZN(n_0_2_15));
   NOR2_X1 i_0_2_17 (.A1(n_0_2_15), .A2(n_0_393), .ZN(n_0_2_16));
   INV_X1 i_0_2_18 (.A(n_0_394), .ZN(n_0_2_17));
   NAND3_X1 i_0_2_19 (.A1(n_0_2_16), .A2(n_0_2_17), .A3(n_0_130), .ZN(n_0_2_18));
   OAI21_X1 i_0_2_20 (.A(n_0_298), .B1(n_0_2_14), .B2(n_0_2_18), .ZN(n_0_232));
   NAND3_X1 i_0_2_21 (.A1(n_0_2_16), .A2(n_0_2_17), .A3(i[0]), .ZN(n_0_2_19));
   OAI21_X1 i_0_2_22 (.A(n_0_298), .B1(n_0_2_14), .B2(n_0_2_19), .ZN(n_0_233));
   AND2_X1 i_0_2_23 (.A1(n_0_393), .A2(state[1]), .ZN(n_0_2_20));
   NAND3_X1 i_0_2_24 (.A1(n_0_2_20), .A2(n_0_2_17), .A3(n_0_130), .ZN(n_0_2_21));
   OAI21_X1 i_0_2_25 (.A(n_0_298), .B1(n_0_2_14), .B2(n_0_2_21), .ZN(n_0_234));
   NAND3_X1 i_0_2_26 (.A1(n_0_2_20), .A2(n_0_2_17), .A3(i[0]), .ZN(n_0_2_22));
   OAI21_X1 i_0_2_27 (.A(n_0_298), .B1(n_0_2_14), .B2(n_0_2_22), .ZN(n_0_235));
   NAND3_X1 i_0_2_28 (.A1(n_0_2_16), .A2(n_0_394), .A3(n_0_130), .ZN(n_0_2_23));
   OAI21_X1 i_0_2_29 (.A(n_0_298), .B1(n_0_2_14), .B2(n_0_2_23), .ZN(n_0_236));
   NAND3_X1 i_0_2_30 (.A1(n_0_2_16), .A2(n_0_394), .A3(i[0]), .ZN(n_0_2_24));
   OAI21_X1 i_0_2_31 (.A(n_0_298), .B1(n_0_2_14), .B2(n_0_2_24), .ZN(n_0_237));
   NAND3_X1 i_0_2_32 (.A1(n_0_2_20), .A2(n_0_394), .A3(n_0_130), .ZN(n_0_2_25));
   OAI21_X1 i_0_2_33 (.A(n_0_298), .B1(n_0_2_14), .B2(n_0_2_25), .ZN(n_0_238));
   NAND3_X1 i_0_2_34 (.A1(n_0_2_20), .A2(n_0_394), .A3(i[0]), .ZN(n_0_2_26));
   OAI21_X1 i_0_2_35 (.A(n_0_298), .B1(n_0_2_14), .B2(n_0_2_26), .ZN(n_0_239));
   INV_X1 i_0_2_36 (.A(n_0_395), .ZN(n_0_2_27));
   NOR2_X1 i_0_2_37 (.A1(n_0_2_11), .A2(n_0_2_27), .ZN(n_0_2_28));
   NAND2_X1 i_0_2_38 (.A1(n_0_2_28), .A2(n_0_2_13), .ZN(n_0_2_29));
   OAI21_X1 i_0_2_39 (.A(n_0_298), .B1(n_0_2_29), .B2(n_0_2_18), .ZN(n_0_240));
   OAI21_X1 i_0_2_40 (.A(n_0_298), .B1(n_0_2_29), .B2(n_0_2_19), .ZN(n_0_241));
   OAI21_X1 i_0_2_41 (.A(n_0_298), .B1(n_0_2_29), .B2(n_0_2_21), .ZN(n_0_242));
   OAI21_X1 i_0_2_42 (.A(n_0_298), .B1(n_0_2_29), .B2(n_0_2_22), .ZN(n_0_243));
   OAI21_X1 i_0_2_43 (.A(n_0_298), .B1(n_0_2_29), .B2(n_0_2_23), .ZN(n_0_244));
   OAI21_X1 i_0_2_44 (.A(n_0_298), .B1(n_0_2_29), .B2(n_0_2_24), .ZN(n_0_245));
   OAI21_X1 i_0_2_45 (.A(n_0_298), .B1(n_0_2_29), .B2(n_0_2_25), .ZN(n_0_246));
   OAI21_X1 i_0_2_46 (.A(n_0_298), .B1(n_0_2_29), .B2(n_0_2_26), .ZN(n_0_247));
   NAND2_X1 i_0_2_47 (.A1(n_0_2_9), .A2(n_0_396), .ZN(n_0_2_30));
   NOR2_X1 i_0_2_48 (.A1(n_0_2_30), .A2(n_0_395), .ZN(n_0_2_31));
   NAND2_X1 i_0_2_49 (.A1(n_0_2_31), .A2(n_0_2_13), .ZN(n_0_2_32));
   OAI21_X1 i_0_2_50 (.A(n_0_298), .B1(n_0_2_32), .B2(n_0_2_18), .ZN(n_0_248));
   OAI21_X1 i_0_2_51 (.A(n_0_298), .B1(n_0_2_32), .B2(n_0_2_19), .ZN(n_0_249));
   OAI21_X1 i_0_2_52 (.A(n_0_298), .B1(n_0_2_32), .B2(n_0_2_21), .ZN(n_0_250));
   OAI21_X1 i_0_2_53 (.A(n_0_298), .B1(n_0_2_32), .B2(n_0_2_22), .ZN(n_0_251));
   OAI21_X1 i_0_2_54 (.A(n_0_298), .B1(n_0_2_32), .B2(n_0_2_23), .ZN(n_0_252));
   OAI21_X1 i_0_2_55 (.A(n_0_298), .B1(n_0_2_32), .B2(n_0_2_24), .ZN(n_0_253));
   OAI21_X1 i_0_2_56 (.A(n_0_298), .B1(n_0_2_32), .B2(n_0_2_25), .ZN(n_0_254));
   OAI21_X1 i_0_2_57 (.A(n_0_298), .B1(n_0_2_32), .B2(n_0_2_26), .ZN(n_0_255));
   NOR2_X1 i_0_2_58 (.A1(n_0_2_30), .A2(n_0_2_27), .ZN(n_0_2_33));
   NAND2_X1 i_0_2_59 (.A1(n_0_2_33), .A2(n_0_2_13), .ZN(n_0_2_34));
   OAI21_X1 i_0_2_60 (.A(n_0_298), .B1(n_0_2_34), .B2(n_0_2_18), .ZN(n_0_256));
   OAI21_X1 i_0_2_61 (.A(n_0_298), .B1(n_0_2_34), .B2(n_0_2_19), .ZN(n_0_257));
   OAI21_X1 i_0_2_62 (.A(n_0_298), .B1(n_0_2_34), .B2(n_0_2_21), .ZN(n_0_258));
   OAI21_X1 i_0_2_63 (.A(n_0_298), .B1(n_0_2_34), .B2(n_0_2_22), .ZN(n_0_259));
   OAI21_X1 i_0_2_64 (.A(n_0_298), .B1(n_0_2_34), .B2(n_0_2_23), .ZN(n_0_260));
   OAI21_X1 i_0_2_65 (.A(n_0_298), .B1(n_0_2_34), .B2(n_0_2_24), .ZN(n_0_261));
   OAI21_X1 i_0_2_66 (.A(n_0_298), .B1(n_0_2_34), .B2(n_0_2_25), .ZN(n_0_262));
   OAI21_X1 i_0_2_67 (.A(n_0_298), .B1(n_0_2_34), .B2(n_0_2_26), .ZN(n_0_263));
   NAND2_X1 i_0_2_68 (.A1(n_0_2_12), .A2(n_0_397), .ZN(n_0_2_35));
   OAI21_X1 i_0_2_69 (.A(n_0_298), .B1(n_0_2_35), .B2(n_0_2_18), .ZN(n_0_264));
   OAI21_X1 i_0_2_70 (.A(n_0_298), .B1(n_0_2_35), .B2(n_0_2_19), .ZN(n_0_265));
   OAI21_X1 i_0_2_71 (.A(n_0_298), .B1(n_0_2_35), .B2(n_0_2_21), .ZN(n_0_266));
   OAI21_X1 i_0_2_72 (.A(n_0_298), .B1(n_0_2_35), .B2(n_0_2_22), .ZN(n_0_267));
   OAI21_X1 i_0_2_73 (.A(n_0_298), .B1(n_0_2_35), .B2(n_0_2_23), .ZN(n_0_268));
   OAI21_X1 i_0_2_74 (.A(n_0_298), .B1(n_0_2_35), .B2(n_0_2_24), .ZN(n_0_269));
   OAI21_X1 i_0_2_75 (.A(n_0_298), .B1(n_0_2_35), .B2(n_0_2_25), .ZN(n_0_270));
   OAI21_X1 i_0_2_76 (.A(n_0_298), .B1(n_0_2_35), .B2(n_0_2_26), .ZN(n_0_271));
   NAND2_X1 i_0_2_77 (.A1(n_0_2_28), .A2(n_0_397), .ZN(n_0_2_36));
   OAI21_X1 i_0_2_78 (.A(n_0_298), .B1(n_0_2_36), .B2(n_0_2_18), .ZN(n_0_272));
   OAI21_X1 i_0_2_79 (.A(n_0_298), .B1(n_0_2_36), .B2(n_0_2_19), .ZN(n_0_273));
   OAI21_X1 i_0_2_80 (.A(n_0_298), .B1(n_0_2_36), .B2(n_0_2_21), .ZN(n_0_274));
   OAI21_X1 i_0_2_81 (.A(n_0_298), .B1(n_0_2_36), .B2(n_0_2_22), .ZN(n_0_275));
   OAI21_X1 i_0_2_82 (.A(n_0_298), .B1(n_0_2_36), .B2(n_0_2_23), .ZN(n_0_276));
   OAI21_X1 i_0_2_83 (.A(n_0_298), .B1(n_0_2_36), .B2(n_0_2_24), .ZN(n_0_277));
   OAI21_X1 i_0_2_84 (.A(n_0_298), .B1(n_0_2_36), .B2(n_0_2_25), .ZN(n_0_278));
   OAI21_X1 i_0_2_85 (.A(n_0_298), .B1(n_0_2_36), .B2(n_0_2_26), .ZN(n_0_279));
   NAND2_X1 i_0_2_86 (.A1(n_0_2_31), .A2(n_0_397), .ZN(n_0_2_37));
   OAI21_X1 i_0_2_87 (.A(n_0_298), .B1(n_0_2_37), .B2(n_0_2_18), .ZN(n_0_280));
   OAI21_X1 i_0_2_88 (.A(n_0_298), .B1(n_0_2_37), .B2(n_0_2_19), .ZN(n_0_281));
   OAI21_X1 i_0_2_89 (.A(n_0_298), .B1(n_0_2_37), .B2(n_0_2_21), .ZN(n_0_282));
   OAI21_X1 i_0_2_90 (.A(n_0_298), .B1(n_0_2_37), .B2(n_0_2_22), .ZN(n_0_283));
   OAI21_X1 i_0_2_91 (.A(n_0_298), .B1(n_0_2_37), .B2(n_0_2_23), .ZN(n_0_284));
   OAI21_X1 i_0_2_92 (.A(n_0_298), .B1(n_0_2_37), .B2(n_0_2_24), .ZN(n_0_285));
   OAI21_X1 i_0_2_93 (.A(n_0_298), .B1(n_0_2_37), .B2(n_0_2_25), .ZN(n_0_286));
   OAI21_X1 i_0_2_94 (.A(n_0_298), .B1(n_0_2_37), .B2(n_0_2_26), .ZN(n_0_287));
   NAND2_X1 i_0_2_95 (.A1(n_0_2_33), .A2(n_0_397), .ZN(n_0_2_38));
   OAI21_X1 i_0_2_96 (.A(n_0_298), .B1(n_0_2_38), .B2(n_0_2_18), .ZN(n_0_288));
   OAI21_X1 i_0_2_97 (.A(n_0_298), .B1(n_0_2_38), .B2(n_0_2_19), .ZN(n_0_289));
   OAI21_X1 i_0_2_98 (.A(n_0_298), .B1(n_0_2_38), .B2(n_0_2_21), .ZN(n_0_290));
   OAI21_X1 i_0_2_99 (.A(n_0_298), .B1(n_0_2_38), .B2(n_0_2_22), .ZN(n_0_291));
   OAI21_X1 i_0_2_100 (.A(n_0_298), .B1(n_0_2_38), .B2(n_0_2_23), .ZN(n_0_292));
   OAI21_X1 i_0_2_101 (.A(n_0_298), .B1(n_0_2_38), .B2(n_0_2_24), .ZN(n_0_293));
   OAI21_X1 i_0_2_102 (.A(n_0_298), .B1(n_0_2_38), .B2(n_0_2_25), .ZN(n_0_294));
   OAI21_X1 i_0_2_103 (.A(n_0_298), .B1(n_0_2_38), .B2(n_0_2_26), .ZN(n_0_295));
   INV_X1 i_0_2_104 (.A(in_b[63]), .ZN(n_0_2_39));
   OAI22_X1 i_0_2_105 (.A1(n_0_2_39), .A2(n_0_11), .B1(in_b[63]), .B2(in_b[1]), 
      .ZN(n_0_2_40));
   INV_X1 i_0_2_106 (.A(n_0_2_40), .ZN(b[1]));
   AOI22_X1 i_0_2_107 (.A1(n_0_2_39), .A2(in_b[3]), .B1(n_0_13), .B2(in_b[63]), 
      .ZN(n_0_2_41));
   INV_X1 i_0_2_108 (.A(n_0_2_41), .ZN(b[3]));
   AOI22_X1 i_0_2_109 (.A1(n_0_2_39), .A2(in_b[2]), .B1(n_0_12), .B2(in_b[63]), 
      .ZN(n_0_2_42));
   INV_X1 i_0_2_110 (.A(n_0_2_42), .ZN(b[2]));
   AOI22_X1 i_0_2_111 (.A1(n_0_2_39), .A2(in_b[4]), .B1(n_0_14), .B2(in_b[63]), 
      .ZN(n_0_2_43));
   INV_X1 i_0_2_112 (.A(n_0_2_43), .ZN(b[4]));
   AOI22_X1 i_0_2_113 (.A1(n_0_2_39), .A2(in_b[6]), .B1(n_0_16), .B2(in_b[63]), 
      .ZN(n_0_2_44));
   INV_X1 i_0_2_114 (.A(n_0_2_44), .ZN(b[6]));
   OAI22_X1 i_0_2_115 (.A1(n_0_2_39), .A2(n_0_15), .B1(in_b[63]), .B2(in_b[5]), 
      .ZN(n_0_2_45));
   INV_X1 i_0_2_116 (.A(n_0_2_45), .ZN(b[5]));
   AOI22_X1 i_0_2_117 (.A1(n_0_2_39), .A2(in_b[8]), .B1(n_0_18), .B2(in_b[63]), 
      .ZN(n_0_2_46));
   INV_X1 i_0_2_118 (.A(n_0_2_46), .ZN(b[8]));
   OAI22_X1 i_0_2_119 (.A1(n_0_2_39), .A2(n_0_17), .B1(in_b[63]), .B2(in_b[7]), 
      .ZN(n_0_2_47));
   INV_X1 i_0_2_120 (.A(n_0_2_47), .ZN(b[7]));
   AOI22_X1 i_0_2_121 (.A1(n_0_2_39), .A2(in_b[10]), .B1(n_0_20), .B2(in_b[63]), 
      .ZN(n_0_2_48));
   INV_X1 i_0_2_122 (.A(n_0_2_48), .ZN(b[10]));
   AOI22_X1 i_0_2_123 (.A1(n_0_2_39), .A2(in_b[9]), .B1(n_0_19), .B2(in_b[63]), 
      .ZN(n_0_2_49));
   INV_X1 i_0_2_124 (.A(n_0_2_49), .ZN(b[9]));
   AOI22_X1 i_0_2_125 (.A1(n_0_2_39), .A2(in_b[11]), .B1(n_0_21), .B2(in_b[63]), 
      .ZN(n_0_2_50));
   INV_X1 i_0_2_126 (.A(n_0_2_50), .ZN(b[11]));
   AOI22_X1 i_0_2_127 (.A1(n_0_2_39), .A2(in_b[12]), .B1(n_0_22), .B2(in_b[63]), 
      .ZN(n_0_2_51));
   INV_X1 i_0_2_128 (.A(n_0_2_51), .ZN(b[12]));
   OAI22_X1 i_0_2_129 (.A1(n_0_2_39), .A2(n_0_23), .B1(in_b[63]), .B2(in_b[13]), 
      .ZN(n_0_2_52));
   INV_X1 i_0_2_130 (.A(n_0_2_52), .ZN(b[13]));
   AOI22_X1 i_0_2_131 (.A1(n_0_2_39), .A2(in_b[14]), .B1(n_0_24), .B2(in_b[63]), 
      .ZN(n_0_2_53));
   INV_X1 i_0_2_132 (.A(n_0_2_53), .ZN(b[14]));
   AOI22_X1 i_0_2_133 (.A1(n_0_2_39), .A2(in_b[16]), .B1(n_0_26), .B2(in_b[63]), 
      .ZN(n_0_2_54));
   INV_X1 i_0_2_134 (.A(n_0_2_54), .ZN(b[16]));
   AOI22_X1 i_0_2_135 (.A1(n_0_2_39), .A2(in_b[15]), .B1(n_0_25), .B2(in_b[63]), 
      .ZN(n_0_2_55));
   INV_X1 i_0_2_136 (.A(n_0_2_55), .ZN(b[15]));
   OAI22_X1 i_0_2_137 (.A1(n_0_2_39), .A2(n_0_27), .B1(in_b[63]), .B2(in_b[17]), 
      .ZN(n_0_2_56));
   INV_X1 i_0_2_138 (.A(n_0_2_56), .ZN(b[17]));
   AOI22_X1 i_0_2_139 (.A1(n_0_2_39), .A2(in_b[18]), .B1(n_0_28), .B2(in_b[63]), 
      .ZN(n_0_2_57));
   INV_X1 i_0_2_140 (.A(n_0_2_57), .ZN(b[18]));
   AOI22_X1 i_0_2_141 (.A1(n_0_2_39), .A2(in_b[20]), .B1(n_0_30), .B2(in_b[63]), 
      .ZN(n_0_2_58));
   INV_X1 i_0_2_142 (.A(n_0_2_58), .ZN(b[20]));
   AOI22_X1 i_0_2_143 (.A1(n_0_2_39), .A2(in_b[19]), .B1(n_0_29), .B2(in_b[63]), 
      .ZN(n_0_2_59));
   INV_X1 i_0_2_144 (.A(n_0_2_59), .ZN(b[19]));
   AOI22_X1 i_0_2_145 (.A1(n_0_2_39), .A2(in_b[21]), .B1(n_0_31), .B2(in_b[63]), 
      .ZN(n_0_2_60));
   INV_X1 i_0_2_146 (.A(n_0_2_60), .ZN(b[21]));
   AOI22_X1 i_0_2_147 (.A1(n_0_2_39), .A2(in_b[22]), .B1(n_0_32), .B2(in_b[63]), 
      .ZN(n_0_2_61));
   INV_X1 i_0_2_148 (.A(n_0_2_61), .ZN(b[22]));
   OAI22_X1 i_0_2_149 (.A1(n_0_2_39), .A2(n_0_33), .B1(in_b[63]), .B2(in_b[23]), 
      .ZN(n_0_2_62));
   INV_X1 i_0_2_150 (.A(n_0_2_62), .ZN(b[23]));
   AOI22_X1 i_0_2_151 (.A1(n_0_2_39), .A2(in_b[24]), .B1(n_0_34), .B2(in_b[63]), 
      .ZN(n_0_2_63));
   INV_X1 i_0_2_152 (.A(n_0_2_63), .ZN(b[24]));
   AOI22_X1 i_0_2_153 (.A1(n_0_2_39), .A2(in_b[26]), .B1(n_0_36), .B2(in_b[63]), 
      .ZN(n_0_2_64));
   INV_X1 i_0_2_154 (.A(n_0_2_64), .ZN(b[26]));
   AOI22_X1 i_0_2_155 (.A1(n_0_2_39), .A2(in_b[25]), .B1(n_0_35), .B2(in_b[63]), 
      .ZN(n_0_2_65));
   INV_X1 i_0_2_156 (.A(n_0_2_65), .ZN(b[25]));
   OAI22_X1 i_0_2_157 (.A1(n_0_2_39), .A2(n_0_38), .B1(in_b[63]), .B2(in_b[28]), 
      .ZN(n_0_2_66));
   INV_X1 i_0_2_158 (.A(n_0_2_66), .ZN(b[28]));
   OAI22_X1 i_0_2_159 (.A1(n_0_2_39), .A2(n_0_37), .B1(in_b[63]), .B2(in_b[27]), 
      .ZN(n_0_2_67));
   INV_X1 i_0_2_160 (.A(n_0_2_67), .ZN(b[27]));
   AOI22_X1 i_0_2_161 (.A1(n_0_2_39), .A2(in_b[29]), .B1(n_0_39), .B2(in_b[63]), 
      .ZN(n_0_2_68));
   INV_X1 i_0_2_162 (.A(n_0_2_68), .ZN(b[29]));
   AOI22_X1 i_0_2_163 (.A1(n_0_2_39), .A2(in_b[30]), .B1(n_0_40), .B2(in_b[63]), 
      .ZN(n_0_2_69));
   INV_X1 i_0_2_164 (.A(n_0_2_69), .ZN(b[30]));
   OAI22_X1 i_0_2_165 (.A1(n_0_2_39), .A2(n_0_42), .B1(in_b[63]), .B2(in_b[32]), 
      .ZN(n_0_2_70));
   INV_X1 i_0_2_166 (.A(n_0_2_70), .ZN(b[32]));
   AOI22_X1 i_0_2_167 (.A1(n_0_2_39), .A2(in_b[31]), .B1(n_0_41), .B2(in_b[63]), 
      .ZN(n_0_2_71));
   INV_X1 i_0_2_168 (.A(n_0_2_71), .ZN(b[31]));
   AOI22_X1 i_0_2_169 (.A1(n_0_2_39), .A2(in_b[34]), .B1(n_0_44), .B2(in_b[63]), 
      .ZN(n_0_2_72));
   INV_X1 i_0_2_170 (.A(n_0_2_72), .ZN(b[34]));
   OAI22_X1 i_0_2_171 (.A1(n_0_2_39), .A2(n_0_43), .B1(in_b[63]), .B2(in_b[33]), 
      .ZN(n_0_2_73));
   INV_X1 i_0_2_172 (.A(n_0_2_73), .ZN(b[33]));
   AOI22_X1 i_0_2_173 (.A1(n_0_2_39), .A2(in_b[35]), .B1(n_0_45), .B2(in_b[63]), 
      .ZN(n_0_2_74));
   INV_X1 i_0_2_174 (.A(n_0_2_74), .ZN(b[35]));
   AOI22_X1 i_0_2_175 (.A1(n_0_2_39), .A2(in_b[36]), .B1(n_0_46), .B2(in_b[63]), 
      .ZN(n_0_2_75));
   INV_X1 i_0_2_176 (.A(n_0_2_75), .ZN(b[36]));
   AOI22_X1 i_0_2_177 (.A1(n_0_2_39), .A2(in_b[38]), .B1(n_0_48), .B2(in_b[63]), 
      .ZN(n_0_2_76));
   INV_X1 i_0_2_178 (.A(n_0_2_76), .ZN(b[38]));
   OAI22_X1 i_0_2_179 (.A1(n_0_2_39), .A2(n_0_47), .B1(in_b[63]), .B2(in_b[37]), 
      .ZN(n_0_2_77));
   INV_X1 i_0_2_180 (.A(n_0_2_77), .ZN(b[37]));
   AOI22_X1 i_0_2_181 (.A1(n_0_2_39), .A2(in_b[39]), .B1(n_0_49), .B2(in_b[63]), 
      .ZN(n_0_2_78));
   INV_X1 i_0_2_182 (.A(n_0_2_78), .ZN(b[39]));
   AOI22_X1 i_0_2_183 (.A1(n_0_2_39), .A2(in_b[40]), .B1(n_0_50), .B2(in_b[63]), 
      .ZN(n_0_2_79));
   INV_X1 i_0_2_184 (.A(n_0_2_79), .ZN(b[40]));
   AOI22_X1 i_0_2_185 (.A1(n_0_2_39), .A2(in_b[42]), .B1(n_0_52), .B2(in_b[63]), 
      .ZN(n_0_2_80));
   INV_X1 i_0_2_186 (.A(n_0_2_80), .ZN(b[42]));
   AOI22_X1 i_0_2_187 (.A1(n_0_2_39), .A2(in_b[41]), .B1(n_0_51), .B2(in_b[63]), 
      .ZN(n_0_2_81));
   INV_X1 i_0_2_188 (.A(n_0_2_81), .ZN(b[41]));
   AOI22_X1 i_0_2_189 (.A1(n_0_2_39), .A2(in_b[44]), .B1(n_0_54), .B2(in_b[63]), 
      .ZN(n_0_2_82));
   INV_X1 i_0_2_190 (.A(n_0_2_82), .ZN(b[44]));
   OAI22_X1 i_0_2_191 (.A1(n_0_2_39), .A2(n_0_53), .B1(in_b[63]), .B2(in_b[43]), 
      .ZN(n_0_2_83));
   INV_X1 i_0_2_192 (.A(n_0_2_83), .ZN(b[43]));
   AOI22_X1 i_0_2_193 (.A1(n_0_2_39), .A2(in_b[45]), .B1(n_0_55), .B2(in_b[63]), 
      .ZN(n_0_2_84));
   INV_X1 i_0_2_194 (.A(n_0_2_84), .ZN(b[45]));
   AOI22_X1 i_0_2_195 (.A1(n_0_2_39), .A2(in_b[46]), .B1(n_0_56), .B2(in_b[63]), 
      .ZN(n_0_2_85));
   INV_X1 i_0_2_196 (.A(n_0_2_85), .ZN(b[46]));
   AOI22_X1 i_0_2_197 (.A1(n_0_2_39), .A2(in_b[47]), .B1(n_0_57), .B2(in_b[63]), 
      .ZN(n_0_2_86));
   INV_X1 i_0_2_198 (.A(n_0_2_86), .ZN(b[47]));
   AOI22_X1 i_0_2_199 (.A1(n_0_2_39), .A2(in_b[48]), .B1(n_0_58), .B2(in_b[63]), 
      .ZN(n_0_2_87));
   INV_X1 i_0_2_200 (.A(n_0_2_87), .ZN(b[48]));
   AOI22_X1 i_0_2_201 (.A1(n_0_2_39), .A2(in_b[49]), .B1(n_0_59), .B2(in_b[63]), 
      .ZN(n_0_2_88));
   INV_X1 i_0_2_202 (.A(n_0_2_88), .ZN(b[49]));
   AOI22_X1 i_0_2_203 (.A1(n_0_2_39), .A2(in_b[50]), .B1(n_0_60), .B2(in_b[63]), 
      .ZN(n_0_2_89));
   INV_X1 i_0_2_204 (.A(n_0_2_89), .ZN(b[50]));
   OAI22_X1 i_0_2_205 (.A1(n_0_2_39), .A2(n_0_61), .B1(in_b[51]), .B2(in_b[63]), 
      .ZN(n_0_2_90));
   INV_X1 i_0_2_206 (.A(n_0_2_90), .ZN(b[51]));
   AOI22_X1 i_0_2_207 (.A1(n_0_2_39), .A2(in_b[52]), .B1(n_0_62), .B2(in_b[63]), 
      .ZN(n_0_2_91));
   INV_X1 i_0_2_208 (.A(n_0_2_91), .ZN(b[52]));
   OAI22_X1 i_0_2_209 (.A1(n_0_2_39), .A2(n_0_63), .B1(in_b[53]), .B2(in_b[63]), 
      .ZN(n_0_2_92));
   INV_X1 i_0_2_210 (.A(n_0_2_92), .ZN(b[53]));
   AOI22_X1 i_0_2_211 (.A1(n_0_2_39), .A2(in_b[54]), .B1(n_0_64), .B2(in_b[63]), 
      .ZN(n_0_2_93));
   INV_X1 i_0_2_212 (.A(n_0_2_93), .ZN(b[54]));
   AOI22_X1 i_0_2_213 (.A1(n_0_2_39), .A2(in_b[55]), .B1(n_0_65), .B2(in_b[63]), 
      .ZN(n_0_2_94));
   INV_X1 i_0_2_214 (.A(n_0_2_94), .ZN(b[55]));
   AOI22_X1 i_0_2_215 (.A1(n_0_2_39), .A2(in_b[56]), .B1(n_0_66), .B2(in_b[63]), 
      .ZN(n_0_2_95));
   INV_X1 i_0_2_216 (.A(n_0_2_95), .ZN(b[56]));
   AOI22_X1 i_0_2_217 (.A1(n_0_2_39), .A2(in_b[57]), .B1(n_0_67), .B2(in_b[63]), 
      .ZN(n_0_2_96));
   INV_X1 i_0_2_218 (.A(n_0_2_96), .ZN(b[57]));
   OAI22_X1 i_0_2_219 (.A1(n_0_2_39), .A2(n_0_68), .B1(in_b[63]), .B2(in_b[58]), 
      .ZN(n_0_2_97));
   INV_X1 i_0_2_220 (.A(n_0_2_97), .ZN(b[58]));
   AOI22_X1 i_0_2_221 (.A1(n_0_2_39), .A2(in_b[60]), .B1(n_0_70), .B2(in_b[63]), 
      .ZN(n_0_2_98));
   INV_X1 i_0_2_222 (.A(n_0_2_98), .ZN(b[60]));
   AOI22_X1 i_0_2_223 (.A1(n_0_2_39), .A2(in_b[59]), .B1(n_0_69), .B2(in_b[63]), 
      .ZN(n_0_2_99));
   INV_X1 i_0_2_224 (.A(n_0_2_99), .ZN(b[59]));
   OAI22_X1 i_0_2_225 (.A1(n_0_2_39), .A2(n_0_72), .B1(in_b[63]), .B2(in_b[62]), 
      .ZN(n_0_2_100));
   INV_X1 i_0_2_226 (.A(n_0_2_100), .ZN(b[62]));
   OAI22_X1 i_0_2_227 (.A1(n_0_2_39), .A2(n_0_71), .B1(in_b[61]), .B2(in_b[63]), 
      .ZN(n_0_2_101));
   INV_X1 i_0_2_228 (.A(n_0_2_101), .ZN(b[61]));
   NOR2_X1 i_0_2_229 (.A1(n_0_2_97), .A2(z[58]), .ZN(n_0_2_102));
   NOR2_X1 i_0_2_230 (.A1(n_0_2_83), .A2(z[43]), .ZN(n_0_2_103));
   NOR2_X1 i_0_2_231 (.A1(n_0_2_77), .A2(z[37]), .ZN(n_0_2_104));
   NOR2_X1 i_0_2_232 (.A1(n_0_2_73), .A2(z[33]), .ZN(n_0_2_105));
   INV_X1 i_0_2_233 (.A(in_b[0]), .ZN(n_0_2_106));
   OAI22_X1 i_0_2_234 (.A1(n_0_2_40), .A2(z[1]), .B1(n_0_2_106), .B2(z[0]), 
      .ZN(n_0_2_107));
   INV_X1 i_0_2_235 (.A(n_0_2_107), .ZN(n_0_2_108));
   AOI221_X1 i_0_2_236 (.A(n_0_2_108), .B1(z[2]), .B2(n_0_2_42), .C1(z[1]), 
      .C2(n_0_2_40), .ZN(n_0_2_109));
   OAI22_X1 i_0_2_237 (.A1(n_0_2_41), .A2(z[3]), .B1(n_0_2_42), .B2(z[2]), 
      .ZN(n_0_2_110));
   INV_X1 i_0_2_238 (.A(z[3]), .ZN(n_0_2_111));
   OAI22_X1 i_0_2_239 (.A1(n_0_2_109), .A2(n_0_2_110), .B1(n_0_2_111), .B2(b[3]), 
      .ZN(n_0_2_112));
   OAI21_X1 i_0_2_240 (.A(n_0_2_112), .B1(z[4]), .B2(n_0_2_43), .ZN(n_0_2_113));
   NAND2_X1 i_0_2_241 (.A1(n_0_2_45), .A2(z[5]), .ZN(n_0_2_114));
   INV_X1 i_0_2_242 (.A(z[4]), .ZN(n_0_2_115));
   OAI211_X1 i_0_2_243 (.A(n_0_2_113), .B(n_0_2_114), .C1(n_0_2_115), .C2(b[4]), 
      .ZN(n_0_2_116));
   OAI221_X1 i_0_2_244 (.A(n_0_2_116), .B1(z[6]), .B2(n_0_2_44), .C1(z[5]), 
      .C2(n_0_2_45), .ZN(n_0_2_117));
   NAND2_X1 i_0_2_245 (.A1(n_0_2_47), .A2(z[7]), .ZN(n_0_2_118));
   INV_X1 i_0_2_246 (.A(z[6]), .ZN(n_0_2_119));
   OAI211_X1 i_0_2_247 (.A(n_0_2_117), .B(n_0_2_118), .C1(n_0_2_119), .C2(b[6]), 
      .ZN(n_0_2_120));
   OAI221_X1 i_0_2_248 (.A(n_0_2_120), .B1(z[8]), .B2(n_0_2_46), .C1(z[7]), 
      .C2(n_0_2_47), .ZN(n_0_2_121));
   INV_X1 i_0_2_249 (.A(z[9]), .ZN(n_0_2_122));
   INV_X1 i_0_2_250 (.A(z[8]), .ZN(n_0_2_123));
   OAI221_X1 i_0_2_251 (.A(n_0_2_121), .B1(n_0_2_122), .B2(b[9]), .C1(n_0_2_123), 
      .C2(b[8]), .ZN(n_0_2_124));
   OAI221_X1 i_0_2_252 (.A(n_0_2_124), .B1(z[10]), .B2(n_0_2_48), .C1(z[9]), 
      .C2(n_0_2_49), .ZN(n_0_2_125));
   INV_X1 i_0_2_253 (.A(z[10]), .ZN(n_0_2_126));
   INV_X1 i_0_2_254 (.A(z[11]), .ZN(n_0_2_127));
   OAI221_X1 i_0_2_255 (.A(n_0_2_125), .B1(n_0_2_126), .B2(b[10]), .C1(n_0_2_127), 
      .C2(b[11]), .ZN(n_0_2_128));
   OAI221_X1 i_0_2_256 (.A(n_0_2_128), .B1(z[11]), .B2(n_0_2_50), .C1(z[12]), 
      .C2(n_0_2_51), .ZN(n_0_2_129));
   NAND2_X1 i_0_2_257 (.A1(n_0_2_52), .A2(z[13]), .ZN(n_0_2_130));
   INV_X1 i_0_2_258 (.A(z[12]), .ZN(n_0_2_131));
   OAI211_X1 i_0_2_259 (.A(n_0_2_129), .B(n_0_2_130), .C1(n_0_2_131), .C2(b[12]), 
      .ZN(n_0_2_132));
   OAI221_X1 i_0_2_260 (.A(n_0_2_132), .B1(z[13]), .B2(n_0_2_52), .C1(z[14]), 
      .C2(n_0_2_53), .ZN(n_0_2_133));
   INV_X1 i_0_2_261 (.A(z[15]), .ZN(n_0_2_134));
   INV_X1 i_0_2_262 (.A(z[14]), .ZN(n_0_2_135));
   OAI221_X1 i_0_2_263 (.A(n_0_2_133), .B1(n_0_2_134), .B2(b[15]), .C1(n_0_2_135), 
      .C2(b[14]), .ZN(n_0_2_136));
   OAI221_X1 i_0_2_264 (.A(n_0_2_136), .B1(z[16]), .B2(n_0_2_54), .C1(z[15]), 
      .C2(n_0_2_55), .ZN(n_0_2_137));
   NAND2_X1 i_0_2_265 (.A1(n_0_2_56), .A2(z[17]), .ZN(n_0_2_138));
   INV_X1 i_0_2_266 (.A(z[16]), .ZN(n_0_2_139));
   OAI211_X1 i_0_2_267 (.A(n_0_2_137), .B(n_0_2_138), .C1(n_0_2_139), .C2(b[16]), 
      .ZN(n_0_2_140));
   OAI221_X1 i_0_2_268 (.A(n_0_2_140), .B1(z[17]), .B2(n_0_2_56), .C1(z[18]), 
      .C2(n_0_2_57), .ZN(n_0_2_141));
   INV_X1 i_0_2_269 (.A(z[19]), .ZN(n_0_2_142));
   INV_X1 i_0_2_270 (.A(z[18]), .ZN(n_0_2_143));
   OAI221_X1 i_0_2_271 (.A(n_0_2_141), .B1(n_0_2_142), .B2(b[19]), .C1(n_0_2_143), 
      .C2(b[18]), .ZN(n_0_2_144));
   OAI221_X1 i_0_2_272 (.A(n_0_2_144), .B1(z[20]), .B2(n_0_2_58), .C1(z[19]), 
      .C2(n_0_2_59), .ZN(n_0_2_145));
   INV_X1 i_0_2_273 (.A(z[20]), .ZN(n_0_2_146));
   INV_X1 i_0_2_274 (.A(z[21]), .ZN(n_0_2_147));
   OAI221_X1 i_0_2_275 (.A(n_0_2_145), .B1(n_0_2_146), .B2(b[20]), .C1(n_0_2_147), 
      .C2(b[21]), .ZN(n_0_2_148));
   OAI221_X1 i_0_2_276 (.A(n_0_2_148), .B1(z[21]), .B2(n_0_2_60), .C1(z[22]), 
      .C2(n_0_2_61), .ZN(n_0_2_149));
   NAND2_X1 i_0_2_277 (.A1(n_0_2_62), .A2(z[23]), .ZN(n_0_2_150));
   INV_X1 i_0_2_278 (.A(z[22]), .ZN(n_0_2_151));
   OAI211_X1 i_0_2_279 (.A(n_0_2_149), .B(n_0_2_150), .C1(n_0_2_151), .C2(b[22]), 
      .ZN(n_0_2_152));
   OAI221_X1 i_0_2_280 (.A(n_0_2_152), .B1(z[23]), .B2(n_0_2_62), .C1(z[24]), 
      .C2(n_0_2_63), .ZN(n_0_2_153));
   INV_X1 i_0_2_281 (.A(z[25]), .ZN(n_0_2_154));
   INV_X1 i_0_2_282 (.A(z[24]), .ZN(n_0_2_155));
   OAI221_X1 i_0_2_283 (.A(n_0_2_153), .B1(n_0_2_154), .B2(b[25]), .C1(n_0_2_155), 
      .C2(b[24]), .ZN(n_0_2_156));
   OAI221_X1 i_0_2_284 (.A(n_0_2_156), .B1(z[26]), .B2(n_0_2_64), .C1(z[25]), 
      .C2(n_0_2_65), .ZN(n_0_2_157));
   NAND2_X1 i_0_2_285 (.A1(n_0_2_67), .A2(z[27]), .ZN(n_0_2_158));
   INV_X1 i_0_2_286 (.A(z[26]), .ZN(n_0_2_159));
   OAI211_X1 i_0_2_287 (.A(n_0_2_157), .B(n_0_2_158), .C1(n_0_2_159), .C2(b[26]), 
      .ZN(n_0_2_160));
   OAI221_X1 i_0_2_288 (.A(n_0_2_160), .B1(z[28]), .B2(n_0_2_66), .C1(z[27]), 
      .C2(n_0_2_67), .ZN(n_0_2_161));
   NAND2_X1 i_0_2_289 (.A1(n_0_2_66), .A2(z[28]), .ZN(n_0_2_162));
   INV_X1 i_0_2_290 (.A(z[29]), .ZN(n_0_2_163));
   OAI211_X1 i_0_2_291 (.A(n_0_2_161), .B(n_0_2_162), .C1(n_0_2_163), .C2(b[29]), 
      .ZN(n_0_2_164));
   OAI221_X1 i_0_2_292 (.A(n_0_2_164), .B1(z[29]), .B2(n_0_2_68), .C1(z[30]), 
      .C2(n_0_2_69), .ZN(n_0_2_165));
   INV_X1 i_0_2_293 (.A(z[31]), .ZN(n_0_2_166));
   INV_X1 i_0_2_294 (.A(z[30]), .ZN(n_0_2_167));
   OAI221_X1 i_0_2_295 (.A(n_0_2_165), .B1(n_0_2_166), .B2(b[31]), .C1(n_0_2_167), 
      .C2(b[30]), .ZN(n_0_2_168));
   OAI221_X1 i_0_2_296 (.A(n_0_2_168), .B1(z[32]), .B2(n_0_2_70), .C1(z[31]), 
      .C2(n_0_2_71), .ZN(n_0_2_169));
   INV_X1 i_0_2_297 (.A(n_0_2_169), .ZN(n_0_2_170));
   AOI221_X1 i_0_2_298 (.A(n_0_2_170), .B1(z[32]), .B2(n_0_2_70), .C1(z[33]), 
      .C2(n_0_2_73), .ZN(n_0_2_171));
   INV_X1 i_0_2_299 (.A(z[34]), .ZN(n_0_2_172));
   AOI211_X1 i_0_2_300 (.A(n_0_2_105), .B(n_0_2_171), .C1(n_0_2_172), .C2(b[34]), 
      .ZN(n_0_2_173));
   AOI221_X1 i_0_2_301 (.A(n_0_2_173), .B1(z[35]), .B2(n_0_2_74), .C1(z[34]), 
      .C2(n_0_2_72), .ZN(n_0_2_174));
   INV_X1 i_0_2_302 (.A(z[35]), .ZN(n_0_2_175));
   INV_X1 i_0_2_303 (.A(z[36]), .ZN(n_0_2_176));
   AOI221_X1 i_0_2_304 (.A(n_0_2_174), .B1(n_0_2_175), .B2(b[35]), .C1(n_0_2_176), 
      .C2(b[36]), .ZN(n_0_2_177));
   AOI221_X1 i_0_2_305 (.A(n_0_2_177), .B1(z[37]), .B2(n_0_2_77), .C1(z[36]), 
      .C2(n_0_2_75), .ZN(n_0_2_178));
   INV_X1 i_0_2_306 (.A(z[38]), .ZN(n_0_2_179));
   AOI211_X1 i_0_2_307 (.A(n_0_2_104), .B(n_0_2_178), .C1(n_0_2_179), .C2(b[38]), 
      .ZN(n_0_2_180));
   AOI221_X1 i_0_2_308 (.A(n_0_2_180), .B1(z[39]), .B2(n_0_2_78), .C1(z[38]), 
      .C2(n_0_2_76), .ZN(n_0_2_181));
   INV_X1 i_0_2_309 (.A(z[39]), .ZN(n_0_2_182));
   INV_X1 i_0_2_310 (.A(z[40]), .ZN(n_0_2_183));
   AOI221_X1 i_0_2_311 (.A(n_0_2_181), .B1(n_0_2_182), .B2(b[39]), .C1(n_0_2_183), 
      .C2(b[40]), .ZN(n_0_2_184));
   AOI221_X1 i_0_2_312 (.A(n_0_2_184), .B1(z[41]), .B2(n_0_2_81), .C1(z[40]), 
      .C2(n_0_2_79), .ZN(n_0_2_185));
   INV_X1 i_0_2_313 (.A(z[42]), .ZN(n_0_2_186));
   INV_X1 i_0_2_314 (.A(z[41]), .ZN(n_0_2_187));
   AOI221_X1 i_0_2_315 (.A(n_0_2_185), .B1(n_0_2_186), .B2(b[42]), .C1(n_0_2_187), 
      .C2(b[41]), .ZN(n_0_2_188));
   AOI221_X1 i_0_2_316 (.A(n_0_2_188), .B1(z[43]), .B2(n_0_2_83), .C1(z[42]), 
      .C2(n_0_2_80), .ZN(n_0_2_189));
   INV_X1 i_0_2_317 (.A(z[44]), .ZN(n_0_2_190));
   AOI211_X1 i_0_2_318 (.A(n_0_2_103), .B(n_0_2_189), .C1(n_0_2_190), .C2(b[44]), 
      .ZN(n_0_2_191));
   AOI221_X1 i_0_2_319 (.A(n_0_2_191), .B1(z[44]), .B2(n_0_2_82), .C1(z[45]), 
      .C2(n_0_2_84), .ZN(n_0_2_192));
   INV_X1 i_0_2_320 (.A(z[45]), .ZN(n_0_2_193));
   INV_X1 i_0_2_321 (.A(z[46]), .ZN(n_0_2_194));
   AOI221_X1 i_0_2_322 (.A(n_0_2_192), .B1(n_0_2_193), .B2(b[45]), .C1(n_0_2_194), 
      .C2(b[46]), .ZN(n_0_2_195));
   AOI221_X1 i_0_2_323 (.A(n_0_2_195), .B1(z[47]), .B2(n_0_2_86), .C1(z[46]), 
      .C2(n_0_2_85), .ZN(n_0_2_196));
   INV_X1 i_0_2_324 (.A(z[47]), .ZN(n_0_2_197));
   INV_X1 i_0_2_325 (.A(z[48]), .ZN(n_0_2_198));
   AOI221_X1 i_0_2_326 (.A(n_0_2_196), .B1(n_0_2_197), .B2(b[47]), .C1(n_0_2_198), 
      .C2(b[48]), .ZN(n_0_2_199));
   AOI221_X1 i_0_2_327 (.A(n_0_2_199), .B1(z[49]), .B2(n_0_2_88), .C1(z[48]), 
      .C2(n_0_2_87), .ZN(n_0_2_200));
   INV_X1 i_0_2_328 (.A(z[49]), .ZN(n_0_2_201));
   INV_X1 i_0_2_329 (.A(z[50]), .ZN(n_0_2_202));
   AOI221_X1 i_0_2_330 (.A(n_0_2_200), .B1(n_0_2_201), .B2(b[49]), .C1(n_0_2_202), 
      .C2(b[50]), .ZN(n_0_2_203));
   AOI221_X1 i_0_2_331 (.A(n_0_2_203), .B1(z[51]), .B2(n_0_2_90), .C1(z[50]), 
      .C2(n_0_2_89), .ZN(n_0_2_204));
   OAI22_X1 i_0_2_332 (.A1(n_0_2_90), .A2(z[51]), .B1(n_0_2_91), .B2(z[52]), 
      .ZN(n_0_2_205));
   INV_X1 i_0_2_333 (.A(z[52]), .ZN(n_0_2_206));
   OAI22_X1 i_0_2_334 (.A1(n_0_2_204), .A2(n_0_2_205), .B1(n_0_2_206), .B2(b[52]), 
      .ZN(n_0_2_207));
   OAI21_X1 i_0_2_335 (.A(n_0_2_207), .B1(z[53]), .B2(n_0_2_92), .ZN(n_0_2_208));
   NAND2_X1 i_0_2_336 (.A1(n_0_2_92), .A2(z[53]), .ZN(n_0_2_209));
   INV_X1 i_0_2_337 (.A(z[54]), .ZN(n_0_2_210));
   OAI211_X1 i_0_2_338 (.A(n_0_2_208), .B(n_0_2_209), .C1(n_0_2_210), .C2(b[54]), 
      .ZN(n_0_2_211));
   OAI221_X1 i_0_2_339 (.A(n_0_2_211), .B1(z[54]), .B2(n_0_2_93), .C1(z[55]), 
      .C2(n_0_2_94), .ZN(n_0_2_212));
   AOI22_X1 i_0_2_340 (.A1(n_0_2_94), .A2(z[55]), .B1(n_0_2_95), .B2(z[56]), 
      .ZN(n_0_2_213));
   INV_X1 i_0_2_341 (.A(z[56]), .ZN(n_0_2_214));
   AOI22_X1 i_0_2_342 (.A1(n_0_2_212), .A2(n_0_2_213), .B1(n_0_2_214), .B2(b[56]), 
      .ZN(n_0_2_215));
   AOI21_X1 i_0_2_343 (.A(n_0_2_215), .B1(z[57]), .B2(n_0_2_96), .ZN(n_0_2_216));
   INV_X1 i_0_2_344 (.A(z[57]), .ZN(n_0_2_217));
   AOI211_X1 i_0_2_345 (.A(n_0_2_102), .B(n_0_2_216), .C1(n_0_2_217), .C2(b[57]), 
      .ZN(n_0_2_218));
   AOI221_X1 i_0_2_346 (.A(n_0_2_218), .B1(z[58]), .B2(n_0_2_97), .C1(z[59]), 
      .C2(n_0_2_99), .ZN(n_0_2_219));
   INV_X1 i_0_2_347 (.A(z[60]), .ZN(n_0_2_220));
   INV_X1 i_0_2_348 (.A(z[59]), .ZN(n_0_2_221));
   AOI221_X1 i_0_2_349 (.A(n_0_2_219), .B1(n_0_2_220), .B2(b[60]), .C1(n_0_2_221), 
      .C2(b[59]), .ZN(n_0_2_222));
   AOI221_X1 i_0_2_350 (.A(n_0_2_222), .B1(z[60]), .B2(n_0_2_98), .C1(z[61]), 
      .C2(n_0_2_101), .ZN(n_0_2_223));
   INV_X1 i_0_2_351 (.A(n_0_2_223), .ZN(n_0_2_224));
   OAI221_X1 i_0_2_352 (.A(n_0_2_224), .B1(z[62]), .B2(n_0_2_100), .C1(z[61]), 
      .C2(n_0_2_101), .ZN(n_0_2_225));
   NAND2_X1 i_0_2_353 (.A1(n_0_73), .A2(in_b[63]), .ZN(n_0_2_226));
   AOI22_X1 i_0_2_354 (.A1(n_0_2_100), .A2(z[62]), .B1(n_0_2_226), .B2(z[63]), 
      .ZN(n_0_2_227));
   NAND2_X1 i_0_2_355 (.A1(n_0_2_225), .A2(n_0_2_227), .ZN(n_0_2_228));
   OAI21_X1 i_0_2_356 (.A(n_0_2_228), .B1(z[63]), .B2(n_0_2_226), .ZN(n_0_2_229));
   NOR2_X1 i_0_2_357 (.A1(n_0_2_229), .A2(n_0_2_0), .ZN(n_0_296));
   NAND2_X1 i_0_2_358 (.A1(sub[0]), .A2(state[1]), .ZN(n_0_2_230));
   INV_X1 i_0_2_359 (.A(in_a[63]), .ZN(n_0_2_231));
   OAI22_X1 i_0_2_360 (.A1(n_0_2_231), .A2(n_0_88), .B1(in_a[63]), .B2(in_a[15]), 
      .ZN(n_0_2_232));
   INV_X1 i_0_2_361 (.A(n_0_229), .ZN(n_0_2_233));
   NOR2_X1 i_0_2_362 (.A1(n_0_130), .A2(i[2]), .ZN(n_0_2_234));
   NOR2_X1 i_0_2_363 (.A1(i[0]), .A2(n_0_227), .ZN(n_0_2_235));
   NOR2_X1 i_0_2_364 (.A1(n_0_130), .A2(n_0_227), .ZN(n_0_2_236));
   AOI222_X1 i_0_2_365 (.A1(n_0_2_234), .A2(n_0_101), .B1(n_0_2_235), .B2(n_0_98), 
      .C1(n_0_2_236), .C2(n_0_97), .ZN(n_0_2_237));
   NAND2_X1 i_0_2_366 (.A1(n_0_130), .A2(n_0_227), .ZN(n_0_2_238));
   INV_X1 i_0_2_367 (.A(n_0_2_238), .ZN(n_0_2_239));
   AOI21_X1 i_0_2_368 (.A(n_0_2_231), .B1(n_0_2_239), .B2(n_0_102), .ZN(
      n_0_2_240));
   AOI221_X1 i_0_2_369 (.A(in_a[63]), .B1(n_0_2_234), .B2(in_a[28]), .C1(
      in_a[24]), .C2(n_0_2_236), .ZN(n_0_2_241));
   AOI22_X1 i_0_2_370 (.A1(n_0_2_239), .A2(in_a[29]), .B1(n_0_2_235), .B2(
      in_a[25]), .ZN(n_0_2_242));
   AOI22_X1 i_0_2_371 (.A1(n_0_2_237), .A2(n_0_2_240), .B1(n_0_2_241), .B2(
      n_0_2_242), .ZN(n_0_2_243));
   NOR2_X1 i_0_2_372 (.A1(n_0_230), .A2(i[3]), .ZN(n_0_2_244));
   INV_X1 i_0_2_373 (.A(i[3]), .ZN(n_0_2_245));
   OR2_X1 i_0_2_374 (.A1(n_0_2_245), .A2(n_0_230), .ZN(n_0_2_246));
   INV_X1 i_0_2_375 (.A(n_0_2_246), .ZN(n_0_2_247));
   AOI222_X1 i_0_2_376 (.A1(n_0_2_239), .A2(n_0_110), .B1(n_0_2_236), .B2(
      n_0_105), .C1(n_0_2_234), .C2(n_0_109), .ZN(n_0_2_248));
   AOI21_X1 i_0_2_377 (.A(n_0_2_231), .B1(n_0_2_235), .B2(n_0_106), .ZN(
      n_0_2_249));
   AOI221_X1 i_0_2_378 (.A(in_a[63]), .B1(n_0_2_234), .B2(in_a[36]), .C1(
      in_a[37]), .C2(n_0_2_239), .ZN(n_0_2_250));
   AOI22_X1 i_0_2_379 (.A1(n_0_2_235), .A2(in_a[33]), .B1(n_0_2_236), .B2(
      in_a[32]), .ZN(n_0_2_251));
   AOI22_X1 i_0_2_380 (.A1(n_0_2_248), .A2(n_0_2_249), .B1(n_0_2_250), .B2(
      n_0_2_251), .ZN(n_0_2_252));
   AOI221_X1 i_0_2_381 (.A(n_0_2_233), .B1(n_0_2_243), .B2(n_0_2_244), .C1(
      n_0_2_247), .C2(n_0_2_252), .ZN(n_0_2_253));
   NAND3_X1 i_0_2_382 (.A1(n_0_2_236), .A2(n_0_230), .A3(n_0_2_245), .ZN(
      n_0_2_254));
   AOI22_X1 i_0_2_383 (.A1(n_0_2_231), .A2(in_a[56]), .B1(n_0_129), .B2(in_a[63]), 
      .ZN(n_0_2_255));
   OAI21_X1 i_0_2_384 (.A(n_0_2_233), .B1(n_0_2_254), .B2(n_0_2_255), .ZN(
      n_0_2_256));
   OAI221_X1 i_0_2_385 (.A(n_0_2_234), .B1(in_a[4]), .B2(in_a[63]), .C1(n_0_77), 
      .C2(n_0_2_231), .ZN(n_0_2_257));
   NAND2_X1 i_0_2_386 (.A1(n_0_2_236), .A2(in_a[0]), .ZN(n_0_2_258));
   AOI221_X1 i_0_2_387 (.A(in_a[63]), .B1(n_0_2_235), .B2(in_a[1]), .C1(in_a[5]), 
      .C2(n_0_2_239), .ZN(n_0_2_259));
   AOI221_X1 i_0_2_388 (.A(n_0_2_231), .B1(n_0_2_235), .B2(n_0_74), .C1(
      n_0_2_239), .C2(n_0_78), .ZN(n_0_2_260));
   OAI211_X1 i_0_2_389 (.A(n_0_2_257), .B(n_0_2_258), .C1(n_0_2_259), .C2(
      n_0_2_260), .ZN(n_0_2_261));
   AOI21_X1 i_0_2_390 (.A(n_0_2_256), .B1(n_0_2_261), .B2(n_0_2_247), .ZN(
      n_0_2_262));
   NOR4_X1 i_0_2_391 (.A1(n_0_2_253), .A2(n_0_226), .A3(n_0_228), .A4(n_0_2_262), 
      .ZN(n_0_2_263));
   AOI22_X1 i_0_2_392 (.A1(n_0_2_239), .A2(n_0_80), .B1(n_0_2_234), .B2(n_0_79), 
      .ZN(n_0_2_264));
   AOI22_X1 i_0_2_393 (.A1(n_0_2_235), .A2(n_0_76), .B1(n_0_2_236), .B2(n_0_75), 
      .ZN(n_0_2_265));
   AOI21_X1 i_0_2_394 (.A(n_0_2_231), .B1(n_0_2_264), .B2(n_0_2_265), .ZN(
      n_0_2_266));
   AOI22_X1 i_0_2_395 (.A1(n_0_2_235), .A2(in_a[3]), .B1(n_0_2_236), .B2(in_a[2]), 
      .ZN(n_0_2_267));
   AOI22_X1 i_0_2_396 (.A1(n_0_2_239), .A2(in_a[7]), .B1(n_0_2_234), .B2(in_a[6]), 
      .ZN(n_0_2_268));
   AOI21_X1 i_0_2_397 (.A(in_a[63]), .B1(n_0_2_267), .B2(n_0_2_268), .ZN(
      n_0_2_269));
   OR3_X1 i_0_2_398 (.A1(n_0_2_266), .A2(n_0_2_269), .A3(n_0_228), .ZN(n_0_2_270));
   AOI21_X1 i_0_2_399 (.A(n_0_229), .B1(n_0_2_270), .B2(n_0_2_247), .ZN(
      n_0_2_271));
   AOI22_X1 i_0_2_400 (.A1(n_0_2_235), .A2(in_a[19]), .B1(n_0_2_234), .B2(
      in_a[22]), .ZN(n_0_2_272));
   AOI22_X1 i_0_2_401 (.A1(n_0_2_239), .A2(in_a[23]), .B1(n_0_2_236), .B2(
      in_a[18]), .ZN(n_0_2_273));
   NAND3_X1 i_0_2_402 (.A1(n_0_2_272), .A2(n_0_2_273), .A3(n_0_2_231), .ZN(
      n_0_2_274));
   AOI22_X1 i_0_2_403 (.A1(n_0_2_235), .A2(n_0_92), .B1(n_0_2_234), .B2(n_0_95), 
      .ZN(n_0_2_275));
   AOI22_X1 i_0_2_404 (.A1(n_0_2_239), .A2(n_0_96), .B1(n_0_2_236), .B2(n_0_91), 
      .ZN(n_0_2_276));
   NAND3_X1 i_0_2_405 (.A1(n_0_2_275), .A2(n_0_2_276), .A3(in_a[63]), .ZN(
      n_0_2_277));
   NAND3_X1 i_0_2_406 (.A1(n_0_2_274), .A2(n_0_2_277), .A3(n_0_2_233), .ZN(
      n_0_2_278));
   AOI21_X1 i_0_2_407 (.A(n_0_2_271), .B1(n_0_228), .B2(n_0_2_278), .ZN(
      n_0_2_279));
   AOI22_X1 i_0_2_408 (.A1(n_0_2_239), .A2(in_a[39]), .B1(n_0_2_236), .B2(
      in_a[34]), .ZN(n_0_2_280));
   AOI22_X1 i_0_2_409 (.A1(n_0_2_234), .A2(in_a[38]), .B1(n_0_2_235), .B2(
      in_a[35]), .ZN(n_0_2_281));
   AND2_X1 i_0_2_410 (.A1(n_0_2_280), .A2(n_0_2_281), .ZN(n_0_2_282));
   OAI21_X1 i_0_2_411 (.A(n_0_229), .B1(n_0_2_282), .B2(in_a[63]), .ZN(n_0_2_283));
   AOI22_X1 i_0_2_412 (.A1(n_0_2_234), .A2(n_0_111), .B1(n_0_2_235), .B2(n_0_108), 
      .ZN(n_0_2_284));
   AOI22_X1 i_0_2_413 (.A1(n_0_2_239), .A2(n_0_112), .B1(n_0_2_236), .B2(n_0_107), 
      .ZN(n_0_2_285));
   AOI21_X1 i_0_2_414 (.A(n_0_2_231), .B1(n_0_2_284), .B2(n_0_2_285), .ZN(
      n_0_2_286));
   OAI21_X1 i_0_2_415 (.A(n_0_2_247), .B1(n_0_2_283), .B2(n_0_2_286), .ZN(
      n_0_2_287));
   AOI22_X1 i_0_2_416 (.A1(n_0_2_239), .A2(n_0_104), .B1(n_0_2_235), .B2(n_0_100), 
      .ZN(n_0_2_288));
   AOI22_X1 i_0_2_417 (.A1(n_0_2_234), .A2(n_0_103), .B1(n_0_2_236), .B2(n_0_99), 
      .ZN(n_0_2_289));
   AOI21_X1 i_0_2_418 (.A(n_0_2_231), .B1(n_0_2_288), .B2(n_0_2_289), .ZN(
      n_0_2_290));
   AOI22_X1 i_0_2_419 (.A1(n_0_2_239), .A2(in_a[31]), .B1(n_0_2_235), .B2(
      in_a[27]), .ZN(n_0_2_291));
   AOI22_X1 i_0_2_420 (.A1(n_0_2_234), .A2(in_a[30]), .B1(n_0_2_236), .B2(
      in_a[26]), .ZN(n_0_2_292));
   AOI21_X1 i_0_2_421 (.A(in_a[63]), .B1(n_0_2_291), .B2(n_0_2_292), .ZN(
      n_0_2_293));
   OAI21_X1 i_0_2_422 (.A(n_0_2_244), .B1(n_0_2_290), .B2(n_0_2_293), .ZN(
      n_0_2_294));
   AOI21_X1 i_0_2_423 (.A(i[1]), .B1(n_0_2_287), .B2(n_0_2_294), .ZN(n_0_2_295));
   AOI221_X1 i_0_2_424 (.A(in_a[63]), .B1(n_0_2_235), .B2(in_a[41]), .C1(
      n_0_2_239), .C2(in_a[45]), .ZN(n_0_2_296));
   AOI22_X1 i_0_2_425 (.A1(n_0_2_234), .A2(in_a[44]), .B1(n_0_2_236), .B2(
      in_a[40]), .ZN(n_0_2_297));
   AOI222_X1 i_0_2_426 (.A1(n_0_2_239), .A2(n_0_118), .B1(n_0_2_236), .B2(
      n_0_113), .C1(n_0_2_235), .C2(n_0_114), .ZN(n_0_2_298));
   AOI21_X1 i_0_2_427 (.A(n_0_2_231), .B1(n_0_2_234), .B2(n_0_117), .ZN(
      n_0_2_299));
   AOI221_X1 i_0_2_428 (.A(n_0_226), .B1(n_0_2_296), .B2(n_0_2_297), .C1(
      n_0_2_298), .C2(n_0_2_299), .ZN(n_0_2_300));
   AOI221_X1 i_0_2_429 (.A(in_a[63]), .B1(n_0_2_235), .B2(in_a[43]), .C1(
      in_a[42]), .C2(n_0_2_236), .ZN(n_0_2_301));
   AOI22_X1 i_0_2_430 (.A1(n_0_2_239), .A2(in_a[47]), .B1(n_0_2_234), .B2(
      in_a[46]), .ZN(n_0_2_302));
   AOI222_X1 i_0_2_431 (.A1(n_0_120), .A2(n_0_2_239), .B1(n_0_2_235), .B2(
      n_0_116), .C1(n_0_2_234), .C2(n_0_119), .ZN(n_0_2_303));
   AOI21_X1 i_0_2_432 (.A(n_0_2_231), .B1(n_0_2_236), .B2(n_0_115), .ZN(
      n_0_2_304));
   AOI221_X1 i_0_2_433 (.A(i[1]), .B1(n_0_2_301), .B2(n_0_2_302), .C1(n_0_2_303), 
      .C2(n_0_2_304), .ZN(n_0_2_305));
   OAI21_X1 i_0_2_434 (.A(n_0_2_244), .B1(n_0_2_300), .B2(n_0_2_305), .ZN(
      n_0_2_306));
   AOI22_X1 i_0_2_435 (.A1(n_0_2_236), .A2(in_a[50]), .B1(n_0_2_234), .B2(
      in_a[54]), .ZN(n_0_2_307));
   INV_X1 i_0_2_436 (.A(n_0_2_307), .ZN(n_0_2_308));
   AOI221_X1 i_0_2_437 (.A(n_0_2_308), .B1(in_a[51]), .B2(n_0_2_235), .C1(
      in_a[55]), .C2(n_0_2_239), .ZN(n_0_2_309));
   AOI22_X1 i_0_2_438 (.A1(n_0_2_239), .A2(n_0_128), .B1(n_0_2_235), .B2(n_0_124), 
      .ZN(n_0_2_310));
   INV_X1 i_0_2_439 (.A(n_0_2_310), .ZN(n_0_2_311));
   AOI221_X1 i_0_2_440 (.A(n_0_2_311), .B1(n_0_123), .B2(n_0_2_236), .C1(n_0_127), 
      .C2(n_0_2_234), .ZN(n_0_2_312));
   AOI221_X1 i_0_2_441 (.A(i[1]), .B1(n_0_2_309), .B2(n_0_2_231), .C1(in_a[63]), 
      .C2(n_0_2_312), .ZN(n_0_2_313));
   AOI22_X1 i_0_2_442 (.A1(n_0_2_235), .A2(n_0_122), .B1(n_0_2_234), .B2(n_0_125), 
      .ZN(n_0_2_314));
   AOI22_X1 i_0_2_443 (.A1(n_0_2_239), .A2(n_0_126), .B1(n_0_2_236), .B2(n_0_121), 
      .ZN(n_0_2_315));
   NAND3_X1 i_0_2_444 (.A1(n_0_2_314), .A2(n_0_2_315), .A3(in_a[63]), .ZN(
      n_0_2_316));
   AOI22_X1 i_0_2_445 (.A1(n_0_2_234), .A2(in_a[52]), .B1(n_0_2_235), .B2(
      in_a[49]), .ZN(n_0_2_317));
   AOI22_X1 i_0_2_446 (.A1(n_0_2_239), .A2(in_a[53]), .B1(n_0_2_236), .B2(
      in_a[48]), .ZN(n_0_2_318));
   NAND3_X1 i_0_2_447 (.A1(n_0_2_317), .A2(n_0_2_318), .A3(n_0_2_231), .ZN(
      n_0_2_319));
   AND2_X1 i_0_2_448 (.A1(n_0_2_316), .A2(n_0_2_319), .ZN(n_0_2_320));
   AOI21_X1 i_0_2_449 (.A(n_0_2_313), .B1(i[1]), .B2(n_0_2_320), .ZN(n_0_2_321));
   OAI21_X1 i_0_2_450 (.A(n_0_2_306), .B1(n_0_2_321), .B2(n_0_2_246), .ZN(
      n_0_2_322));
   AOI22_X1 i_0_2_451 (.A1(n_0_2_235), .A2(n_0_90), .B1(n_0_2_234), .B2(n_0_93), 
      .ZN(n_0_2_323));
   AOI22_X1 i_0_2_452 (.A1(n_0_2_239), .A2(n_0_94), .B1(n_0_2_236), .B2(n_0_89), 
      .ZN(n_0_2_324));
   AOI21_X1 i_0_2_453 (.A(n_0_2_231), .B1(n_0_2_323), .B2(n_0_2_324), .ZN(
      n_0_2_325));
   AOI22_X1 i_0_2_454 (.A1(n_0_2_239), .A2(in_a[21]), .B1(n_0_2_235), .B2(
      in_a[17]), .ZN(n_0_2_326));
   AOI22_X1 i_0_2_455 (.A1(n_0_2_234), .A2(in_a[20]), .B1(n_0_2_236), .B2(
      in_a[16]), .ZN(n_0_2_327));
   AOI21_X1 i_0_2_456 (.A(in_a[63]), .B1(n_0_2_326), .B2(n_0_2_327), .ZN(
      n_0_2_328));
   OAI211_X1 i_0_2_457 (.A(i[1]), .B(n_0_2_247), .C1(n_0_2_325), .C2(n_0_2_328), 
      .ZN(n_0_2_329));
   AOI221_X1 i_0_2_458 (.A(n_0_2_231), .B1(n_0_2_234), .B2(n_0_85), .C1(n_0_82), 
      .C2(n_0_2_235), .ZN(n_0_2_330));
   AOI22_X1 i_0_2_459 (.A1(n_0_2_239), .A2(n_0_86), .B1(n_0_2_236), .B2(n_0_81), 
      .ZN(n_0_2_331));
   AOI222_X1 i_0_2_460 (.A1(n_0_2_239), .A2(in_a[13]), .B1(n_0_2_234), .B2(
      in_a[12]), .C1(n_0_2_235), .C2(in_a[9]), .ZN(n_0_2_332));
   AOI21_X1 i_0_2_461 (.A(in_a[63]), .B1(n_0_2_236), .B2(in_a[8]), .ZN(n_0_2_333));
   AOI221_X1 i_0_2_462 (.A(n_0_226), .B1(n_0_2_330), .B2(n_0_2_331), .C1(
      n_0_2_332), .C2(n_0_2_333), .ZN(n_0_2_334));
   AOI222_X1 i_0_2_463 (.A1(n_0_2_236), .A2(in_a[10]), .B1(n_0_2_234), .B2(
      in_a[14]), .C1(n_0_2_235), .C2(in_a[11]), .ZN(n_0_2_335));
   AOI21_X1 i_0_2_464 (.A(n_0_2_231), .B1(n_0_2_235), .B2(n_0_84), .ZN(n_0_2_336));
   AOI22_X1 i_0_2_465 (.A1(n_0_2_236), .A2(n_0_83), .B1(n_0_2_234), .B2(n_0_87), 
      .ZN(n_0_2_337));
   AOI22_X1 i_0_2_466 (.A1(n_0_2_335), .A2(n_0_2_231), .B1(n_0_2_336), .B2(
      n_0_2_337), .ZN(n_0_2_338));
   INV_X1 i_0_2_467 (.A(n_0_2_338), .ZN(n_0_2_339));
   OAI21_X1 i_0_2_468 (.A(n_0_2_339), .B1(n_0_2_232), .B2(n_0_2_238), .ZN(
      n_0_2_340));
   AOI21_X1 i_0_2_469 (.A(n_0_2_334), .B1(n_0_2_340), .B2(n_0_226), .ZN(
      n_0_2_341));
   INV_X1 i_0_2_470 (.A(n_0_2_244), .ZN(n_0_2_342));
   OAI21_X1 i_0_2_471 (.A(n_0_2_329), .B1(n_0_2_341), .B2(n_0_2_342), .ZN(
      n_0_2_343));
   AOI22_X1 i_0_2_472 (.A1(n_0_2_322), .A2(n_0_229), .B1(n_0_2_343), .B2(
      n_0_2_233), .ZN(n_0_2_344));
   INV_X1 i_0_2_473 (.A(n_0_2_344), .ZN(n_0_2_345));
   AOI221_X1 i_0_2_474 (.A(n_0_2_263), .B1(n_0_2_279), .B2(n_0_2_295), .C1(
      n_0_2_345), .C2(n_0_228), .ZN(n_0_2_346));
   INV_X1 i_0_2_475 (.A(state[0]), .ZN(n_0_2_347));
   OAI221_X1 i_0_2_476 (.A(n_0_2_230), .B1(n_0_2_232), .B2(n_0_298), .C1(
      n_0_2_346), .C2(n_0_2_347), .ZN(z_next_reg[0]));
   OAI22_X1 i_0_2_477 (.A1(n_0_2_15), .A2(sub[1]), .B1(z[0]), .B2(state[1]), 
      .ZN(n_0_2_348));
   INV_X1 i_0_2_478 (.A(n_0_2_348), .ZN(z_next_reg[1]));
   OAI22_X1 i_0_2_479 (.A1(n_0_2_15), .A2(sub[2]), .B1(z[1]), .B2(state[1]), 
      .ZN(n_0_2_349));
   INV_X1 i_0_2_480 (.A(n_0_2_349), .ZN(z_next_reg[2]));
   OAI22_X1 i_0_2_481 (.A1(n_0_2_15), .A2(sub[3]), .B1(z[2]), .B2(state[1]), 
      .ZN(n_0_2_350));
   INV_X1 i_0_2_482 (.A(n_0_2_350), .ZN(z_next_reg[3]));
   OAI22_X1 i_0_2_483 (.A1(n_0_2_15), .A2(sub[4]), .B1(z[3]), .B2(state[1]), 
      .ZN(n_0_2_351));
   INV_X1 i_0_2_484 (.A(n_0_2_351), .ZN(z_next_reg[4]));
   OAI22_X1 i_0_2_485 (.A1(n_0_2_15), .A2(sub[5]), .B1(z[4]), .B2(state[1]), 
      .ZN(n_0_2_352));
   INV_X1 i_0_2_486 (.A(n_0_2_352), .ZN(z_next_reg[5]));
   OAI22_X1 i_0_2_487 (.A1(n_0_2_15), .A2(sub[6]), .B1(z[5]), .B2(state[1]), 
      .ZN(n_0_2_353));
   INV_X1 i_0_2_488 (.A(n_0_2_353), .ZN(z_next_reg[6]));
   OAI22_X1 i_0_2_489 (.A1(n_0_2_15), .A2(sub[7]), .B1(z[6]), .B2(state[1]), 
      .ZN(n_0_2_354));
   INV_X1 i_0_2_490 (.A(n_0_2_354), .ZN(z_next_reg[7]));
   OAI22_X1 i_0_2_491 (.A1(n_0_2_15), .A2(sub[8]), .B1(z[7]), .B2(state[1]), 
      .ZN(n_0_2_355));
   INV_X1 i_0_2_492 (.A(n_0_2_355), .ZN(z_next_reg[8]));
   OAI22_X1 i_0_2_493 (.A1(n_0_2_15), .A2(sub[9]), .B1(z[8]), .B2(state[1]), 
      .ZN(n_0_2_356));
   INV_X1 i_0_2_494 (.A(n_0_2_356), .ZN(z_next_reg[9]));
   OAI22_X1 i_0_2_495 (.A1(n_0_2_15), .A2(sub[10]), .B1(z[9]), .B2(state[1]), 
      .ZN(n_0_2_357));
   INV_X1 i_0_2_496 (.A(n_0_2_357), .ZN(z_next_reg[10]));
   OAI22_X1 i_0_2_497 (.A1(n_0_2_15), .A2(sub[11]), .B1(z[10]), .B2(state[1]), 
      .ZN(n_0_2_358));
   INV_X1 i_0_2_498 (.A(n_0_2_358), .ZN(z_next_reg[11]));
   OAI22_X1 i_0_2_499 (.A1(n_0_2_15), .A2(sub[12]), .B1(z[11]), .B2(state[1]), 
      .ZN(n_0_2_359));
   INV_X1 i_0_2_500 (.A(n_0_2_359), .ZN(z_next_reg[12]));
   OAI22_X1 i_0_2_501 (.A1(n_0_2_15), .A2(sub[13]), .B1(z[12]), .B2(state[1]), 
      .ZN(n_0_2_360));
   INV_X1 i_0_2_502 (.A(n_0_2_360), .ZN(z_next_reg[13]));
   OAI22_X1 i_0_2_503 (.A1(n_0_2_15), .A2(sub[14]), .B1(z[13]), .B2(state[1]), 
      .ZN(n_0_2_361));
   INV_X1 i_0_2_504 (.A(n_0_2_361), .ZN(z_next_reg[14]));
   OAI22_X1 i_0_2_505 (.A1(n_0_2_15), .A2(sub[15]), .B1(z[14]), .B2(state[1]), 
      .ZN(n_0_2_362));
   INV_X1 i_0_2_506 (.A(n_0_2_362), .ZN(z_next_reg[15]));
   OAI22_X1 i_0_2_507 (.A1(n_0_2_15), .A2(sub[16]), .B1(z[15]), .B2(state[1]), 
      .ZN(n_0_2_363));
   INV_X1 i_0_2_508 (.A(n_0_2_363), .ZN(z_next_reg[16]));
   OAI22_X1 i_0_2_509 (.A1(n_0_2_15), .A2(sub[17]), .B1(z[16]), .B2(state[1]), 
      .ZN(n_0_2_364));
   INV_X1 i_0_2_510 (.A(n_0_2_364), .ZN(z_next_reg[17]));
   OAI22_X1 i_0_2_511 (.A1(n_0_2_15), .A2(sub[18]), .B1(z[17]), .B2(state[1]), 
      .ZN(n_0_2_365));
   INV_X1 i_0_2_512 (.A(n_0_2_365), .ZN(z_next_reg[18]));
   OAI22_X1 i_0_2_513 (.A1(n_0_2_15), .A2(sub[19]), .B1(z[18]), .B2(state[1]), 
      .ZN(n_0_2_366));
   INV_X1 i_0_2_514 (.A(n_0_2_366), .ZN(z_next_reg[19]));
   OAI22_X1 i_0_2_515 (.A1(n_0_2_15), .A2(sub[20]), .B1(z[19]), .B2(state[1]), 
      .ZN(n_0_2_367));
   INV_X1 i_0_2_516 (.A(n_0_2_367), .ZN(z_next_reg[20]));
   OAI22_X1 i_0_2_517 (.A1(n_0_2_15), .A2(sub[21]), .B1(z[20]), .B2(state[1]), 
      .ZN(n_0_2_368));
   INV_X1 i_0_2_518 (.A(n_0_2_368), .ZN(z_next_reg[21]));
   OAI22_X1 i_0_2_519 (.A1(n_0_2_15), .A2(sub[22]), .B1(z[21]), .B2(state[1]), 
      .ZN(n_0_2_369));
   INV_X1 i_0_2_520 (.A(n_0_2_369), .ZN(z_next_reg[22]));
   OAI22_X1 i_0_2_521 (.A1(n_0_2_15), .A2(sub[23]), .B1(z[22]), .B2(state[1]), 
      .ZN(n_0_2_370));
   INV_X1 i_0_2_522 (.A(n_0_2_370), .ZN(z_next_reg[23]));
   OAI22_X1 i_0_2_523 (.A1(n_0_2_15), .A2(sub[24]), .B1(z[23]), .B2(state[1]), 
      .ZN(n_0_2_371));
   INV_X1 i_0_2_524 (.A(n_0_2_371), .ZN(z_next_reg[24]));
   OAI22_X1 i_0_2_525 (.A1(n_0_2_15), .A2(sub[25]), .B1(z[24]), .B2(state[1]), 
      .ZN(n_0_2_372));
   INV_X1 i_0_2_526 (.A(n_0_2_372), .ZN(z_next_reg[25]));
   OAI22_X1 i_0_2_527 (.A1(n_0_2_15), .A2(sub[26]), .B1(z[25]), .B2(state[1]), 
      .ZN(n_0_2_373));
   INV_X1 i_0_2_528 (.A(n_0_2_373), .ZN(z_next_reg[26]));
   OAI22_X1 i_0_2_529 (.A1(n_0_2_15), .A2(sub[27]), .B1(z[26]), .B2(state[1]), 
      .ZN(n_0_2_374));
   INV_X1 i_0_2_530 (.A(n_0_2_374), .ZN(z_next_reg[27]));
   OAI22_X1 i_0_2_531 (.A1(n_0_2_15), .A2(sub[28]), .B1(z[27]), .B2(state[1]), 
      .ZN(n_0_2_375));
   INV_X1 i_0_2_532 (.A(n_0_2_375), .ZN(z_next_reg[28]));
   OAI22_X1 i_0_2_533 (.A1(n_0_2_15), .A2(sub[29]), .B1(z[28]), .B2(state[1]), 
      .ZN(n_0_2_376));
   INV_X1 i_0_2_534 (.A(n_0_2_376), .ZN(z_next_reg[29]));
   OAI22_X1 i_0_2_535 (.A1(n_0_2_15), .A2(sub[30]), .B1(z[29]), .B2(state[1]), 
      .ZN(n_0_2_377));
   INV_X1 i_0_2_536 (.A(n_0_2_377), .ZN(z_next_reg[30]));
   OAI22_X1 i_0_2_537 (.A1(n_0_2_15), .A2(sub[31]), .B1(z[30]), .B2(state[1]), 
      .ZN(n_0_2_378));
   INV_X1 i_0_2_538 (.A(n_0_2_378), .ZN(z_next_reg[31]));
   OAI22_X1 i_0_2_539 (.A1(n_0_2_15), .A2(sub[32]), .B1(z[31]), .B2(state[1]), 
      .ZN(n_0_2_379));
   INV_X1 i_0_2_540 (.A(n_0_2_379), .ZN(z_next_reg[32]));
   OAI22_X1 i_0_2_541 (.A1(n_0_2_15), .A2(sub[33]), .B1(z[32]), .B2(state[1]), 
      .ZN(n_0_2_380));
   INV_X1 i_0_2_542 (.A(n_0_2_380), .ZN(z_next_reg[33]));
   OAI22_X1 i_0_2_543 (.A1(n_0_2_15), .A2(sub[34]), .B1(z[33]), .B2(state[1]), 
      .ZN(n_0_2_381));
   INV_X1 i_0_2_544 (.A(n_0_2_381), .ZN(z_next_reg[34]));
   OAI22_X1 i_0_2_545 (.A1(n_0_2_15), .A2(sub[35]), .B1(z[34]), .B2(state[1]), 
      .ZN(n_0_2_382));
   INV_X1 i_0_2_546 (.A(n_0_2_382), .ZN(z_next_reg[35]));
   OAI22_X1 i_0_2_547 (.A1(n_0_2_15), .A2(sub[36]), .B1(z[35]), .B2(state[1]), 
      .ZN(n_0_2_383));
   INV_X1 i_0_2_548 (.A(n_0_2_383), .ZN(z_next_reg[36]));
   OAI22_X1 i_0_2_549 (.A1(n_0_2_15), .A2(sub[37]), .B1(z[36]), .B2(state[1]), 
      .ZN(n_0_2_384));
   INV_X1 i_0_2_550 (.A(n_0_2_384), .ZN(z_next_reg[37]));
   OAI22_X1 i_0_2_551 (.A1(n_0_2_15), .A2(sub[38]), .B1(z[37]), .B2(state[1]), 
      .ZN(n_0_2_385));
   INV_X1 i_0_2_552 (.A(n_0_2_385), .ZN(z_next_reg[38]));
   OAI22_X1 i_0_2_553 (.A1(n_0_2_15), .A2(sub[39]), .B1(z[38]), .B2(state[1]), 
      .ZN(n_0_2_386));
   INV_X1 i_0_2_554 (.A(n_0_2_386), .ZN(z_next_reg[39]));
   OAI22_X1 i_0_2_555 (.A1(n_0_2_15), .A2(sub[40]), .B1(z[39]), .B2(state[1]), 
      .ZN(n_0_2_387));
   INV_X1 i_0_2_556 (.A(n_0_2_387), .ZN(z_next_reg[40]));
   OAI22_X1 i_0_2_557 (.A1(n_0_2_15), .A2(sub[41]), .B1(z[40]), .B2(state[1]), 
      .ZN(n_0_2_388));
   INV_X1 i_0_2_558 (.A(n_0_2_388), .ZN(z_next_reg[41]));
   OAI22_X1 i_0_2_559 (.A1(n_0_2_15), .A2(sub[42]), .B1(z[41]), .B2(state[1]), 
      .ZN(n_0_2_389));
   INV_X1 i_0_2_560 (.A(n_0_2_389), .ZN(z_next_reg[42]));
   OAI22_X1 i_0_2_561 (.A1(n_0_2_15), .A2(sub[43]), .B1(z[42]), .B2(state[1]), 
      .ZN(n_0_2_390));
   INV_X1 i_0_2_562 (.A(n_0_2_390), .ZN(z_next_reg[43]));
   OAI22_X1 i_0_2_563 (.A1(n_0_2_15), .A2(sub[44]), .B1(z[43]), .B2(state[1]), 
      .ZN(n_0_2_391));
   INV_X1 i_0_2_564 (.A(n_0_2_391), .ZN(z_next_reg[44]));
   OAI22_X1 i_0_2_565 (.A1(n_0_2_15), .A2(sub[45]), .B1(z[44]), .B2(state[1]), 
      .ZN(n_0_2_392));
   INV_X1 i_0_2_566 (.A(n_0_2_392), .ZN(z_next_reg[45]));
   OAI22_X1 i_0_2_567 (.A1(n_0_2_15), .A2(sub[46]), .B1(z[45]), .B2(state[1]), 
      .ZN(n_0_2_393));
   INV_X1 i_0_2_568 (.A(n_0_2_393), .ZN(z_next_reg[46]));
   OAI22_X1 i_0_2_569 (.A1(n_0_2_15), .A2(sub[47]), .B1(z[46]), .B2(state[1]), 
      .ZN(n_0_2_394));
   INV_X1 i_0_2_570 (.A(n_0_2_394), .ZN(z_next_reg[47]));
   OAI22_X1 i_0_2_571 (.A1(n_0_2_15), .A2(sub[48]), .B1(z[47]), .B2(state[1]), 
      .ZN(n_0_2_395));
   INV_X1 i_0_2_572 (.A(n_0_2_395), .ZN(z_next_reg[48]));
   OAI22_X1 i_0_2_573 (.A1(n_0_2_15), .A2(sub[49]), .B1(z[48]), .B2(state[1]), 
      .ZN(n_0_2_396));
   INV_X1 i_0_2_574 (.A(n_0_2_396), .ZN(z_next_reg[49]));
   OAI22_X1 i_0_2_575 (.A1(n_0_2_15), .A2(sub[50]), .B1(z[49]), .B2(state[1]), 
      .ZN(n_0_2_397));
   INV_X1 i_0_2_576 (.A(n_0_2_397), .ZN(z_next_reg[50]));
   OAI22_X1 i_0_2_577 (.A1(n_0_2_15), .A2(sub[51]), .B1(z[50]), .B2(state[1]), 
      .ZN(n_0_2_398));
   INV_X1 i_0_2_578 (.A(n_0_2_398), .ZN(z_next_reg[51]));
   OAI22_X1 i_0_2_579 (.A1(n_0_2_15), .A2(sub[52]), .B1(z[51]), .B2(state[1]), 
      .ZN(n_0_2_399));
   INV_X1 i_0_2_580 (.A(n_0_2_399), .ZN(z_next_reg[52]));
   OAI22_X1 i_0_2_581 (.A1(n_0_2_15), .A2(sub[53]), .B1(z[52]), .B2(state[1]), 
      .ZN(n_0_2_400));
   INV_X1 i_0_2_582 (.A(n_0_2_400), .ZN(z_next_reg[53]));
   OAI22_X1 i_0_2_583 (.A1(n_0_2_15), .A2(sub[54]), .B1(z[53]), .B2(state[1]), 
      .ZN(n_0_2_401));
   INV_X1 i_0_2_584 (.A(n_0_2_401), .ZN(z_next_reg[54]));
   OAI22_X1 i_0_2_585 (.A1(n_0_2_15), .A2(sub[55]), .B1(z[54]), .B2(state[1]), 
      .ZN(n_0_2_402));
   INV_X1 i_0_2_586 (.A(n_0_2_402), .ZN(z_next_reg[55]));
   OAI22_X1 i_0_2_587 (.A1(n_0_2_15), .A2(sub[56]), .B1(z[55]), .B2(state[1]), 
      .ZN(n_0_2_403));
   INV_X1 i_0_2_588 (.A(n_0_2_403), .ZN(z_next_reg[56]));
   OAI22_X1 i_0_2_589 (.A1(n_0_2_15), .A2(sub[57]), .B1(z[56]), .B2(state[1]), 
      .ZN(n_0_2_404));
   INV_X1 i_0_2_590 (.A(n_0_2_404), .ZN(z_next_reg[57]));
   OAI22_X1 i_0_2_591 (.A1(n_0_2_15), .A2(sub[58]), .B1(z[57]), .B2(state[1]), 
      .ZN(n_0_2_405));
   INV_X1 i_0_2_592 (.A(n_0_2_405), .ZN(z_next_reg[58]));
   OAI22_X1 i_0_2_593 (.A1(n_0_2_15), .A2(sub[59]), .B1(z[58]), .B2(state[1]), 
      .ZN(n_0_2_406));
   INV_X1 i_0_2_594 (.A(n_0_2_406), .ZN(z_next_reg[59]));
   OAI22_X1 i_0_2_595 (.A1(n_0_2_15), .A2(sub[60]), .B1(z[59]), .B2(state[1]), 
      .ZN(n_0_2_407));
   INV_X1 i_0_2_596 (.A(n_0_2_407), .ZN(z_next_reg[60]));
   OAI22_X1 i_0_2_597 (.A1(n_0_2_15), .A2(sub[61]), .B1(z[60]), .B2(state[1]), 
      .ZN(n_0_2_408));
   INV_X1 i_0_2_598 (.A(n_0_2_408), .ZN(z_next_reg[61]));
   OAI22_X1 i_0_2_599 (.A1(n_0_2_15), .A2(sub[62]), .B1(z[61]), .B2(state[1]), 
      .ZN(n_0_2_409));
   INV_X1 i_0_2_600 (.A(n_0_2_409), .ZN(z_next_reg[62]));
   OAI22_X1 i_0_2_601 (.A1(n_0_2_15), .A2(sub[63]), .B1(z[62]), .B2(state[1]), 
      .ZN(n_0_2_410));
   INV_X1 i_0_2_602 (.A(n_0_2_410), .ZN(z_next_reg[63]));
   NAND2_X1 i_0_2_603 (.A1(n_0_2_229), .A2(state[1]), .ZN(n_0_297));
   AOI22_X1 i_0_2_604 (.A1(n_0_132), .A2(state[1]), .B1(i[2]), .B2(state[0]), 
      .ZN(n_0_2_411));
   INV_X1 i_0_2_605 (.A(n_0_2_411), .ZN(i_next_reg[2]));
   AOI22_X1 i_0_2_606 (.A1(n_0_131), .A2(state[1]), .B1(i[1]), .B2(state[0]), 
      .ZN(n_0_2_412));
   INV_X1 i_0_2_607 (.A(n_0_2_412), .ZN(i_next_reg[1]));
   AOI22_X1 i_0_2_608 (.A1(n_0_130), .A2(state[1]), .B1(i[0]), .B2(state[0]), 
      .ZN(n_0_2_413));
   INV_X1 i_0_2_609 (.A(n_0_2_413), .ZN(i_next_reg[0]));
   AOI22_X1 i_0_2_610 (.A1(n_0_137), .A2(state[1]), .B1(i[7]), .B2(state[0]), 
      .ZN(n_0_2_414));
   INV_X1 i_0_2_611 (.A(n_0_2_414), .ZN(i_next_reg[7]));
   AOI22_X1 i_0_2_612 (.A1(n_0_136), .A2(state[1]), .B1(i[6]), .B2(state[0]), 
      .ZN(n_0_2_415));
   INV_X1 i_0_2_613 (.A(n_0_2_415), .ZN(i_next_reg[6]));
   AOI22_X1 i_0_2_614 (.A1(n_0_135), .A2(state[1]), .B1(i[5]), .B2(state[0]), 
      .ZN(n_0_2_416));
   INV_X1 i_0_2_615 (.A(n_0_2_416), .ZN(i_next_reg[5]));
   AOI22_X1 i_0_2_616 (.A1(n_0_142), .A2(state[1]), .B1(i[12]), .B2(state[0]), 
      .ZN(n_0_2_417));
   INV_X1 i_0_2_617 (.A(n_0_2_417), .ZN(i_next_reg[12]));
   AOI22_X1 i_0_2_618 (.A1(n_0_138), .A2(state[1]), .B1(i[8]), .B2(state[0]), 
      .ZN(n_0_2_418));
   INV_X1 i_0_2_619 (.A(n_0_2_418), .ZN(i_next_reg[8]));
   AOI22_X1 i_0_2_620 (.A1(i[20]), .A2(state[0]), .B1(n_0_150), .B2(state[1]), 
      .ZN(n_0_2_419));
   INV_X1 i_0_2_621 (.A(n_0_2_419), .ZN(i_next_reg[20]));
   AOI22_X1 i_0_2_622 (.A1(n_0_161), .A2(state[1]), .B1(i[31]), .B2(state[0]), 
      .ZN(n_0_2_420));
   INV_X1 i_0_2_623 (.A(n_0_2_420), .ZN(i_next_reg[31]));
   AOI22_X1 i_0_2_624 (.A1(n_0_160), .A2(state[1]), .B1(i[30]), .B2(state[0]), 
      .ZN(n_0_2_421));
   INV_X1 i_0_2_625 (.A(n_0_2_421), .ZN(i_next_reg[30]));
   AOI22_X1 i_0_2_626 (.A1(n_0_159), .A2(state[1]), .B1(i[29]), .B2(state[0]), 
      .ZN(n_0_2_422));
   INV_X1 i_0_2_627 (.A(n_0_2_422), .ZN(i_next_reg[29]));
   AOI22_X1 i_0_2_628 (.A1(n_0_158), .A2(state[1]), .B1(i[28]), .B2(state[0]), 
      .ZN(n_0_2_423));
   INV_X1 i_0_2_629 (.A(n_0_2_423), .ZN(i_next_reg[28]));
   AOI22_X1 i_0_2_630 (.A1(n_0_157), .A2(state[1]), .B1(i[27]), .B2(state[0]), 
      .ZN(n_0_2_424));
   INV_X1 i_0_2_631 (.A(n_0_2_424), .ZN(i_next_reg[27]));
   AOI22_X1 i_0_2_632 (.A1(n_0_156), .A2(state[1]), .B1(i[26]), .B2(state[0]), 
      .ZN(n_0_2_425));
   INV_X1 i_0_2_633 (.A(n_0_2_425), .ZN(i_next_reg[26]));
   AOI22_X1 i_0_2_634 (.A1(n_0_155), .A2(state[1]), .B1(i[25]), .B2(state[0]), 
      .ZN(n_0_2_426));
   INV_X1 i_0_2_635 (.A(n_0_2_426), .ZN(i_next_reg[25]));
   AOI22_X1 i_0_2_636 (.A1(n_0_154), .A2(state[1]), .B1(i[24]), .B2(state[0]), 
      .ZN(n_0_2_427));
   INV_X1 i_0_2_637 (.A(n_0_2_427), .ZN(i_next_reg[24]));
   NAND4_X1 i_0_2_638 (.A1(n_0_2_420), .A2(n_0_2_421), .A3(n_0_2_422), .A4(
      n_0_2_423), .ZN(n_0_2_428));
   NAND4_X1 i_0_2_639 (.A1(n_0_2_424), .A2(n_0_2_425), .A3(n_0_2_426), .A4(
      n_0_2_427), .ZN(n_0_2_429));
   NOR2_X1 i_0_2_640 (.A1(n_0_2_428), .A2(n_0_2_429), .ZN(n_0_2_430));
   AOI22_X1 i_0_2_641 (.A1(n_0_153), .A2(state[1]), .B1(i[23]), .B2(state[0]), 
      .ZN(n_0_2_431));
   INV_X1 i_0_2_642 (.A(n_0_2_431), .ZN(i_next_reg[23]));
   AOI22_X1 i_0_2_643 (.A1(n_0_152), .A2(state[1]), .B1(i[22]), .B2(state[0]), 
      .ZN(n_0_2_432));
   INV_X1 i_0_2_644 (.A(n_0_2_432), .ZN(i_next_reg[22]));
   AOI22_X1 i_0_2_645 (.A1(n_0_151), .A2(state[1]), .B1(i[21]), .B2(state[0]), 
      .ZN(n_0_2_433));
   INV_X1 i_0_2_646 (.A(n_0_2_433), .ZN(i_next_reg[21]));
   NOR3_X1 i_0_2_647 (.A1(i_next_reg[23]), .A2(i_next_reg[22]), .A3(
      i_next_reg[21]), .ZN(n_0_2_434));
   AOI22_X1 i_0_2_648 (.A1(n_0_149), .A2(state[1]), .B1(i[19]), .B2(state[0]), 
      .ZN(n_0_2_435));
   INV_X1 i_0_2_649 (.A(n_0_2_435), .ZN(i_next_reg[19]));
   AOI22_X1 i_0_2_650 (.A1(n_0_148), .A2(state[1]), .B1(i[18]), .B2(state[0]), 
      .ZN(n_0_2_436));
   INV_X1 i_0_2_651 (.A(n_0_2_436), .ZN(i_next_reg[18]));
   AOI22_X1 i_0_2_652 (.A1(n_0_147), .A2(state[1]), .B1(i[17]), .B2(state[0]), 
      .ZN(n_0_2_437));
   INV_X1 i_0_2_653 (.A(n_0_2_437), .ZN(i_next_reg[17]));
   AOI22_X1 i_0_2_654 (.A1(n_0_146), .A2(state[1]), .B1(i[16]), .B2(state[0]), 
      .ZN(n_0_2_438));
   INV_X1 i_0_2_655 (.A(n_0_2_438), .ZN(i_next_reg[16]));
   NOR4_X1 i_0_2_656 (.A1(i_next_reg[19]), .A2(i_next_reg[18]), .A3(
      i_next_reg[17]), .A4(i_next_reg[16]), .ZN(n_0_2_439));
   NAND4_X1 i_0_2_657 (.A1(n_0_2_430), .A2(n_0_2_419), .A3(n_0_2_434), .A4(
      n_0_2_439), .ZN(n_0_2_440));
   AOI22_X1 i_0_2_658 (.A1(n_0_133), .A2(state[1]), .B1(i[3]), .B2(state[0]), 
      .ZN(n_0_2_441));
   NAND4_X1 i_0_2_659 (.A1(n_0_2_441), .A2(i_next_reg[2]), .A3(i_next_reg[1]), 
      .A4(i_next_reg[0]), .ZN(n_0_2_442));
   AOI22_X1 i_0_2_660 (.A1(n_0_141), .A2(state[1]), .B1(i[11]), .B2(state[0]), 
      .ZN(n_0_2_443));
   INV_X1 i_0_2_661 (.A(n_0_2_443), .ZN(i_next_reg[11]));
   AOI22_X1 i_0_2_662 (.A1(n_0_140), .A2(state[1]), .B1(i[10]), .B2(state[0]), 
      .ZN(n_0_2_444));
   INV_X1 i_0_2_663 (.A(n_0_2_444), .ZN(i_next_reg[10]));
   AOI22_X1 i_0_2_664 (.A1(n_0_139), .A2(state[1]), .B1(i[9]), .B2(state[0]), 
      .ZN(n_0_2_445));
   INV_X1 i_0_2_665 (.A(n_0_2_445), .ZN(i_next_reg[9]));
   NOR3_X1 i_0_2_666 (.A1(i_next_reg[11]), .A2(i_next_reg[10]), .A3(
      i_next_reg[9]), .ZN(n_0_2_446));
   AOI22_X1 i_0_2_667 (.A1(n_0_145), .A2(state[1]), .B1(i[15]), .B2(state[0]), 
      .ZN(n_0_2_447));
   INV_X1 i_0_2_668 (.A(n_0_2_447), .ZN(i_next_reg[15]));
   AOI22_X1 i_0_2_669 (.A1(n_0_144), .A2(state[1]), .B1(i[14]), .B2(state[0]), 
      .ZN(n_0_2_448));
   INV_X1 i_0_2_670 (.A(n_0_2_448), .ZN(i_next_reg[14]));
   AOI22_X1 i_0_2_671 (.A1(n_0_143), .A2(state[1]), .B1(i[13]), .B2(state[0]), 
      .ZN(n_0_2_449));
   INV_X1 i_0_2_672 (.A(n_0_2_449), .ZN(i_next_reg[13]));
   NOR3_X1 i_0_2_673 (.A1(i_next_reg[15]), .A2(i_next_reg[14]), .A3(
      i_next_reg[13]), .ZN(n_0_2_450));
   NAND4_X1 i_0_2_674 (.A1(n_0_2_446), .A2(n_0_2_450), .A3(n_0_2_417), .A4(
      n_0_2_418), .ZN(n_0_2_451));
   AOI22_X1 i_0_2_675 (.A1(i[4]), .A2(state[0]), .B1(n_0_134), .B2(state[1]), 
      .ZN(n_0_2_452));
   INV_X1 i_0_2_676 (.A(n_0_2_452), .ZN(i_next_reg[4]));
   NAND4_X1 i_0_2_677 (.A1(i_next_reg[4]), .A2(n_0_2_414), .A3(n_0_2_415), 
      .A4(n_0_2_416), .ZN(n_0_2_453));
   NOR4_X1 i_0_2_678 (.A1(n_0_2_440), .A2(n_0_2_442), .A3(n_0_2_451), .A4(
      n_0_2_453), .ZN(n_0_2_454));
   INV_X1 i_0_2_679 (.A(enbl), .ZN(n_0_2_455));
   NOR2_X1 i_0_2_680 (.A1(n_0_2_454), .A2(n_0_2_455), .ZN(n_0_2_456));
   AOI22_X1 i_0_2_681 (.A1(n_0_2_456), .A2(out_sig[0]), .B1(n_0_2_454), .B2(
      quotient[0]), .ZN(n_0_2_457));
   NOR2_X1 i_0_2_682 (.A1(n_0_2_457), .A2(n_0_2_0), .ZN(n_0_299));
   XOR2_X1 i_0_2_683 (.A(in_a[15]), .B(in_b[15]), .Z(n_0_2_458));
   AND2_X1 i_0_2_684 (.A1(n_0_2_454), .A2(n_0_2_458), .ZN(n_0_2_459));
   INV_X1 i_0_2_685 (.A(n_0_2_454), .ZN(n_0_2_460));
   NOR2_X1 i_0_2_686 (.A1(n_0_2_460), .A2(n_0_2_458), .ZN(n_0_2_461));
   AOI222_X1 i_0_2_687 (.A1(n_0_2_456), .A2(out_sig[1]), .B1(n_0_2_459), 
      .B2(n_0_162), .C1(n_0_2_461), .C2(quotient[1]), .ZN(n_0_2_462));
   NOR2_X1 i_0_2_688 (.A1(n_0_2_462), .A2(n_0_2_0), .ZN(n_0_300));
   AOI222_X1 i_0_2_689 (.A1(n_0_2_456), .A2(out_sig[2]), .B1(n_0_2_459), 
      .B2(n_0_163), .C1(n_0_2_461), .C2(quotient[2]), .ZN(n_0_2_463));
   NOR2_X1 i_0_2_690 (.A1(n_0_2_463), .A2(n_0_2_0), .ZN(n_0_301));
   AOI222_X1 i_0_2_691 (.A1(n_0_2_456), .A2(out_sig[3]), .B1(n_0_2_459), 
      .B2(n_0_164), .C1(n_0_2_461), .C2(quotient[3]), .ZN(n_0_2_464));
   NOR2_X1 i_0_2_692 (.A1(n_0_2_464), .A2(n_0_2_0), .ZN(n_0_302));
   AOI222_X1 i_0_2_693 (.A1(n_0_2_456), .A2(out_sig[4]), .B1(n_0_2_459), 
      .B2(n_0_165), .C1(n_0_2_461), .C2(quotient[4]), .ZN(n_0_2_465));
   NOR2_X1 i_0_2_694 (.A1(n_0_2_465), .A2(n_0_2_0), .ZN(n_0_303));
   AOI222_X1 i_0_2_695 (.A1(n_0_2_456), .A2(out_sig[5]), .B1(n_0_2_459), 
      .B2(n_0_166), .C1(n_0_2_461), .C2(quotient[5]), .ZN(n_0_2_466));
   NOR2_X1 i_0_2_696 (.A1(n_0_2_466), .A2(n_0_2_0), .ZN(n_0_304));
   AOI222_X1 i_0_2_697 (.A1(n_0_2_456), .A2(out_sig[6]), .B1(n_0_2_459), 
      .B2(n_0_167), .C1(n_0_2_461), .C2(quotient[6]), .ZN(n_0_2_467));
   NOR2_X1 i_0_2_698 (.A1(n_0_2_467), .A2(n_0_2_0), .ZN(n_0_305));
   AOI222_X1 i_0_2_699 (.A1(n_0_2_456), .A2(out_sig[7]), .B1(n_0_2_459), 
      .B2(n_0_168), .C1(n_0_2_461), .C2(quotient[7]), .ZN(n_0_2_468));
   NOR2_X1 i_0_2_700 (.A1(n_0_2_468), .A2(n_0_2_0), .ZN(n_0_306));
   AOI222_X1 i_0_2_701 (.A1(n_0_2_456), .A2(out_sig[8]), .B1(n_0_2_459), 
      .B2(n_0_169), .C1(n_0_2_461), .C2(quotient[8]), .ZN(n_0_2_469));
   NOR2_X1 i_0_2_702 (.A1(n_0_2_469), .A2(n_0_2_0), .ZN(n_0_307));
   AOI222_X1 i_0_2_703 (.A1(n_0_2_456), .A2(out_sig[9]), .B1(n_0_2_459), 
      .B2(n_0_170), .C1(n_0_2_461), .C2(quotient[9]), .ZN(n_0_2_470));
   NOR2_X1 i_0_2_704 (.A1(n_0_2_470), .A2(n_0_2_0), .ZN(n_0_308));
   AOI222_X1 i_0_2_705 (.A1(n_0_2_456), .A2(out_sig[10]), .B1(n_0_2_459), 
      .B2(n_0_171), .C1(n_0_2_461), .C2(quotient[10]), .ZN(n_0_2_471));
   NOR2_X1 i_0_2_706 (.A1(n_0_2_471), .A2(n_0_2_0), .ZN(n_0_309));
   AOI222_X1 i_0_2_707 (.A1(n_0_2_456), .A2(out_sig[11]), .B1(n_0_2_459), 
      .B2(n_0_172), .C1(n_0_2_461), .C2(quotient[11]), .ZN(n_0_2_472));
   NOR2_X1 i_0_2_708 (.A1(n_0_2_472), .A2(n_0_2_0), .ZN(n_0_310));
   AOI222_X1 i_0_2_709 (.A1(n_0_2_456), .A2(out_sig[12]), .B1(n_0_2_459), 
      .B2(n_0_173), .C1(n_0_2_461), .C2(quotient[12]), .ZN(n_0_2_473));
   NOR2_X1 i_0_2_710 (.A1(n_0_2_473), .A2(n_0_2_0), .ZN(n_0_311));
   AOI222_X1 i_0_2_711 (.A1(n_0_2_456), .A2(out_sig[13]), .B1(n_0_2_459), 
      .B2(n_0_174), .C1(n_0_2_461), .C2(quotient[13]), .ZN(n_0_2_474));
   NOR2_X1 i_0_2_712 (.A1(n_0_2_474), .A2(n_0_2_0), .ZN(n_0_312));
   AOI222_X1 i_0_2_713 (.A1(n_0_2_456), .A2(out_sig[14]), .B1(n_0_2_459), 
      .B2(n_0_175), .C1(n_0_2_461), .C2(quotient[14]), .ZN(n_0_2_475));
   NOR2_X1 i_0_2_714 (.A1(n_0_2_475), .A2(n_0_2_0), .ZN(n_0_313));
   AOI222_X1 i_0_2_715 (.A1(n_0_2_456), .A2(out_sig[15]), .B1(n_0_2_459), 
      .B2(n_0_176), .C1(n_0_2_461), .C2(quotient[15]), .ZN(n_0_2_476));
   NOR2_X1 i_0_2_716 (.A1(n_0_2_476), .A2(n_0_2_0), .ZN(n_0_314));
   AOI222_X1 i_0_2_717 (.A1(n_0_2_456), .A2(out_sig[16]), .B1(n_0_2_459), 
      .B2(n_0_177), .C1(n_0_2_461), .C2(quotient[16]), .ZN(n_0_2_477));
   NOR2_X1 i_0_2_718 (.A1(n_0_2_477), .A2(n_0_2_0), .ZN(n_0_315));
   AOI222_X1 i_0_2_719 (.A1(n_0_2_456), .A2(out_sig[17]), .B1(n_0_2_459), 
      .B2(n_0_178), .C1(n_0_2_461), .C2(quotient[17]), .ZN(n_0_2_478));
   NOR2_X1 i_0_2_720 (.A1(n_0_2_478), .A2(n_0_2_0), .ZN(n_0_316));
   AOI222_X1 i_0_2_721 (.A1(n_0_2_456), .A2(out_sig[18]), .B1(n_0_2_459), 
      .B2(n_0_179), .C1(n_0_2_461), .C2(quotient[18]), .ZN(n_0_2_479));
   NOR2_X1 i_0_2_722 (.A1(n_0_2_479), .A2(n_0_2_0), .ZN(n_0_317));
   AOI222_X1 i_0_2_723 (.A1(n_0_2_456), .A2(out_sig[19]), .B1(n_0_2_459), 
      .B2(n_0_180), .C1(n_0_2_461), .C2(quotient[19]), .ZN(n_0_2_480));
   NOR2_X1 i_0_2_724 (.A1(n_0_2_480), .A2(n_0_2_0), .ZN(n_0_318));
   AOI222_X1 i_0_2_725 (.A1(n_0_2_456), .A2(out_sig[20]), .B1(n_0_2_459), 
      .B2(n_0_181), .C1(n_0_2_461), .C2(quotient[20]), .ZN(n_0_2_481));
   NOR2_X1 i_0_2_726 (.A1(n_0_2_481), .A2(n_0_2_0), .ZN(n_0_319));
   AOI222_X1 i_0_2_727 (.A1(n_0_2_456), .A2(out_sig[21]), .B1(n_0_2_459), 
      .B2(n_0_182), .C1(n_0_2_461), .C2(quotient[21]), .ZN(n_0_2_482));
   NOR2_X1 i_0_2_728 (.A1(n_0_2_482), .A2(n_0_2_0), .ZN(n_0_320));
   AOI222_X1 i_0_2_729 (.A1(n_0_2_456), .A2(out_sig[22]), .B1(n_0_2_459), 
      .B2(n_0_183), .C1(n_0_2_461), .C2(quotient[22]), .ZN(n_0_2_483));
   NOR2_X1 i_0_2_730 (.A1(n_0_2_483), .A2(n_0_2_0), .ZN(n_0_321));
   AOI222_X1 i_0_2_731 (.A1(n_0_2_456), .A2(out_sig[23]), .B1(n_0_2_459), 
      .B2(n_0_184), .C1(n_0_2_461), .C2(quotient[23]), .ZN(n_0_2_484));
   NOR2_X1 i_0_2_732 (.A1(n_0_2_484), .A2(n_0_2_0), .ZN(n_0_322));
   AOI222_X1 i_0_2_733 (.A1(n_0_2_456), .A2(out_sig[24]), .B1(n_0_2_459), 
      .B2(n_0_185), .C1(n_0_2_461), .C2(quotient[24]), .ZN(n_0_2_485));
   NOR2_X1 i_0_2_734 (.A1(n_0_2_485), .A2(n_0_2_0), .ZN(n_0_323));
   AOI222_X1 i_0_2_735 (.A1(n_0_2_456), .A2(out_sig[25]), .B1(n_0_2_459), 
      .B2(n_0_186), .C1(n_0_2_461), .C2(quotient[25]), .ZN(n_0_2_486));
   NOR2_X1 i_0_2_736 (.A1(n_0_2_486), .A2(n_0_2_0), .ZN(n_0_324));
   AOI222_X1 i_0_2_737 (.A1(n_0_2_456), .A2(out_sig[26]), .B1(n_0_2_459), 
      .B2(n_0_187), .C1(n_0_2_461), .C2(quotient[26]), .ZN(n_0_2_487));
   NOR2_X1 i_0_2_738 (.A1(n_0_2_487), .A2(n_0_2_0), .ZN(n_0_325));
   AOI222_X1 i_0_2_739 (.A1(n_0_2_456), .A2(out_sig[27]), .B1(n_0_2_459), 
      .B2(n_0_188), .C1(n_0_2_461), .C2(quotient[27]), .ZN(n_0_2_488));
   NOR2_X1 i_0_2_740 (.A1(n_0_2_488), .A2(n_0_2_0), .ZN(n_0_326));
   AOI222_X1 i_0_2_741 (.A1(n_0_2_456), .A2(out_sig[28]), .B1(n_0_2_459), 
      .B2(n_0_189), .C1(n_0_2_461), .C2(quotient[28]), .ZN(n_0_2_489));
   NOR2_X1 i_0_2_742 (.A1(n_0_2_489), .A2(n_0_2_0), .ZN(n_0_327));
   AOI222_X1 i_0_2_743 (.A1(n_0_2_456), .A2(out_sig[29]), .B1(n_0_2_459), 
      .B2(n_0_190), .C1(n_0_2_461), .C2(quotient[29]), .ZN(n_0_2_490));
   NOR2_X1 i_0_2_744 (.A1(n_0_2_490), .A2(n_0_2_0), .ZN(n_0_328));
   AOI222_X1 i_0_2_745 (.A1(n_0_2_456), .A2(out_sig[30]), .B1(n_0_2_459), 
      .B2(n_0_191), .C1(n_0_2_461), .C2(quotient[30]), .ZN(n_0_2_491));
   NOR2_X1 i_0_2_746 (.A1(n_0_2_491), .A2(n_0_2_0), .ZN(n_0_329));
   AOI222_X1 i_0_2_747 (.A1(n_0_2_456), .A2(out_sig[31]), .B1(n_0_2_459), 
      .B2(n_0_192), .C1(n_0_2_461), .C2(quotient[31]), .ZN(n_0_2_492));
   NOR2_X1 i_0_2_748 (.A1(n_0_2_492), .A2(n_0_2_0), .ZN(n_0_330));
   AOI222_X1 i_0_2_749 (.A1(n_0_2_456), .A2(out_sig[32]), .B1(n_0_2_459), 
      .B2(n_0_193), .C1(n_0_2_461), .C2(quotient[32]), .ZN(n_0_2_493));
   NOR2_X1 i_0_2_750 (.A1(n_0_2_493), .A2(n_0_2_0), .ZN(n_0_331));
   AOI222_X1 i_0_2_751 (.A1(n_0_2_456), .A2(out_sig[33]), .B1(n_0_2_459), 
      .B2(n_0_194), .C1(n_0_2_461), .C2(quotient[33]), .ZN(n_0_2_494));
   NOR2_X1 i_0_2_752 (.A1(n_0_2_494), .A2(n_0_2_0), .ZN(n_0_332));
   AOI222_X1 i_0_2_753 (.A1(n_0_2_456), .A2(out_sig[34]), .B1(n_0_2_459), 
      .B2(n_0_195), .C1(n_0_2_461), .C2(quotient[34]), .ZN(n_0_2_495));
   NOR2_X1 i_0_2_754 (.A1(n_0_2_495), .A2(n_0_2_0), .ZN(n_0_333));
   AOI222_X1 i_0_2_755 (.A1(n_0_2_456), .A2(out_sig[35]), .B1(n_0_2_459), 
      .B2(n_0_196), .C1(n_0_2_461), .C2(quotient[35]), .ZN(n_0_2_496));
   NOR2_X1 i_0_2_756 (.A1(n_0_2_496), .A2(n_0_2_0), .ZN(n_0_334));
   AOI222_X1 i_0_2_757 (.A1(n_0_2_456), .A2(out_sig[36]), .B1(n_0_2_459), 
      .B2(n_0_197), .C1(n_0_2_461), .C2(quotient[36]), .ZN(n_0_2_497));
   NOR2_X1 i_0_2_758 (.A1(n_0_2_497), .A2(n_0_2_0), .ZN(n_0_335));
   AOI222_X1 i_0_2_759 (.A1(n_0_2_456), .A2(out_sig[37]), .B1(n_0_2_459), 
      .B2(n_0_198), .C1(n_0_2_461), .C2(quotient[37]), .ZN(n_0_2_498));
   NOR2_X1 i_0_2_760 (.A1(n_0_2_498), .A2(n_0_2_0), .ZN(n_0_336));
   AOI222_X1 i_0_2_761 (.A1(n_0_2_456), .A2(out_sig[38]), .B1(n_0_2_459), 
      .B2(n_0_199), .C1(n_0_2_461), .C2(quotient[38]), .ZN(n_0_2_499));
   NOR2_X1 i_0_2_762 (.A1(n_0_2_499), .A2(n_0_2_0), .ZN(n_0_337));
   AOI222_X1 i_0_2_763 (.A1(n_0_2_456), .A2(out_sig[39]), .B1(n_0_2_459), 
      .B2(n_0_200), .C1(n_0_2_461), .C2(quotient[39]), .ZN(n_0_2_500));
   NOR2_X1 i_0_2_764 (.A1(n_0_2_500), .A2(n_0_2_0), .ZN(n_0_338));
   AOI222_X1 i_0_2_765 (.A1(n_0_2_456), .A2(out_sig[40]), .B1(n_0_2_459), 
      .B2(n_0_201), .C1(n_0_2_461), .C2(quotient[40]), .ZN(n_0_2_501));
   NOR2_X1 i_0_2_766 (.A1(n_0_2_501), .A2(n_0_2_0), .ZN(n_0_339));
   AOI222_X1 i_0_2_767 (.A1(n_0_2_456), .A2(out_sig[41]), .B1(n_0_2_459), 
      .B2(n_0_202), .C1(n_0_2_461), .C2(quotient[41]), .ZN(n_0_2_502));
   NOR2_X1 i_0_2_768 (.A1(n_0_2_502), .A2(n_0_2_0), .ZN(n_0_340));
   AOI222_X1 i_0_2_769 (.A1(n_0_2_456), .A2(out_sig[42]), .B1(n_0_2_459), 
      .B2(n_0_203), .C1(n_0_2_461), .C2(quotient[42]), .ZN(n_0_2_503));
   NOR2_X1 i_0_2_770 (.A1(n_0_2_503), .A2(n_0_2_0), .ZN(n_0_341));
   AOI222_X1 i_0_2_771 (.A1(n_0_2_456), .A2(out_sig[43]), .B1(n_0_2_459), 
      .B2(n_0_204), .C1(n_0_2_461), .C2(quotient[43]), .ZN(n_0_2_504));
   NOR2_X1 i_0_2_772 (.A1(n_0_2_504), .A2(n_0_2_0), .ZN(n_0_342));
   AOI222_X1 i_0_2_773 (.A1(n_0_2_456), .A2(out_sig[44]), .B1(n_0_2_459), 
      .B2(n_0_205), .C1(n_0_2_461), .C2(quotient[44]), .ZN(n_0_2_505));
   NOR2_X1 i_0_2_774 (.A1(n_0_2_505), .A2(n_0_2_0), .ZN(n_0_343));
   AOI222_X1 i_0_2_775 (.A1(n_0_2_456), .A2(out_sig[45]), .B1(n_0_2_459), 
      .B2(n_0_206), .C1(n_0_2_461), .C2(quotient[45]), .ZN(n_0_2_506));
   NOR2_X1 i_0_2_776 (.A1(n_0_2_506), .A2(n_0_2_0), .ZN(n_0_344));
   AOI222_X1 i_0_2_777 (.A1(n_0_2_456), .A2(out_sig[46]), .B1(n_0_2_459), 
      .B2(n_0_207), .C1(n_0_2_461), .C2(quotient[46]), .ZN(n_0_2_507));
   NOR2_X1 i_0_2_778 (.A1(n_0_2_507), .A2(n_0_2_0), .ZN(n_0_345));
   AOI222_X1 i_0_2_779 (.A1(n_0_2_456), .A2(out_sig[47]), .B1(n_0_2_459), 
      .B2(n_0_208), .C1(n_0_2_461), .C2(quotient[47]), .ZN(n_0_2_508));
   NOR2_X1 i_0_2_780 (.A1(n_0_2_508), .A2(n_0_2_0), .ZN(n_0_346));
   AOI222_X1 i_0_2_781 (.A1(n_0_2_456), .A2(out_sig[48]), .B1(n_0_2_459), 
      .B2(n_0_209), .C1(n_0_2_461), .C2(quotient[48]), .ZN(n_0_2_509));
   NOR2_X1 i_0_2_782 (.A1(n_0_2_509), .A2(n_0_2_0), .ZN(n_0_347));
   AOI222_X1 i_0_2_783 (.A1(n_0_2_456), .A2(out_sig[49]), .B1(n_0_2_459), 
      .B2(n_0_210), .C1(n_0_2_461), .C2(quotient[49]), .ZN(n_0_2_510));
   NOR2_X1 i_0_2_784 (.A1(n_0_2_510), .A2(n_0_2_0), .ZN(n_0_348));
   AOI222_X1 i_0_2_785 (.A1(n_0_2_456), .A2(out_sig[50]), .B1(n_0_2_459), 
      .B2(n_0_211), .C1(n_0_2_461), .C2(quotient[50]), .ZN(n_0_2_511));
   NOR2_X1 i_0_2_786 (.A1(n_0_2_511), .A2(n_0_2_0), .ZN(n_0_349));
   AOI222_X1 i_0_2_787 (.A1(n_0_2_456), .A2(out_sig[51]), .B1(n_0_2_459), 
      .B2(n_0_212), .C1(n_0_2_461), .C2(quotient[51]), .ZN(n_0_2_512));
   NOR2_X1 i_0_2_788 (.A1(n_0_2_512), .A2(n_0_2_0), .ZN(n_0_350));
   AOI222_X1 i_0_2_789 (.A1(n_0_2_456), .A2(out_sig[52]), .B1(n_0_2_459), 
      .B2(n_0_213), .C1(n_0_2_461), .C2(quotient[52]), .ZN(n_0_2_513));
   NOR2_X1 i_0_2_790 (.A1(n_0_2_513), .A2(n_0_2_0), .ZN(n_0_351));
   AOI222_X1 i_0_2_791 (.A1(n_0_2_456), .A2(out_sig[53]), .B1(n_0_2_459), 
      .B2(n_0_214), .C1(n_0_2_461), .C2(quotient[53]), .ZN(n_0_2_514));
   NOR2_X1 i_0_2_792 (.A1(n_0_2_514), .A2(n_0_2_0), .ZN(n_0_352));
   AOI222_X1 i_0_2_793 (.A1(n_0_2_456), .A2(out_sig[54]), .B1(n_0_2_459), 
      .B2(n_0_215), .C1(n_0_2_461), .C2(quotient[54]), .ZN(n_0_2_515));
   NOR2_X1 i_0_2_794 (.A1(n_0_2_515), .A2(n_0_2_0), .ZN(n_0_353));
   AOI222_X1 i_0_2_795 (.A1(n_0_2_456), .A2(out_sig[55]), .B1(n_0_2_459), 
      .B2(n_0_216), .C1(n_0_2_461), .C2(quotient[55]), .ZN(n_0_2_516));
   NOR2_X1 i_0_2_796 (.A1(n_0_2_516), .A2(n_0_2_0), .ZN(n_0_354));
   AOI222_X1 i_0_2_797 (.A1(n_0_2_456), .A2(out_sig[56]), .B1(n_0_2_459), 
      .B2(n_0_218), .C1(n_0_2_461), .C2(quotient[56]), .ZN(n_0_2_517));
   NOR2_X1 i_0_2_798 (.A1(n_0_2_517), .A2(n_0_2_0), .ZN(n_0_355));
   AOI222_X1 i_0_2_799 (.A1(n_0_2_456), .A2(out_sig[57]), .B1(n_0_2_459), 
      .B2(n_0_219), .C1(n_0_2_461), .C2(quotient[57]), .ZN(n_0_2_518));
   NOR2_X1 i_0_2_800 (.A1(n_0_2_518), .A2(n_0_2_0), .ZN(n_0_356));
   AOI222_X1 i_0_2_801 (.A1(n_0_2_456), .A2(out_sig[58]), .B1(n_0_2_459), 
      .B2(n_0_220), .C1(n_0_2_461), .C2(quotient[58]), .ZN(n_0_2_519));
   NOR2_X1 i_0_2_802 (.A1(n_0_2_519), .A2(n_0_2_0), .ZN(n_0_357));
   AOI222_X1 i_0_2_803 (.A1(n_0_2_456), .A2(out_sig[59]), .B1(n_0_2_459), 
      .B2(n_0_221), .C1(n_0_2_461), .C2(quotient[59]), .ZN(n_0_2_520));
   NOR2_X1 i_0_2_804 (.A1(n_0_2_520), .A2(n_0_2_0), .ZN(n_0_358));
   AOI222_X1 i_0_2_805 (.A1(n_0_2_456), .A2(out_sig[60]), .B1(n_0_2_459), 
      .B2(n_0_222), .C1(n_0_2_461), .C2(quotient[60]), .ZN(n_0_2_521));
   NOR2_X1 i_0_2_806 (.A1(n_0_2_521), .A2(n_0_2_0), .ZN(n_0_359));
   AOI222_X1 i_0_2_807 (.A1(n_0_2_456), .A2(out_sig[61]), .B1(n_0_2_459), 
      .B2(n_0_223), .C1(n_0_2_461), .C2(quotient[61]), .ZN(n_0_2_522));
   NOR2_X1 i_0_2_808 (.A1(n_0_2_522), .A2(n_0_2_0), .ZN(n_0_360));
   AOI222_X1 i_0_2_809 (.A1(n_0_2_456), .A2(out_sig[62]), .B1(n_0_2_459), 
      .B2(n_0_224), .C1(n_0_2_461), .C2(quotient[62]), .ZN(n_0_2_523));
   NOR2_X1 i_0_2_810 (.A1(n_0_2_523), .A2(n_0_2_0), .ZN(n_0_361));
   AOI222_X1 i_0_2_811 (.A1(n_0_2_456), .A2(out_sig[63]), .B1(n_0_2_459), 
      .B2(n_0_225), .C1(n_0_2_461), .C2(quotient[63]), .ZN(n_0_2_524));
   NOR2_X1 i_0_2_812 (.A1(n_0_2_524), .A2(n_0_2_0), .ZN(n_0_362));
   NOR4_X1 i_0_2_813 (.A1(in_b[11]), .A2(in_b[10]), .A3(in_b[9]), .A4(in_b[8]), 
      .ZN(n_0_2_525));
   NOR4_X1 i_0_2_814 (.A1(in_b[15]), .A2(in_b[14]), .A3(in_b[13]), .A4(in_b[12]), 
      .ZN(n_0_2_526));
   NOR4_X1 i_0_2_815 (.A1(in_b[7]), .A2(in_b[6]), .A3(in_b[5]), .A4(in_b[4]), 
      .ZN(n_0_2_527));
   NOR4_X1 i_0_2_816 (.A1(in_b[3]), .A2(in_b[2]), .A3(in_b[1]), .A4(in_b[0]), 
      .ZN(n_0_2_528));
   NAND4_X1 i_0_2_817 (.A1(n_0_2_525), .A2(n_0_2_526), .A3(n_0_2_527), .A4(
      n_0_2_528), .ZN(n_0_2_529));
   NOR4_X1 i_0_2_818 (.A1(in_b[27]), .A2(in_b[26]), .A3(in_b[25]), .A4(in_b[24]), 
      .ZN(n_0_2_530));
   NOR4_X1 i_0_2_819 (.A1(in_b[31]), .A2(in_b[30]), .A3(in_b[29]), .A4(in_b[28]), 
      .ZN(n_0_2_531));
   NOR4_X1 i_0_2_820 (.A1(in_b[23]), .A2(in_b[22]), .A3(in_b[21]), .A4(in_b[20]), 
      .ZN(n_0_2_532));
   NOR4_X1 i_0_2_821 (.A1(in_b[19]), .A2(in_b[18]), .A3(in_b[17]), .A4(in_b[16]), 
      .ZN(n_0_2_533));
   NAND4_X1 i_0_2_822 (.A1(n_0_2_530), .A2(n_0_2_531), .A3(n_0_2_532), .A4(
      n_0_2_533), .ZN(n_0_2_534));
   OR2_X1 i_0_2_823 (.A1(n_0_2_529), .A2(n_0_2_534), .ZN(n_0_2_535));
   NOR4_X1 i_0_2_824 (.A1(in_b[43]), .A2(in_b[42]), .A3(in_b[41]), .A4(in_b[40]), 
      .ZN(n_0_2_536));
   NOR4_X1 i_0_2_825 (.A1(in_b[47]), .A2(in_b[46]), .A3(in_b[45]), .A4(in_b[44]), 
      .ZN(n_0_2_537));
   NOR4_X1 i_0_2_826 (.A1(in_b[35]), .A2(in_b[34]), .A3(in_b[33]), .A4(in_b[32]), 
      .ZN(n_0_2_538));
   NOR4_X1 i_0_2_827 (.A1(in_b[39]), .A2(in_b[38]), .A3(in_b[37]), .A4(in_b[36]), 
      .ZN(n_0_2_539));
   NAND4_X1 i_0_2_828 (.A1(n_0_2_536), .A2(n_0_2_537), .A3(n_0_2_538), .A4(
      n_0_2_539), .ZN(n_0_2_540));
   OR4_X1 i_0_2_829 (.A1(in_b[51]), .A2(in_b[50]), .A3(in_b[49]), .A4(in_b[48]), 
      .ZN(n_0_2_541));
   NOR4_X1 i_0_2_830 (.A1(n_0_2_541), .A2(in_b[55]), .A3(in_b[54]), .A4(in_b[53]), 
      .ZN(n_0_2_542));
   NOR4_X1 i_0_2_831 (.A1(in_b[59]), .A2(in_b[56]), .A3(in_b[61]), .A4(in_b[60]), 
      .ZN(n_0_2_543));
   NOR4_X1 i_0_2_832 (.A1(in_b[63]), .A2(in_b[62]), .A3(in_b[58]), .A4(in_b[57]), 
      .ZN(n_0_2_544));
   NAND3_X1 i_0_2_833 (.A1(n_0_2_542), .A2(n_0_2_543), .A3(n_0_2_544), .ZN(
      n_0_2_545));
   NOR4_X1 i_0_2_834 (.A1(n_0_2_535), .A2(n_0_2_540), .A3(n_0_2_545), .A4(
      in_b[52]), .ZN(n_0_2_546));
   AOI22_X1 i_0_2_835 (.A1(n_0_2_456), .A2(div_by_zero_sig), .B1(n_0_2_454), 
      .B2(n_0_2_546), .ZN(n_0_2_547));
   NOR2_X1 i_0_2_836 (.A1(n_0_2_547), .A2(n_0_2_0), .ZN(n_0_363));
   OR4_X1 i_0_2_837 (.A1(quotient[22]), .A2(quotient[21]), .A3(quotient[20]), 
      .A4(quotient[19]), .ZN(n_0_2_548));
   OR4_X1 i_0_2_838 (.A1(n_0_2_548), .A2(quotient[18]), .A3(quotient[17]), 
      .A4(quotient[16]), .ZN(n_0_2_549));
   AOI22_X1 i_0_2_839 (.A1(n_0_2_456), .A2(ovfl_sig), .B1(n_0_2_454), .B2(
      n_0_2_549), .ZN(n_0_2_550));
   NOR2_X1 i_0_2_840 (.A1(n_0_2_550), .A2(n_0_2_0), .ZN(n_0_364));
   INV_X1 i_0_2_841 (.A(n_0_2_524), .ZN(out_c[63]));
   INV_X1 i_0_2_842 (.A(n_0_2_457), .ZN(out_c[0]));
   INV_X1 i_0_2_843 (.A(n_0_2_523), .ZN(out_c[62]));
   INV_X1 i_0_2_844 (.A(n_0_2_522), .ZN(out_c[61]));
   INV_X1 i_0_2_845 (.A(n_0_2_519), .ZN(out_c[58]));
   INV_X1 i_0_2_846 (.A(n_0_2_518), .ZN(out_c[57]));
   INV_X1 i_0_2_847 (.A(n_0_2_521), .ZN(out_c[60]));
   INV_X1 i_0_2_848 (.A(n_0_2_520), .ZN(out_c[59]));
   INV_X1 i_0_2_849 (.A(n_0_2_511), .ZN(out_c[50]));
   INV_X1 i_0_2_850 (.A(n_0_2_510), .ZN(out_c[49]));
   INV_X1 i_0_2_851 (.A(n_0_2_513), .ZN(out_c[52]));
   INV_X1 i_0_2_852 (.A(n_0_2_512), .ZN(out_c[51]));
   INV_X1 i_0_2_853 (.A(n_0_2_515), .ZN(out_c[54]));
   INV_X1 i_0_2_854 (.A(n_0_2_514), .ZN(out_c[53]));
   INV_X1 i_0_2_855 (.A(n_0_2_517), .ZN(out_c[56]));
   INV_X1 i_0_2_856 (.A(n_0_2_516), .ZN(out_c[55]));
   INV_X1 i_0_2_857 (.A(n_0_2_464), .ZN(out_c[3]));
   INV_X1 i_0_2_858 (.A(n_0_2_466), .ZN(out_c[5]));
   INV_X1 i_0_2_859 (.A(n_0_2_465), .ZN(out_c[4]));
   INV_X1 i_0_2_860 (.A(n_0_2_468), .ZN(out_c[7]));
   INV_X1 i_0_2_861 (.A(n_0_2_467), .ZN(out_c[6]));
   INV_X1 i_0_2_862 (.A(n_0_2_472), .ZN(out_c[11]));
   INV_X1 i_0_2_863 (.A(n_0_2_471), .ZN(out_c[10]));
   INV_X1 i_0_2_864 (.A(n_0_2_470), .ZN(out_c[9]));
   INV_X1 i_0_2_865 (.A(n_0_2_469), .ZN(out_c[8]));
   INV_X1 i_0_2_866 (.A(n_0_2_481), .ZN(out_c[20]));
   INV_X1 i_0_2_867 (.A(n_0_2_480), .ZN(out_c[19]));
   INV_X1 i_0_2_868 (.A(n_0_2_479), .ZN(out_c[18]));
   INV_X1 i_0_2_869 (.A(n_0_2_478), .ZN(out_c[17]));
   INV_X1 i_0_2_870 (.A(n_0_2_487), .ZN(out_c[26]));
   INV_X1 i_0_2_871 (.A(n_0_2_486), .ZN(out_c[25]));
   INV_X1 i_0_2_872 (.A(n_0_2_489), .ZN(out_c[28]));
   INV_X1 i_0_2_873 (.A(n_0_2_488), .ZN(out_c[27]));
   INV_X1 i_0_2_874 (.A(n_0_2_503), .ZN(out_c[42]));
   INV_X1 i_0_2_875 (.A(n_0_2_502), .ZN(out_c[41]));
   INV_X1 i_0_2_876 (.A(n_0_2_505), .ZN(out_c[44]));
   INV_X1 i_0_2_877 (.A(n_0_2_504), .ZN(out_c[43]));
   INV_X1 i_0_2_878 (.A(n_0_2_495), .ZN(out_c[34]));
   INV_X1 i_0_2_879 (.A(n_0_2_494), .ZN(out_c[33]));
   INV_X1 i_0_2_880 (.A(n_0_2_497), .ZN(out_c[36]));
   INV_X1 i_0_2_881 (.A(n_0_2_496), .ZN(out_c[35]));
   NOR4_X1 i_0_2_882 (.A1(out_c[33]), .A2(out_c[34]), .A3(out_c[35]), .A4(
      out_c[36]), .ZN(n_0_2_551));
   NAND3_X1 i_0_2_883 (.A1(n_0_2_551), .A2(n_0_2_498), .A3(n_0_2_501), .ZN(
      n_0_2_552));
   NAND4_X1 i_0_2_884 (.A1(n_0_2_499), .A2(n_0_2_500), .A3(n_0_2_506), .A4(
      n_0_2_509), .ZN(n_0_2_553));
   NOR2_X1 i_0_2_885 (.A1(n_0_2_552), .A2(n_0_2_553), .ZN(n_0_2_554));
   NOR4_X1 i_0_2_886 (.A1(out_c[41]), .A2(out_c[42]), .A3(out_c[43]), .A4(
      out_c[44]), .ZN(n_0_2_555));
   NAND4_X1 i_0_2_887 (.A1(n_0_2_554), .A2(n_0_2_507), .A3(n_0_2_508), .A4(
      n_0_2_555), .ZN(n_0_2_556));
   NOR4_X1 i_0_2_888 (.A1(out_c[17]), .A2(out_c[18]), .A3(out_c[19]), .A4(
      out_c[20]), .ZN(n_0_2_557));
   NAND3_X1 i_0_2_889 (.A1(n_0_2_557), .A2(n_0_2_483), .A3(n_0_2_484), .ZN(
      n_0_2_558));
   NAND4_X1 i_0_2_890 (.A1(n_0_2_482), .A2(n_0_2_485), .A3(n_0_2_491), .A4(
      n_0_2_492), .ZN(n_0_2_559));
   NOR4_X1 i_0_2_891 (.A1(out_c[25]), .A2(out_c[26]), .A3(out_c[27]), .A4(
      out_c[28]), .ZN(n_0_2_560));
   NAND3_X1 i_0_2_892 (.A1(n_0_2_560), .A2(n_0_2_490), .A3(n_0_2_493), .ZN(
      n_0_2_561));
   NOR4_X1 i_0_2_893 (.A1(n_0_2_556), .A2(n_0_2_558), .A3(n_0_2_559), .A4(
      n_0_2_561), .ZN(n_0_2_562));
   NOR4_X1 i_0_2_894 (.A1(out_c[63]), .A2(out_c[61]), .A3(out_c[62]), .A4(
      out_c[0]), .ZN(n_0_2_563));
   NAND4_X1 i_0_2_895 (.A1(n_0_2_518), .A2(n_0_2_519), .A3(n_0_2_520), .A4(
      n_0_2_521), .ZN(n_0_2_564));
   NAND4_X1 i_0_2_896 (.A1(n_0_2_510), .A2(n_0_2_511), .A3(n_0_2_512), .A4(
      n_0_2_513), .ZN(n_0_2_565));
   NAND4_X1 i_0_2_897 (.A1(n_0_2_514), .A2(n_0_2_515), .A3(n_0_2_516), .A4(
      n_0_2_517), .ZN(n_0_2_566));
   NOR3_X1 i_0_2_898 (.A1(n_0_2_564), .A2(n_0_2_565), .A3(n_0_2_566), .ZN(
      n_0_2_567));
   NOR4_X1 i_0_2_899 (.A1(out_c[8]), .A2(out_c[9]), .A3(out_c[10]), .A4(
      out_c[11]), .ZN(n_0_2_568));
   NAND3_X1 i_0_2_900 (.A1(n_0_2_568), .A2(n_0_2_474), .A3(n_0_2_475), .ZN(
      n_0_2_569));
   NOR4_X1 i_0_2_901 (.A1(out_c[4]), .A2(out_c[5]), .A3(out_c[6]), .A4(out_c[7]), 
      .ZN(n_0_2_570));
   NAND3_X1 i_0_2_902 (.A1(n_0_2_570), .A2(n_0_2_462), .A3(n_0_2_463), .ZN(
      n_0_2_571));
   NAND2_X1 i_0_2_903 (.A1(n_0_2_473), .A2(n_0_2_477), .ZN(n_0_2_572));
   NOR4_X1 i_0_2_904 (.A1(n_0_2_569), .A2(n_0_2_571), .A3(out_c[3]), .A4(
      n_0_2_572), .ZN(n_0_2_573));
   NAND4_X1 i_0_2_905 (.A1(n_0_2_562), .A2(n_0_2_563), .A3(n_0_2_567), .A4(
      n_0_2_573), .ZN(n_0_2_574));
   INV_X1 i_0_2_906 (.A(n_0_2_574), .ZN(n_0_2_575));
   INV_X1 i_0_2_907 (.A(n_0_2_476), .ZN(out_c[15]));
   NOR2_X1 i_0_2_908 (.A1(out_c[15]), .A2(n_0_2_460), .ZN(n_0_2_576));
   AOI22_X1 i_0_2_909 (.A1(n_0_2_575), .A2(n_0_2_576), .B1(n_0_2_456), .B2(
      zero_sig), .ZN(n_0_2_577));
   INV_X1 i_0_2_910 (.A(n_0_2_577), .ZN(zero));
   NOR2_X1 i_0_2_911 (.A1(n_0_2_577), .A2(n_0_2_0), .ZN(n_0_365));
   NAND2_X1 i_0_2_912 (.A1(n_0_2_454), .A2(state[1]), .ZN(n_0_2_578));
   OAI21_X1 i_0_2_913 (.A(n_0_2_578), .B1(enbl), .B2(n_0_298), .ZN(n_0_391));
   AOI22_X1 i_0_2_914 (.A1(n_0_2_574), .A2(n_0_2_576), .B1(n_0_2_456), .B2(
      posv_sig), .ZN(n_0_2_579));
   NOR2_X1 i_0_2_915 (.A1(n_0_2_579), .A2(n_0_2_0), .ZN(n_0_392));
   INV_X1 i_0_2_916 (.A(n_0_2_579), .ZN(posv));
   INV_X1 i_0_2_917 (.A(n_0_2_578), .ZN(n_0_2_580));
   INV_X1 i_0_2_918 (.A(done_sig), .ZN(n_0_2_581));
   OAI211_X1 i_0_2_919 (.A(n_0_2_347), .B(enbl), .C1(n_0_2_454), .C2(n_0_2_581), 
      .ZN(n_0_2_582));
   AOI21_X1 i_0_2_920 (.A(n_0_2_580), .B1(n_0_2_582), .B2(n_0_2_15), .ZN(
      state_next_reg[0]));
   INV_X1 i_0_2_921 (.A(n_0_2_462), .ZN(out_c[1]));
   INV_X1 i_0_2_922 (.A(n_0_2_463), .ZN(out_c[2]));
   INV_X1 i_0_2_923 (.A(n_0_2_473), .ZN(out_c[12]));
   INV_X1 i_0_2_924 (.A(n_0_2_474), .ZN(out_c[13]));
   INV_X1 i_0_2_925 (.A(n_0_2_475), .ZN(out_c[14]));
   INV_X1 i_0_2_926 (.A(n_0_2_477), .ZN(out_c[16]));
   INV_X1 i_0_2_927 (.A(n_0_2_482), .ZN(out_c[21]));
   INV_X1 i_0_2_928 (.A(n_0_2_483), .ZN(out_c[22]));
   INV_X1 i_0_2_929 (.A(n_0_2_484), .ZN(out_c[23]));
   INV_X1 i_0_2_930 (.A(n_0_2_485), .ZN(out_c[24]));
   INV_X1 i_0_2_931 (.A(n_0_2_490), .ZN(out_c[29]));
   INV_X1 i_0_2_932 (.A(n_0_2_491), .ZN(out_c[30]));
   INV_X1 i_0_2_933 (.A(n_0_2_492), .ZN(out_c[31]));
   INV_X1 i_0_2_934 (.A(n_0_2_493), .ZN(out_c[32]));
   INV_X1 i_0_2_935 (.A(n_0_2_498), .ZN(out_c[37]));
   INV_X1 i_0_2_936 (.A(n_0_2_499), .ZN(out_c[38]));
   INV_X1 i_0_2_937 (.A(n_0_2_500), .ZN(out_c[39]));
   INV_X1 i_0_2_938 (.A(n_0_2_501), .ZN(out_c[40]));
   INV_X1 i_0_2_939 (.A(n_0_2_506), .ZN(out_c[45]));
   INV_X1 i_0_2_940 (.A(n_0_2_507), .ZN(out_c[46]));
   INV_X1 i_0_2_941 (.A(n_0_2_508), .ZN(out_c[47]));
   INV_X1 i_0_2_942 (.A(n_0_2_509), .ZN(out_c[48]));
   OAI21_X1 i_0_2_943 (.A(n_0_2_460), .B1(n_0_2_455), .B2(n_0_2_581), .ZN(done));
   NAND2_X1 i_0_2_944 (.A1(n_0_2_547), .A2(n_0_2_550), .ZN(err));
   INV_X1 i_0_2_945 (.A(n_0_2_226), .ZN(b[63]));
   INV_X1 i_0_2_946 (.A(n_0_2_441), .ZN(i_next_reg[3]));
endmodule
