/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sat Apr 25 22:01:01 2020
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 3930312276 */

module datapath(in_b, p_0);
   input [22:0]in_b;
   output [22:0]p_0;

   XOR2_X1 i_0 (.A(in_b[1]), .B(in_b[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_20), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(in_b[2]), .B1(in_b[1]), .B2(in_b[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(in_b[3]), .B(n_20), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(in_b[4]), .B(n_19), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(in_b[5]), .B(n_18), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_17), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(in_b[6]), .B1(n_18), .B2(in_b[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(in_b[7]), .B(n_17), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(in_b[8]), .B(n_16), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_15), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(in_b[9]), .B1(n_16), .B2(in_b[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(in_b[10]), .B(n_15), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(in_b[11]), .B(n_14), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(in_b[12]), .B(n_13), .Z(p_0[12]));
   XOR2_X1 i_15 (.A(in_b[13]), .B(n_12), .Z(p_0[13]));
   XNOR2_X1 i_16 (.A(in_b[14]), .B(n_11), .ZN(p_0[14]));
   XNOR2_X1 i_17 (.A(in_b[15]), .B(n_10), .ZN(p_0[15]));
   XOR2_X1 i_18 (.A(in_b[16]), .B(n_9), .Z(p_0[16]));
   XOR2_X1 i_19 (.A(in_b[17]), .B(n_8), .Z(p_0[17]));
   XNOR2_X1 i_20 (.A(in_b[18]), .B(n_7), .ZN(p_0[18]));
   XNOR2_X1 i_21 (.A(in_b[19]), .B(n_6), .ZN(p_0[19]));
   XOR2_X1 i_22 (.A(in_b[20]), .B(n_5), .Z(p_0[20]));
   XNOR2_X1 i_23 (.A(in_b[21]), .B(n_4), .ZN(p_0[21]));
   XNOR2_X1 i_24 (.A(in_b[22]), .B(n_3), .ZN(p_0[22]));
   NOR3_X1 i_25 (.A1(n_5), .A2(in_b[20]), .A3(in_b[21]), .ZN(n_3));
   NOR2_X1 i_26 (.A1(n_5), .A2(in_b[20]), .ZN(n_4));
   NAND2_X1 i_27 (.A1(n_6), .A2(n_23), .ZN(n_5));
   NOR3_X1 i_28 (.A1(n_8), .A2(in_b[17]), .A3(in_b[18]), .ZN(n_6));
   NOR2_X1 i_29 (.A1(n_8), .A2(in_b[17]), .ZN(n_7));
   OR2_X1 i_30 (.A1(n_9), .A2(in_b[16]), .ZN(n_8));
   NAND2_X1 i_31 (.A1(n_10), .A2(n_22), .ZN(n_9));
   NOR3_X1 i_32 (.A1(n_12), .A2(in_b[13]), .A3(in_b[14]), .ZN(n_10));
   NOR2_X1 i_33 (.A1(n_12), .A2(in_b[13]), .ZN(n_11));
   OR2_X1 i_34 (.A1(n_13), .A2(in_b[12]), .ZN(n_12));
   NAND2_X1 i_35 (.A1(n_14), .A2(n_21), .ZN(n_13));
   NOR2_X1 i_36 (.A1(n_15), .A2(in_b[10]), .ZN(n_14));
   OR3_X1 i_37 (.A1(n_16), .A2(in_b[8]), .A3(in_b[9]), .ZN(n_15));
   OR2_X1 i_38 (.A1(n_17), .A2(in_b[7]), .ZN(n_16));
   OR3_X1 i_39 (.A1(n_18), .A2(in_b[5]), .A3(in_b[6]), .ZN(n_17));
   OR2_X1 i_40 (.A1(n_19), .A2(in_b[4]), .ZN(n_18));
   OR2_X1 i_41 (.A1(n_20), .A2(in_b[3]), .ZN(n_19));
   OR3_X1 i_42 (.A1(in_b[2]), .A2(in_b[1]), .A3(in_b[0]), .ZN(n_20));
   INV_X1 i_43 (.A(in_b[11]), .ZN(n_21));
   INV_X1 i_44 (.A(in_b[15]), .ZN(n_22));
   INV_X1 i_45 (.A(in_b[19]), .ZN(n_23));
endmodule

module datapath__0_10(plus, p_0);
   output [63:0]plus;
   input [63:0]p_0;

   XOR2_X1 i_0 (.A(p_0[1]), .B(p_0[0]), .Z(plus[1]));
   AND2_X1 i_1 (.A1(n_13), .A2(n_0), .ZN(plus[2]));
   OAI21_X1 i_2 (.A(p_0[2]), .B1(p_0[1]), .B2(p_0[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(p_0[3]), .B(n_13), .Z(plus[3]));
   XOR2_X1 i_4 (.A(p_0[4]), .B(n_12), .Z(plus[4]));
   XOR2_X1 i_5 (.A(p_0[5]), .B(n_11), .Z(plus[5]));
   AND2_X1 i_6 (.A1(n_10), .A2(n_1), .ZN(plus[6]));
   OAI21_X1 i_7 (.A(p_0[6]), .B1(n_11), .B2(p_0[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(p_0[7]), .B(n_10), .Z(plus[7]));
   XOR2_X1 i_9 (.A(p_0[8]), .B(n_9), .Z(plus[8]));
   AND2_X1 i_10 (.A1(n_8), .A2(n_2), .ZN(plus[9]));
   OAI21_X1 i_11 (.A(p_0[9]), .B1(n_9), .B2(p_0[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(p_0[10]), .B(n_8), .Z(plus[10]));
   XOR2_X1 i_13 (.A(p_0[11]), .B(n_7), .Z(plus[11]));
   XOR2_X1 i_14 (.A(p_0[12]), .B(n_6), .Z(plus[12]));
   XNOR2_X1 i_15 (.A(p_0[13]), .B(n_5), .ZN(plus[13]));
   XOR2_X1 i_16 (.A(p_0[14]), .B(n_4), .Z(plus[14]));
   AND2_X1 i_17 (.A1(plus[63]), .A2(n_3), .ZN(plus[15]));
   OAI21_X1 i_18 (.A(p_0[15]), .B1(n_4), .B2(p_0[14]), .ZN(n_3));
   OR3_X1 i_19 (.A1(n_4), .A2(p_0[14]), .A3(p_0[15]), .ZN(plus[63]));
   NAND2_X1 i_20 (.A1(n_5), .A2(n_14), .ZN(n_4));
   NOR2_X1 i_21 (.A1(n_6), .A2(p_0[12]), .ZN(n_5));
   OR2_X1 i_22 (.A1(n_7), .A2(p_0[11]), .ZN(n_6));
   OR2_X1 i_23 (.A1(n_8), .A2(p_0[10]), .ZN(n_7));
   OR3_X1 i_24 (.A1(n_9), .A2(p_0[8]), .A3(p_0[9]), .ZN(n_8));
   OR2_X1 i_25 (.A1(n_10), .A2(p_0[7]), .ZN(n_9));
   OR3_X1 i_26 (.A1(n_11), .A2(p_0[5]), .A3(p_0[6]), .ZN(n_10));
   OR2_X1 i_27 (.A1(n_12), .A2(p_0[4]), .ZN(n_11));
   OR2_X1 i_28 (.A1(n_13), .A2(p_0[3]), .ZN(n_12));
   OR3_X1 i_29 (.A1(p_0[2]), .A2(p_0[1]), .A3(p_0[0]), .ZN(n_13));
   INV_X1 i_30 (.A(p_0[13]), .ZN(n_14));
endmodule

module fpu_divider(mode, clk, rst, enbl, in_a, in_b, out_c, done, err, zero, 
      posv);
   input [1:0]mode;
   input clk;
   input rst;
   input enbl;
   input [63:0]in_a;
   input [63:0]in_b;
   output [63:0]out_c;
   output done;
   output err;
   output zero;
   output posv;

   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire ovfl_flag;
   wire divide_by_zero_error;
   wire n_0_39;
   wire n_0_0;
   wire n_0_2_57;
   wire n_0_2_58;
   wire n_0_2_59;
   wire n_0_2_60;
   wire n_0_2_61;
   wire n_0_2_62;
   wire n_0_2_63;
   wire n_0_2_64;
   wire n_0_2_65;
   wire n_0_2_66;
   wire n_0_2_67;
   wire n_0_2_68;
   wire n_0_2_69;
   wire n_0_2_70;
   wire n_0_2_71;
   wire n_0_2_72;
   wire n_0_2_73;
   wire n_0_2_74;
   wire n_0_2_75;
   wire n_0_2_76;
   wire n_0_2_77;
   wire n_0_2_78;
   wire n_0_2_79;
   wire n_0_2_80;
   wire n_0_2_81;
   wire n_0_2_82;
   wire n_0_2_83;
   wire n_0_2_84;
   wire n_0_2_85;
   wire n_0_2_86;
   wire n_0_2_87;
   wire n_0_2_88;
   wire n_0_2_89;
   wire n_0_2_90;
   wire n_0_2_91;
   wire n_0_2_92;
   wire n_0_2_93;
   wire n_0_2_94;
   wire n_0_2_95;
   wire n_0_2_97;
   wire n_0_2_98;
   wire n_0_2_99;
   wire n_0_2_100;
   wire n_0_2_101;
   wire n_0_2_102;
   wire n_0_2_103;
   wire n_0_2_104;
   wire n_0_2_105;
   wire n_0_2_106;
   wire n_0_2_107;
   wire n_0_2_108;
   wire n_0_2_109;
   wire n_0_2_110;
   wire n_0_2_111;
   wire n_0_2_112;
   wire n_0_2_113;
   wire n_0_2_114;
   wire n_0_2_115;
   wire n_0_2_116;
   wire n_0_2_117;
   wire n_0_2_118;
   wire n_0_2_119;
   wire n_0_2_120;
   wire n_0_2_121;
   wire n_0_2_122;
   wire n_0_2_123;
   wire n_0_2_124;
   wire n_0_2_125;
   wire n_0_2_126;
   wire n_0_2_127;
   wire n_0_2_128;
   wire n_0_2_129;
   wire n_0_2_130;
   wire n_0_2_131;
   wire n_0_2_132;
   wire n_0_2_133;
   wire n_0_2_134;
   wire n_0_2_135;
   wire n_0_2_136;
   wire n_0_2_137;
   wire n_0_2_138;
   wire n_0_2_139;
   wire n_0_2_140;
   wire n_0_2_141;
   wire n_0_2_142;
   wire n_0_2_143;
   wire n_0_2_144;
   wire n_0_2_145;
   wire n_0_2_146;
   wire n_0_2_148;
   wire n_0_2_149;
   wire n_0_2_150;
   wire n_0_2_151;
   wire n_0_2_152;
   wire n_0_2_153;
   wire n_0_2_155;
   wire n_0_2_156;
   wire n_0_2_157;
   wire n_0_2_158;
   wire n_0_2_159;
   wire n_0_2_160;
   wire n_0_2_161;
   wire n_0_2_162;
   wire n_0_2_163;
   wire n_0_2_164;
   wire n_0_2_165;
   wire n_0_2_166;
   wire n_0_2_167;
   wire n_0_2_168;
   wire n_0_2_169;
   wire n_0_2_170;
   wire n_0_2_171;
   wire n_0_2_172;
   wire n_0_2_173;
   wire n_0_2_174;
   wire n_0_2_175;
   wire n_0_2_176;
   wire n_0_2_177;
   wire n_0_2_178;
   wire n_0_2_179;
   wire n_0_2_180;
   wire n_0_2_181;
   wire n_0_2_182;
   wire n_0_2_183;
   wire n_0_2_184;
   wire n_0_2_185;
   wire n_0_2_186;
   wire n_0_2_187;
   wire n_0_2_188;
   wire n_0_2_189;
   wire n_0_2_190;
   wire n_0_2_191;
   wire n_0_2_192;
   wire n_0_2_193;
   wire n_0_2_194;
   wire n_0_2_195;
   wire n_0_2_196;
   wire n_0_2_197;
   wire n_0_2_198;
   wire n_0_2_199;
   wire n_0_2_200;
   wire n_0_2_201;
   wire n_0_2_202;
   wire n_0_2_203;
   wire n_0_2_204;
   wire n_0_2_205;
   wire n_0_2_206;
   wire n_0_2_207;
   wire n_0_2_208;
   wire n_0_2_210;
   wire n_0_2_211;
   wire n_0_2_212;
   wire n_0_2_213;
   wire n_0_2_214;
   wire n_0_2_215;
   wire n_0_2_216;
   wire n_0_2_217;
   wire n_0_2_218;
   wire n_0_2_219;
   wire n_0_2_220;
   wire n_0_2_221;
   wire n_0_2_1522;
   wire n_0_2_222;
   wire n_0_2_223;
   wire n_0_2_224;
   wire n_0_2_225;
   wire n_0_2_226;
   wire n_0_2_1525;
   wire n_0_2_227;
   wire n_0_2_228;
   wire n_0_2_229;
   wire n_0_2_1579;
   wire n_0_2_1573;
   wire n_0_2_230;
   wire n_0_2_231;
   wire n_0_2_1570;
   wire n_0_2_0;
   wire n_0_2_1;
   wire n_0_2_232;
   wire n_0_2_233;
   wire n_0_2_1567;
   wire n_0_2_2;
   wire n_0_2_3;
   wire n_0_2_234;
   wire n_0_2_235;
   wire n_0_2_236;
   wire n_0_2_1564;
   wire n_0_2_4;
   wire n_0_2_5;
   wire n_0_2_237;
   wire n_0_2_238;
   wire n_0_2_239;
   wire n_0_2_1561;
   wire n_0_2_6;
   wire n_0_2_7;
   wire n_0_2_240;
   wire n_0_2_241;
   wire n_0_2_1558;
   wire n_0_2_8;
   wire n_0_2_9;
   wire n_0_2_242;
   wire n_0_2_243;
   wire n_0_2_244;
   wire n_0_2_1555;
   wire n_0_2_10;
   wire n_0_2_11;
   wire n_0_2_245;
   wire n_0_2_246;
   wire n_0_2_247;
   wire n_0_2_1552;
   wire n_0_2_12;
   wire n_0_2_13;
   wire n_0_2_248;
   wire n_0_2_249;
   wire n_0_2_1549;
   wire n_0_2_14;
   wire n_0_2_15;
   wire n_0_2_250;
   wire n_0_2_251;
   wire n_0_2_252;
   wire n_0_2_1546;
   wire n_0_2_16;
   wire n_0_2_17;
   wire n_0_2_253;
   wire n_0_2_254;
   wire n_0_2_1543;
   wire n_0_2_18;
   wire n_0_2_19;
   wire n_0_2_255;
   wire n_0_2_256;
   wire n_0_2_257;
   wire n_0_2_1540;
   wire n_0_2_20;
   wire n_0_2_21;
   wire n_0_2_258;
   wire n_0_2_259;
   wire n_0_2_260;
   wire n_0_2_1537;
   wire n_0_2_22;
   wire n_0_2_23;
   wire n_0_2_261;
   wire n_0_2_262;
   wire n_0_2_263;
   wire n_0_2_1534;
   wire n_0_2_1602;
   wire n_0_2_1598;
   wire n_0_2_264;
   wire n_0_2_265;
   wire n_0_2_266;
   wire n_0_2_1531;
   wire n_0_2_1595;
   wire n_0_2_1591;
   wire n_0_2_267;
   wire n_0_2_268;
   wire n_0_2_1590;
   wire n_0_2_269;
   wire n_0_2_270;
   wire n_0_2_271;
   wire n_0_2_1528;
   wire n_0_2_1588;
   wire n_0_2_1589;
   wire n_0_2_272;
   wire n_0_2_1585;
   wire n_0_2_273;
   wire [22:0]quotient;
   wire n_0_49;
   wire n_0_2_274;
   wire n_0_48;
   wire n_0_2_275;
   wire n_0_2_276;
   wire n_0_41;
   wire n_0_40;
   wire n_0_2_277;
   wire n_0_47;
   wire n_0_2_278;
   wire n_0_2_279;
   wire n_0_2_280;
   wire n_0_2_282;
   wire n_0_2_283;
   wire n_0_2_284;
   wire n_0_2_285;
   wire n_0_2_286;
   wire n_0_2_288;
   wire n_0_2_289;
   wire n_0_2_290;
   wire n_0_2_291;
   wire n_0_2_292;
   wire n_0_2_293;
   wire n_0_2_294;
   wire n_0_2_295;
   wire n_0_2_296;
   wire n_0_2_297;
   wire n_0_2_298;
   wire n_0_2_299;
   wire n_0_2_300;
   wire n_0_2_301;
   wire n_0_2_302;
   wire n_0_2_303;
   wire n_0_2_304;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_2_305;
   wire n_0_2_306;
   wire n_0_2_24;
   wire n_0_2_307;
   wire n_0_2_308;
   wire n_0_2_309;
   wire n_0_2_310;
   wire n_0_2_311;
   wire n_0_2_312;
   wire n_0_2_313;
   wire n_0_2_314;
   wire n_0_2_315;
   wire n_0_2_316;
   wire n_0_2_317;
   wire n_0_2_318;
   wire n_0_2_319;
   wire n_0_2_320;
   wire n_0_2_321;
   wire n_0_2_322;
   wire n_0_2_323;
   wire n_0_2_324;
   wire n_0_2_325;
   wire n_0_2_326;
   wire n_0_2_25;
   wire n_0_2_327;
   wire n_0_2_26;
   wire n_0_2_328;
   wire n_0_2_329;
   wire n_0_2_330;
   wire n_0_2_27;
   wire n_0_2_331;
   wire n_0_2_332;
   wire n_0_2_28;
   wire n_0_2_333;
   wire n_0_2_334;
   wire n_0_2_335;
   wire n_0_2_29;
   wire n_0_2_336;
   wire n_0_2_337;
   wire n_0_2_30;
   wire n_0_2_338;
   wire n_0_2_339;
   wire n_0_2_340;
   wire n_0_2_31;
   wire n_0_2_341;
   wire n_0_2_342;
   wire n_0_2_32;
   wire n_0_2_343;
   wire n_0_2_344;
   wire n_0_2_345;
   wire n_0_2_33;
   wire n_0_2_346;
   wire n_0_2_347;
   wire n_0_2_34;
   wire n_0_2_348;
   wire n_0_2_349;
   wire n_0_2_350;
   wire n_0_2_35;
   wire n_0_2_351;
   wire n_0_2_352;
   wire n_0_2_36;
   wire n_0_2_353;
   wire n_0_2_354;
   wire n_0_2_355;
   wire n_0_2_37;
   wire n_0_2_356;
   wire n_0_2_357;
   wire n_0_2_38;
   wire n_0_2_358;
   wire n_0_2_359;
   wire n_0_2_360;
   wire n_0_2_39;
   wire n_0_2_361;
   wire n_0_2_362;
   wire n_0_2_40;
   wire n_0_2_364;
   wire n_0_2_365;
   wire n_0_2_366;
   wire n_0_2_41;
   wire n_0_2_367;
   wire n_0_2_368;
   wire n_0_2_42;
   wire n_0_2_369;
   wire n_0_2_370;
   wire n_0_2_371;
   wire n_0_2_43;
   wire n_0_2_372;
   wire n_0_2_373;
   wire n_0_2_44;
   wire n_0_2_374;
   wire n_0_2_375;
   wire n_0_2_376;
   wire n_0_2_377;
   wire n_0_2_378;
   wire n_0_2_379;
   wire n_0_2_380;
   wire n_0_2_381;
   wire n_0_2_382;
   wire n_0_2_383;
   wire n_0_2_384;
   wire n_0_2_385;
   wire n_0_2_386;
   wire n_0_2_387;
   wire n_0_2_388;
   wire n_0_2_389;
   wire n_0_2_390;
   wire n_0_2_391;
   wire n_0_2_392;
   wire n_0_2_393;
   wire n_0_2_394;
   wire n_0_2_395;
   wire n_0_2_396;
   wire n_0_2_397;
   wire n_0_2_398;
   wire n_0_2_399;
   wire n_0_2_400;
   wire n_0_2_401;
   wire n_0_2_402;
   wire n_0_2_403;
   wire n_0_2_404;
   wire n_0_2_405;
   wire n_0_2_406;
   wire n_0_2_407;
   wire n_0_2_408;
   wire n_0_2_409;
   wire n_0_2_410;
   wire n_0_2_411;
   wire n_0_2_412;
   wire n_0_2_413;
   wire n_0_2_414;
   wire n_0_2_415;
   wire n_0_2_416;
   wire n_0_2_417;
   wire n_0_2_418;
   wire n_0_2_419;
   wire n_0_2_420;
   wire n_0_2_421;
   wire n_0_2_422;
   wire n_0_2_423;
   wire n_0_2_424;
   wire n_0_2_425;
   wire n_0_2_426;
   wire n_0_2_427;
   wire n_0_2_428;
   wire n_0_2_429;
   wire n_0_2_430;
   wire n_0_2_431;
   wire n_0_2_432;
   wire n_0_2_433;
   wire n_0_2_434;
   wire n_0_2_435;
   wire n_0_2_436;
   wire n_0_2_437;
   wire n_0_2_438;
   wire n_0_2_439;
   wire n_0_2_440;
   wire n_0_2_441;
   wire n_0_2_442;
   wire n_0_2_443;
   wire n_0_2_444;
   wire n_0_2_445;
   wire n_0_2_446;
   wire n_0_2_447;
   wire n_0_2_448;
   wire n_0_2_449;
   wire n_0_2_450;
   wire n_0_2_451;
   wire n_0_2_452;
   wire n_0_2_454;
   wire n_0_2_455;
   wire n_0_2_456;
   wire n_0_2_457;
   wire n_0_2_459;
   wire n_0_2_460;
   wire n_0_2_461;
   wire n_0_2_462;
   wire n_0_2_463;
   wire n_0_2_464;
   wire n_0_2_465;
   wire n_0_2_466;
   wire n_0_2_467;
   wire n_0_2_468;
   wire n_0_2_469;
   wire n_0_2_470;
   wire n_0_2_471;
   wire n_0_2_472;
   wire n_0_2_473;
   wire n_0_2_474;
   wire n_0_2_475;
   wire n_0_2_476;
   wire n_0_2_477;
   wire n_0_2_478;
   wire n_0_2_479;
   wire n_0_2_480;
   wire n_0_2_481;
   wire n_0_2_482;
   wire n_0_2_483;
   wire n_0_2_484;
   wire n_0_2_485;
   wire n_0_2_486;
   wire n_0_2_487;
   wire n_0_2_488;
   wire n_0_2_489;
   wire n_0_2_490;
   wire n_0_2_491;
   wire n_0_2_492;
   wire n_0_2_493;
   wire n_0_2_494;
   wire n_0_2_495;
   wire n_0_2_496;
   wire n_0_2_497;
   wire n_0_2_498;
   wire n_0_2_499;
   wire n_0_2_500;
   wire n_0_2_501;
   wire n_0_2_502;
   wire n_0_2_503;
   wire n_0_2_504;
   wire n_0_2_505;
   wire n_0_2_506;
   wire n_0_2_507;
   wire n_0_2_508;
   wire n_0_2_509;
   wire n_0_2_510;
   wire n_0_2_511;
   wire n_0_2_512;
   wire n_0_2_513;
   wire n_0_2_514;
   wire n_0_2_515;
   wire n_0_2_516;
   wire n_0_2_517;
   wire n_0_2_518;
   wire n_0_2_519;
   wire n_0_2_520;
   wire n_0_2_521;
   wire n_0_2_522;
   wire n_0_2_523;
   wire n_0_2_524;
   wire n_0_2_525;
   wire n_0_2_526;
   wire n_0_2_527;
   wire n_0_2_528;
   wire n_0_2_529;
   wire n_0_2_530;
   wire n_0_2_531;
   wire n_0_2_532;
   wire n_0_2_533;
   wire n_0_2_534;
   wire n_0_2_535;
   wire n_0_2_536;
   wire n_0_2_537;
   wire n_0_2_538;
   wire n_0_2_539;
   wire n_0_2_540;
   wire n_0_2_541;
   wire n_0_2_542;
   wire n_0_2_543;
   wire n_0_2_544;
   wire n_0_2_545;
   wire n_0_2_546;
   wire n_0_2_547;
   wire n_0_2_548;
   wire n_0_2_549;
   wire n_0_2_550;
   wire n_0_2_551;
   wire n_0_2_552;
   wire n_0_2_553;
   wire n_0_2_554;
   wire n_0_2_555;
   wire n_0_2_556;
   wire n_0_2_557;
   wire n_0_2_558;
   wire n_0_2_559;
   wire n_0_2_560;
   wire n_0_2_561;
   wire n_0_2_562;
   wire n_0_2_563;
   wire n_0_2_564;
   wire n_0_2_565;
   wire n_0_2_566;
   wire n_0_2_567;
   wire n_0_2_568;
   wire n_0_2_569;
   wire n_0_2_570;
   wire n_0_2_571;
   wire n_0_2_572;
   wire n_0_2_573;
   wire n_0_2_574;
   wire n_0_2_575;
   wire n_0_2_576;
   wire n_0_2_577;
   wire n_0_2_578;
   wire n_0_2_579;
   wire n_0_2_580;
   wire n_0_2_581;
   wire n_0_2_582;
   wire n_0_2_583;
   wire n_0_2_584;
   wire n_0_2_585;
   wire n_0_2_586;
   wire n_0_2_587;
   wire n_0_2_588;
   wire n_0_2_589;
   wire n_0_2_590;
   wire n_0_2_591;
   wire n_0_2_592;
   wire n_0_2_593;
   wire n_0_2_594;
   wire n_0_2_595;
   wire n_0_2_596;
   wire n_0_2_597;
   wire n_0_2_598;
   wire n_0_2_599;
   wire n_0_2_600;
   wire n_0_2_601;
   wire n_0_2_602;
   wire n_0_2_603;
   wire n_0_2_604;
   wire n_0_2_605;
   wire n_0_2_606;
   wire n_0_2_607;
   wire n_0_2_608;
   wire n_0_2_609;
   wire n_0_2_610;
   wire n_0_2_611;
   wire n_0_2_612;
   wire n_0_2_613;
   wire n_0_2_614;
   wire n_0_2_615;
   wire n_0_2_616;
   wire n_0_2_617;
   wire n_0_2_618;
   wire n_0_2_619;
   wire n_0_2_620;
   wire n_0_2_621;
   wire n_0_2_622;
   wire n_0_2_623;
   wire n_0_2_624;
   wire n_0_2_625;
   wire n_0_2_626;
   wire n_0_2_627;
   wire n_0_2_628;
   wire n_0_2_629;
   wire n_0_2_630;
   wire n_0_2_631;
   wire n_0_2_632;
   wire n_0_2_633;
   wire n_0_2_634;
   wire n_0_2_635;
   wire n_0_2_636;
   wire n_0_2_637;
   wire n_0_2_638;
   wire n_0_2_639;
   wire n_0_2_640;
   wire n_0_2_641;
   wire n_0_2_642;
   wire n_0_2_643;
   wire n_0_2_644;
   wire n_0_2_645;
   wire n_0_2_646;
   wire n_0_2_647;
   wire n_0_2_648;
   wire n_0_2_649;
   wire n_0_2_650;
   wire n_0_2_651;
   wire n_0_2_652;
   wire n_0_2_653;
   wire n_0_2_654;
   wire n_0_2_655;
   wire n_0_2_656;
   wire n_0_2_657;
   wire n_0_2_658;
   wire n_0_2_659;
   wire n_0_2_661;
   wire n_0_2_662;
   wire n_0_2_663;
   wire n_0_2_664;
   wire n_0_2_665;
   wire n_0_2_666;
   wire n_0_2_668;
   wire n_0_2_669;
   wire n_0_2_670;
   wire n_0_2_671;
   wire n_0_2_672;
   wire n_0_2_673;
   wire n_0_2_674;
   wire n_0_2_675;
   wire n_0_2_676;
   wire n_0_2_677;
   wire n_0_2_678;
   wire n_0_2_679;
   wire n_0_2_680;
   wire n_0_2_681;
   wire n_0_2_682;
   wire n_0_2_683;
   wire n_0_2_684;
   wire n_0_2_685;
   wire n_0_2_686;
   wire n_0_2_687;
   wire n_0_2_688;
   wire n_0_2_689;
   wire n_0_2_690;
   wire n_0_2_691;
   wire n_0_2_692;
   wire n_0_2_693;
   wire n_0_2_694;
   wire n_0_2_695;
   wire n_0_2_696;
   wire n_0_2_697;
   wire n_0_2_698;
   wire n_0_2_699;
   wire n_0_2_700;
   wire n_0_2_701;
   wire n_0_2_702;
   wire n_0_2_703;
   wire n_0_2_704;
   wire n_0_2_705;
   wire n_0_2_706;
   wire n_0_2_707;
   wire n_0_2_708;
   wire n_0_2_709;
   wire n_0_2_710;
   wire n_0_2_711;
   wire n_0_2_712;
   wire n_0_2_713;
   wire n_0_2_714;
   wire n_0_2_715;
   wire n_0_2_716;
   wire n_0_2_717;
   wire n_0_2_718;
   wire n_0_2_719;
   wire n_0_2_720;
   wire n_0_2_721;
   wire n_0_2_722;
   wire n_0_2_723;
   wire n_0_2_724;
   wire n_0_2_725;
   wire n_0_2_726;
   wire n_0_2_727;
   wire n_0_2_728;
   wire n_0_2_729;
   wire n_0_2_730;
   wire n_0_2_731;
   wire n_0_2_732;
   wire n_0_2_733;
   wire n_0_2_734;
   wire n_0_2_735;
   wire n_0_2_736;
   wire n_0_2_737;
   wire n_0_2_738;
   wire n_0_2_739;
   wire n_0_2_740;
   wire n_0_2_741;
   wire n_0_2_742;
   wire n_0_2_743;
   wire n_0_2_45;
   wire n_0_2_46;
   wire n_0_2_47;
   wire n_0_2_744;
   wire n_0_2_745;
   wire n_0_2_746;
   wire n_0_2_48;
   wire n_0_2_747;
   wire n_0_2_748;
   wire n_0_2_749;
   wire n_0_2_1246;
   wire n_0_2_750;
   wire n_0_2_751;
   wire n_0_2_752;
   wire n_0_2_753;
   wire n_0_2_754;
   wire n_0_2_755;
   wire n_0_2_756;
   wire n_0_2_757;
   wire n_0_2_758;
   wire n_0_2_759;
   wire n_0_2_760;
   wire n_0_2_761;
   wire n_0_2_762;
   wire n_0_2_763;
   wire n_0_2_764;
   wire n_0_2_765;
   wire n_0_2_766;
   wire n_0_2_1255;
   wire n_0_2_767;
   wire n_0_2_1247;
   wire n_0_2_1091;
   wire n_0_2_768;
   wire n_0_2_287;
   wire n_0_2_1196;
   wire n_0_2_769;
   wire n_0_2_770;
   wire n_0_2_771;
   wire n_0_2_772;
   wire n_0_2_773;
   wire n_0_2_774;
   wire n_0_2_775;
   wire n_0_2_776;
   wire n_0_2_777;
   wire n_0_2_778;
   wire n_0_2_779;
   wire n_0_2_781;
   wire n_0_2_782;
   wire n_0_2_783;
   wire n_0_2_784;
   wire n_0_2_785;
   wire n_0_2_786;
   wire n_0_2_787;
   wire n_0_2_788;
   wire n_0_2_789;
   wire n_0_2_790;
   wire n_0_2_791;
   wire n_0_2_792;
   wire n_0_2_793;
   wire n_0_2_794;
   wire n_0_2_795;
   wire n_0_2_796;
   wire n_0_2_797;
   wire n_0_2_798;
   wire n_0_2_799;
   wire n_0_2_800;
   wire n_0_2_801;
   wire n_0_2_802;
   wire n_0_2_803;
   wire n_0_2_804;
   wire n_0_2_805;
   wire n_0_2_806;
   wire n_0_2_807;
   wire n_0_2_808;
   wire n_0_2_809;
   wire n_0_2_810;
   wire n_0_2_811;
   wire n_0_2_812;
   wire n_0_2_813;
   wire n_0_2_814;
   wire n_0_2_815;
   wire n_0_2_816;
   wire n_0_2_817;
   wire n_0_2_818;
   wire n_0_2_819;
   wire n_0_2_820;
   wire n_0_2_821;
   wire n_0_2_822;
   wire n_0_2_823;
   wire n_0_2_824;
   wire n_0_2_825;
   wire n_0_2_826;
   wire n_0_2_827;
   wire n_0_2_828;
   wire n_0_2_829;
   wire n_0_2_830;
   wire n_0_2_831;
   wire n_0_2_832;
   wire n_0_2_833;
   wire n_0_2_834;
   wire n_0_2_835;
   wire n_0_2_836;
   wire n_0_2_837;
   wire n_0_2_838;
   wire n_0_50;
   wire n_0_2_839;
   wire n_0_51;
   wire n_0_2_840;
   wire n_0_52;
   wire n_0_2_841;
   wire n_0_53;
   wire n_0_2_842;
   wire n_0_54;
   wire n_0_2_843;
   wire n_0_55;
   wire n_0_2_844;
   wire n_0_56;
   wire n_0_2_845;
   wire n_0_57;
   wire n_0_2_846;
   wire n_0_2_847;
   wire n_0_58;
   wire n_0_2_848;
   wire n_0_2_849;
   wire n_0_2_850;
   wire n_0_2_851;
   wire n_0_2_852;
   wire n_0_2_853;
   wire n_0_2_854;
   wire n_0_2_855;
   wire n_0_2_856;
   wire n_0_2_857;
   wire n_0_2_858;
   wire n_0_2_859;
   wire n_0_2_860;
   wire n_0_2_861;
   wire n_0_2_862;
   wire n_0_2_863;
   wire n_0_2_864;
   wire n_0_2_865;
   wire n_0_2_866;
   wire n_0_2_867;
   wire n_0_2_868;
   wire n_0_2_869;
   wire n_0_2_870;
   wire n_0_2_871;
   wire n_0_59;
   wire n_0_2_872;
   wire n_0_2_873;
   wire n_0_2_874;
   wire n_0_2_875;
   wire n_0_2_876;
   wire n_0_2_877;
   wire n_0_2_878;
   wire n_0_2_879;
   wire n_0_2_880;
   wire n_0_2_881;
   wire n_0_2_882;
   wire n_0_2_883;
   wire n_0_2_884;
   wire n_0_2_885;
   wire n_0_2_886;
   wire n_0_2_887;
   wire n_0_2_888;
   wire n_0_2_889;
   wire n_0_2_890;
   wire n_0_2_891;
   wire n_0_2_892;
   wire n_0_2_893;
   wire n_0_2_894;
   wire n_0_2_895;
   wire n_0_2_896;
   wire n_0_2_897;
   wire n_0_2_898;
   wire n_0_2_899;
   wire n_0_2_900;
   wire n_0_2_901;
   wire n_0_2_902;
   wire n_0_2_903;
   wire n_0_2_904;
   wire n_0_2_905;
   wire n_0_2_906;
   wire n_0_2_908;
   wire n_0_2_909;
   wire n_0_2_910;
   wire n_0_2_911;
   wire n_0_2_912;
   wire n_0_2_913;
   wire n_0_2_914;
   wire n_0_2_915;
   wire n_0_2_916;
   wire n_0_2_917;
   wire n_0_2_918;
   wire n_0_2_919;
   wire n_0_2_920;
   wire n_0_2_921;
   wire n_0_2_922;
   wire n_0_2_923;
   wire n_0_2_924;
   wire n_0_2_925;
   wire n_0_2_926;
   wire n_0_2_927;
   wire n_0_2_928;
   wire n_0_2_929;
   wire n_0_2_930;
   wire n_0_2_931;
   wire n_0_2_932;
   wire n_0_2_933;
   wire n_0_2_934;
   wire n_0_2_935;
   wire n_0_2_936;
   wire n_0_2_937;
   wire n_0_2_938;
   wire n_0_2_939;
   wire n_0_2_940;
   wire n_0_2_941;
   wire n_0_2_942;
   wire n_0_2_943;
   wire n_0_2_944;
   wire n_0_2_945;
   wire n_0_2_946;
   wire n_0_2_947;
   wire n_0_2_948;
   wire n_0_2_949;
   wire n_0_2_950;
   wire n_0_2_951;
   wire n_0_2_952;
   wire n_0_2_953;
   wire n_0_2_954;
   wire n_0_2_955;
   wire n_0_2_956;
   wire n_0_2_957;
   wire n_0_2_958;
   wire n_0_2_959;
   wire n_0_2_960;
   wire n_0_2_961;
   wire n_0_2_962;
   wire n_0_2_963;
   wire n_0_2_964;
   wire n_0_2_965;
   wire n_0_2_966;
   wire n_0_2_967;
   wire n_0_2_968;
   wire n_0_2_969;
   wire n_0_2_970;
   wire n_0_2_971;
   wire n_0_2_972;
   wire n_0_2_973;
   wire n_0_2_974;
   wire n_0_2_975;
   wire n_0_2_976;
   wire n_0_2_977;
   wire n_0_2_978;
   wire n_0_2_979;
   wire n_0_2_980;
   wire n_0_2_981;
   wire n_0_2_982;
   wire n_0_2_983;
   wire n_0_2_984;
   wire n_0_2_985;
   wire n_0_2_986;
   wire n_0_2_987;
   wire n_0_2_988;
   wire n_0_2_989;
   wire n_0_2_990;
   wire n_0_2_991;
   wire n_0_2_992;
   wire n_0_2_993;
   wire n_0_2_994;
   wire n_0_2_995;
   wire n_0_2_996;
   wire n_0_2_997;
   wire n_0_2_998;
   wire n_0_2_999;
   wire n_0_2_1000;
   wire n_0_2_1001;
   wire n_0_2_1002;
   wire n_0_2_1003;
   wire n_0_2_1004;
   wire n_0_2_1005;
   wire n_0_2_1006;
   wire n_0_2_1007;
   wire n_0_2_1008;
   wire n_0_2_1009;
   wire n_0_2_1010;
   wire n_0_2_1011;
   wire n_0_2_1012;
   wire n_0_2_1013;
   wire n_0_2_1014;
   wire n_0_2_1015;
   wire n_0_2_1016;
   wire n_0_2_1017;
   wire n_0_2_1018;
   wire n_0_2_1019;
   wire n_0_2_1020;
   wire n_0_2_1021;
   wire n_0_2_1022;
   wire n_0_2_1023;
   wire n_0_2_1024;
   wire n_0_2_1025;
   wire n_0_2_1026;
   wire n_0_2_1027;
   wire n_0_2_1028;
   wire n_0_2_1029;
   wire n_0_2_1030;
   wire n_0_2_1031;
   wire n_0_2_1032;
   wire n_0_2_1033;
   wire n_0_2_1034;
   wire n_0_2_1035;
   wire n_0_2_1036;
   wire n_0_2_1037;
   wire n_0_2_1038;
   wire n_0_2_1039;
   wire n_0_2_1040;
   wire n_0_2_1041;
   wire n_0_2_1042;
   wire n_0_2_1043;
   wire n_0_2_1045;
   wire n_0_2_1046;
   wire n_0_2_1047;
   wire n_0_2_1048;
   wire n_0_2_1049;
   wire n_0_2_1050;
   wire n_0_2_1051;
   wire n_0_2_1052;
   wire n_0_2_1053;
   wire n_0_2_1054;
   wire n_0_2_1055;
   wire n_0_2_1056;
   wire n_0_2_1057;
   wire n_0_2_1058;
   wire n_0_2_1059;
   wire n_0_2_1060;
   wire n_0_2_1061;
   wire n_0_2_1062;
   wire n_0_2_1063;
   wire n_0_2_1064;
   wire n_0_2_1065;
   wire n_0_2_1066;
   wire n_0_2_1067;
   wire n_0_2_1068;
   wire n_0_2_1069;
   wire n_0_2_1070;
   wire n_0_2_1071;
   wire n_0_2_1072;
   wire n_0_2_1073;
   wire n_0_2_1074;
   wire n_0_2_1075;
   wire n_0_2_1076;
   wire n_0_2_1077;
   wire n_0_2_1078;
   wire n_0_2_1079;
   wire n_0_2_1080;
   wire n_0_2_1081;
   wire n_0_2_1082;
   wire n_0_2_1083;
   wire n_0_2_1084;
   wire n_0_2_1085;
   wire n_0_2_1086;
   wire n_0_2_1087;
   wire n_0_2_1088;
   wire n_0_2_1089;
   wire n_0_2_1090;
   wire n_0_2_1092;
   wire n_0_2_1093;
   wire n_0_2_1094;
   wire n_0_2_1095;
   wire n_0_2_1096;
   wire n_0_2_1097;
   wire n_0_2_1098;
   wire n_0_2_1099;
   wire n_0_2_1100;
   wire n_0_2_1101;
   wire n_0_2_1102;
   wire n_0_2_1103;
   wire n_0_2_1104;
   wire n_0_2_1105;
   wire n_0_2_1106;
   wire n_0_2_1107;
   wire n_0_2_1108;
   wire n_0_2_1109;
   wire n_0_2_1110;
   wire n_0_2_1111;
   wire n_0_2_1112;
   wire n_0_2_1113;
   wire n_0_2_1114;
   wire n_0_2_1115;
   wire n_0_2_1116;
   wire n_0_2_1117;
   wire n_0_2_1118;
   wire n_0_2_1119;
   wire n_0_2_1120;
   wire n_0_2_1121;
   wire n_0_2_1122;
   wire n_0_2_1123;
   wire n_0_2_1124;
   wire n_0_2_1125;
   wire n_0_2_1126;
   wire n_0_2_1127;
   wire n_0_2_1128;
   wire n_0_2_1129;
   wire n_0_2_1130;
   wire n_0_2_1131;
   wire n_0_2_1132;
   wire n_0_2_1133;
   wire n_0_2_1134;
   wire n_0_2_1135;
   wire n_0_2_1136;
   wire n_0_2_1137;
   wire n_0_2_1138;
   wire n_0_2_1139;
   wire n_0_2_1140;
   wire n_0_2_1141;
   wire n_0_2_1142;
   wire n_0_2_1143;
   wire n_0_2_1144;
   wire n_0_2_1145;
   wire n_0_2_1146;
   wire n_0_2_1147;
   wire n_0_2_1148;
   wire n_0_2_1149;
   wire n_0_2_1150;
   wire n_0_2_1151;
   wire n_0_2_1152;
   wire n_0_2_1153;
   wire n_0_2_1154;
   wire n_0_2_1155;
   wire n_0_2_1156;
   wire n_0_2_1157;
   wire n_0_2_1158;
   wire n_0_2_1159;
   wire n_0_2_1160;
   wire n_0_2_1161;
   wire n_0_2_1162;
   wire n_0_2_1163;
   wire n_0_2_1164;
   wire n_0_2_1165;
   wire n_0_2_1166;
   wire n_0_2_1167;
   wire n_0_2_1168;
   wire n_0_2_1169;
   wire n_0_2_1170;
   wire n_0_2_1171;
   wire n_0_2_1172;
   wire n_0_2_1173;
   wire n_0_2_1174;
   wire n_0_2_1175;
   wire n_0_2_1176;
   wire n_0_2_1177;
   wire n_0_2_1178;
   wire n_0_2_1179;
   wire n_0_2_1180;
   wire n_0_2_1181;
   wire n_0_2_1182;
   wire n_0_2_1183;
   wire n_0_2_1184;
   wire n_0_2_1185;
   wire n_0_2_1186;
   wire n_0_2_1187;
   wire n_0_2_1188;
   wire n_0_2_1189;
   wire n_0_2_1191;
   wire n_0_2_1192;
   wire n_0_2_1193;
   wire n_0_2_1194;
   wire n_0_2_1195;
   wire n_0_2_1198;
   wire n_0_2_1199;
   wire n_0_2_1200;
   wire n_0_2_1201;
   wire n_0_2_1202;
   wire n_0_2_1203;
   wire n_0_2_1204;
   wire n_0_2_1205;
   wire n_0_2_1206;
   wire n_0_2_1207;
   wire n_0_2_1208;
   wire n_0_2_1209;
   wire n_0_2_1210;
   wire n_0_2_1211;
   wire n_0_2_1212;
   wire n_0_2_1213;
   wire n_0_2_1214;
   wire n_0_2_1215;
   wire n_0_2_1216;
   wire n_0_2_1217;
   wire n_0_2_1218;
   wire n_0_2_1219;
   wire n_0_2_1220;
   wire n_0_2_1221;
   wire n_0_2_1222;
   wire n_0_2_1223;
   wire n_0_2_1224;
   wire n_0_2_1225;
   wire n_0_2_1226;
   wire n_0_2_1227;
   wire n_0_2_1228;
   wire n_0_2_1229;
   wire n_0_2_1230;
   wire n_0_2_1231;
   wire n_0_2_1232;
   wire n_0_2_1233;
   wire n_0_2_1234;
   wire n_0_2_1235;
   wire n_0_2_1236;
   wire n_0_2_1237;
   wire n_0_2_1238;
   wire n_0_2_1239;
   wire n_0_2_1240;
   wire n_0_2_1241;
   wire n_0_2_1242;
   wire n_0_2_1243;
   wire n_0_2_1244;
   wire n_0_2_1245;
   wire n_0_2_1248;
   wire n_0_2_1249;
   wire n_0_2_1250;
   wire n_0_2_1251;
   wire n_0_2_1252;
   wire n_0_2_1253;
   wire n_0_2_1254;
   wire n_0_2_1256;
   wire n_0_2_1257;
   wire n_0_2_1258;
   wire n_0_2_1259;
   wire n_0_2_1260;
   wire n_0_2_1261;
   wire n_0_2_1262;
   wire n_0_2_1263;
   wire n_0_2_1264;
   wire n_0_2_1265;
   wire n_0_2_1266;
   wire n_0_2_1267;
   wire n_0_2_1268;
   wire n_0_2_1269;
   wire n_0_2_1270;
   wire n_0_2_1271;
   wire n_0_2_1272;
   wire n_0_2_1273;
   wire n_0_2_1274;
   wire n_0_2_1275;
   wire n_0_2_1276;
   wire n_0_2_1277;
   wire n_0_2_1278;
   wire n_0_2_1279;
   wire n_0_2_1280;
   wire n_0_2_1281;
   wire n_0_2_1282;
   wire n_0_2_1283;
   wire n_0_2_1284;
   wire n_0_2_1285;
   wire n_0_2_1286;
   wire n_0_2_1287;
   wire n_0_2_1288;
   wire n_0_2_1289;
   wire n_0_2_1290;
   wire n_0_2_1291;
   wire n_0_2_1292;
   wire n_0_2_1293;
   wire n_0_2_1294;
   wire n_0_2_1295;
   wire n_0_2_1296;
   wire n_0_2_1297;
   wire n_0_2_1298;
   wire n_0_2_1299;
   wire n_0_2_1300;
   wire n_0_2_1301;
   wire n_0_2_1302;
   wire n_0_2_1303;
   wire n_0_2_1304;
   wire n_0_2_1305;
   wire n_0_2_1306;
   wire n_0_2_1307;
   wire n_0_2_1308;
   wire n_0_2_1309;
   wire n_0_2_1310;
   wire n_0_2_1311;
   wire n_0_2_1312;
   wire n_0_2_1313;
   wire n_0_2_1314;
   wire n_0_2_1315;
   wire n_0_2_1316;
   wire n_0_2_1317;
   wire n_0_2_1318;
   wire n_0_2_1319;
   wire n_0_2_1320;
   wire n_0_2_1321;
   wire n_0_2_1322;
   wire n_0_2_1323;
   wire n_0_2_1324;
   wire n_0_2_1325;
   wire n_0_2_1326;
   wire n_0_2_1327;
   wire n_0_2_1328;
   wire n_0_2_1329;
   wire n_0_2_1330;
   wire n_0_2_1331;
   wire n_0_2_1332;
   wire n_0_2_1333;
   wire n_0_2_1334;
   wire n_0_2_1335;
   wire n_0_2_1336;
   wire n_0_2_1337;
   wire n_0_2_1338;
   wire n_0_2_1339;
   wire n_0_2_1340;
   wire n_0_2_1341;
   wire n_0_2_1342;
   wire n_0_2_1343;
   wire n_0_2_1344;
   wire n_0_2_1345;
   wire n_0_2_1346;
   wire n_0_2_1347;
   wire n_0_2_1348;
   wire n_0_2_1349;
   wire n_0_2_1350;
   wire n_0_2_1351;
   wire n_0_2_1353;
   wire n_0_2_1354;
   wire n_0_2_1355;
   wire n_0_2_1356;
   wire n_0_2_1357;
   wire n_0_2_1358;
   wire n_0_2_1359;
   wire n_0_2_1360;
   wire n_0_2_1361;
   wire n_0_2_1362;
   wire n_0_2_1363;
   wire n_0_2_1364;
   wire n_0_2_1365;
   wire n_0_2_1366;
   wire n_0_2_1367;
   wire n_0_2_1368;
   wire n_0_2_1369;
   wire n_0_2_1370;
   wire n_0_2_1371;
   wire n_0_2_1372;
   wire n_0_2_1373;
   wire n_0_2_1374;
   wire n_0_2_1375;
   wire n_0_2_1376;
   wire n_0_2_1377;
   wire n_0_2_1378;
   wire n_0_2_1379;
   wire n_0_2_1380;
   wire n_0_2_1381;
   wire n_0_2_1382;
   wire n_0_2_1383;
   wire n_0_2_1384;
   wire n_0_2_1385;
   wire n_0_2_1386;
   wire n_0_2_1387;
   wire n_0_2_1388;
   wire n_0_2_1389;
   wire n_0_2_1390;
   wire n_0_2_1391;
   wire n_0_2_1392;
   wire n_0_2_1393;
   wire n_0_2_1394;
   wire n_0_2_1395;
   wire n_0_2_1396;
   wire n_0_2_1397;
   wire n_0_2_1412;
   wire n_0_2_1398;
   wire n_0_2_49;
   wire n_0_2_1399;
   wire n_0_2_1400;
   wire n_0_2_54;
   wire n_0_2_1401;
   wire n_0_2_1402;
   wire n_0_2_1403;
   wire n_0_2_96;
   wire n_0_2_1404;
   wire n_0_2_1406;
   wire n_0_2_147;
   wire n_0_2_1407;
   wire n_0_2_1408;
   wire n_0_2_209;
   wire n_0_2_1409;
   wire n_0_2_1410;
   wire n_0_2_281;
   wire n_0_2_1411;
   wire n_0_2_1413;
   wire n_0_2_363;
   wire n_0_2_1414;
   wire n_0_2_1415;
   wire n_0_2_453;
   wire n_0_2_1416;
   wire n_0_2_1417;
   wire n_0_2_458;
   wire n_0_2_1418;
   wire n_0_2_660;
   wire n_0_2_1419;
   wire n_0_2_1420;
   wire n_0_2_1421;
   wire n_0_2_907;
   wire n_0_2_1422;
   wire n_0_2_1423;
   wire n_0_2_1424;
   wire n_0_2_1044;
   wire n_0_2_1425;
   wire n_0_2_1426;
   wire n_0_2_1427;
   wire n_0_2_1352;
   wire n_0_2_1428;
   wire n_0_2_1516;
   wire n_0_2_1429;
   wire n_0_2_1190;
   wire n_0_2_1430;
   wire n_0_2_1431;
   wire n_0_2_1432;
   wire n_0_2_667;
   wire n_0_2_1433;
   wire n_0_2_50;
   wire n_0_2_154;
   wire n_0_2_51;
   wire n_0_2_1434;
   wire n_0_2_52;
   wire n_0_2_1197;
   wire n_0_2_1435;
   wire n_0_2_1436;
   wire n_0_2_53;
   wire n_0_2_1437;
   wire n_0_2_1438;
   wire n_0_2_55;
   wire n_0_2_1439;
   wire n_0_2_56;
   wire n_0_2_1440;
   wire n_0_2_780;
   wire n_0_2_1441;
   wire n_0_2_1442;
   wire n_0_2_1443;
   wire n_0_2_1444;
   wire n_0_2_1445;
   wire n_0_2_1446;
   wire n_0_2_1447;
   wire n_0_2_1448;
   wire n_0_2_1449;
   wire n_0_2_1450;
   wire n_0_2_1451;
   wire n_0_2_1452;
   wire n_0_2_1405;
   wire n_0_2_1453;
   wire n_0_2_1454;
   wire n_0_2_1455;
   wire n_0_2_1456;
   wire n_0_2_1457;
   wire n_0_2_1458;
   wire n_0_2_1459;
   wire n_0_2_1460;
   wire n_0_2_1461;
   wire n_0_2_1462;
   wire n_0_2_1463;
   wire n_0_2_1464;
   wire n_0_2_1465;
   wire n_0_2_1466;
   wire n_0_2_1467;
   wire n_0_2_1468;
   wire n_0_2_1469;
   wire n_0_2_1470;
   wire n_0_2_1471;
   wire n_0_2_1472;
   wire n_0_2_1473;
   wire n_0_2_1474;
   wire n_0_2_1475;
   wire n_0_2_1476;
   wire n_0_2_1477;
   wire n_0_2_1478;
   wire n_0_2_1479;
   wire n_0_2_1480;
   wire n_0_2_1481;
   wire n_0_2_1482;
   wire n_0_2_1483;
   wire n_0_42;
   wire n_0_2_1484;
   wire n_0_2_1485;
   wire n_0_2_1486;
   wire n_0_2_1487;
   wire n_0_2_1488;
   wire n_0_2_1489;
   wire n_0_2_1490;
   wire n_0_2_1491;
   wire n_0_2_1492;
   wire n_0_2_1493;
   wire n_0_2_1494;
   wire n_0_2_1495;
   wire n_0_2_1496;
   wire n_0_2_1497;
   wire n_0_2_1498;
   wire n_0_2_1499;
   wire n_0_2_1500;
   wire n_0_2_1501;
   wire n_0_2_1502;
   wire n_0_2_1503;
   wire n_0_2_1504;
   wire n_0_2_1505;
   wire n_0_2_1506;
   wire n_0_2_1507;
   wire n_0_2_1508;
   wire n_0_2_1509;
   wire n_0_2_1510;
   wire n_0_2_1511;
   wire n_0_2_1512;
   wire n_0_2_1513;
   wire n_0_2_1514;
   wire n_0_2_1515;
   wire n_0_2_1517;
   wire n_0_2_1518;
   wire n_0_2_1519;
   wire n_0_2_1520;
   wire n_0_2_1521;
   wire n_0_2_1523;
   wire n_0_2_1524;
   wire n_0_2_1526;
   wire n_0_2_1527;
   wire n_0_2_1529;
   wire n_0_2_1530;
   wire n_0_2_1532;
   wire n_0_2_1533;
   wire n_0_2_1535;
   wire n_0_2_1536;
   wire n_0_2_1538;
   wire n_0_2_1539;
   wire n_0_2_1541;
   wire n_0_2_1542;
   wire n_0_2_1544;
   wire n_0_2_1545;
   wire n_0_2_1547;
   wire n_0_2_1548;
   wire n_0_2_1550;
   wire n_0_2_1551;
   wire n_0_2_1553;
   wire n_0_2_1554;
   wire n_0_2_1556;
   wire n_0_2_1557;
   wire n_0_2_1559;
   wire n_0_2_1560;
   wire n_0_2_1562;
   wire n_0_2_1563;
   wire n_0_2_1565;
   wire n_0_2_1566;
   wire n_0_2_1568;
   wire n_0_2_1569;
   wire n_0_2_1571;
   wire n_0_2_1572;
   wire n_0_2_1574;
   wire n_0_2_1575;
   wire n_0_2_1576;
   wire n_0_2_1577;
   wire n_0_2_1578;
   wire n_0_2_1580;
   wire n_0_2_1581;
   wire n_0_2_1582;
   wire n_0_2_1583;
   wire n_0_2_1584;
   wire n_0_2_1586;
   wire n_0_2_1587;
   wire n_0_2_1592;
   wire n_0_2_1593;
   wire n_0_2_1594;
   wire n_0_2_1596;
   wire n_0_2_1597;
   wire n_0_2_1599;
   wire n_0_2_1600;
   wire n_0_2_1601;
   wire n_0_2_1603;

   assign out_c[63] = out_c[16];
   assign out_c[62] = out_c[16];
   assign out_c[61] = out_c[16];
   assign out_c[60] = out_c[16];
   assign out_c[59] = out_c[16];
   assign out_c[58] = out_c[16];
   assign out_c[57] = out_c[16];
   assign out_c[56] = out_c[16];
   assign out_c[55] = out_c[16];
   assign out_c[54] = out_c[16];
   assign out_c[53] = out_c[16];
   assign out_c[52] = out_c[16];
   assign out_c[51] = out_c[16];
   assign out_c[50] = out_c[16];
   assign out_c[49] = out_c[16];
   assign out_c[48] = out_c[16];
   assign out_c[47] = out_c[16];
   assign out_c[46] = out_c[16];
   assign out_c[45] = out_c[16];
   assign out_c[44] = out_c[16];
   assign out_c[43] = out_c[16];
   assign out_c[42] = out_c[16];
   assign out_c[41] = out_c[16];
   assign out_c[40] = out_c[16];
   assign out_c[39] = out_c[16];
   assign out_c[38] = out_c[16];
   assign out_c[37] = out_c[16];
   assign out_c[36] = out_c[16];
   assign out_c[35] = out_c[16];
   assign out_c[34] = out_c[16];
   assign out_c[33] = out_c[16];
   assign out_c[32] = out_c[16];
   assign out_c[31] = out_c[16];
   assign out_c[30] = out_c[16];
   assign out_c[29] = out_c[16];
   assign out_c[28] = out_c[16];
   assign out_c[27] = out_c[16];
   assign out_c[26] = out_c[16];
   assign out_c[25] = out_c[16];
   assign out_c[24] = out_c[16];
   assign out_c[23] = out_c[16];
   assign out_c[22] = out_c[16];
   assign out_c[21] = out_c[16];
   assign out_c[20] = out_c[16];
   assign out_c[19] = out_c[16];
   assign out_c[18] = out_c[16];
   assign out_c[17] = out_c[16];

   DFFR_X1 posv_flag_reg (.D(n_0_40), .RN(n_0_39), .CK(n_0_0), .Q(posv), .QN());
   datapath i_0_1 (.in_b({in_b[22], in_b[21], in_b[20], in_b[19], in_b[18], 
      in_b[17], in_b[16], in_b[15], in_b[14], in_b[13], in_b[12], in_b[11], 
      in_b[10], in_b[9], in_b[8], in_b[7], in_b[6], in_b[5], in_b[4], in_b[3], 
      in_b[2], in_b[1], in_b[0]}), .p_0({n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, 
      n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, 
      n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, uc_0}));
   datapath__0_10 i_0_12 (.plus({n_0_38, uc_1, uc_2, uc_3, uc_4, uc_5, uc_6, 
      uc_7, uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, uc_15, uc_16, uc_17, 
      uc_18, uc_19, uc_20, uc_21, uc_22, uc_23, uc_24, uc_25, uc_26, uc_27, 
      uc_28, uc_29, uc_30, uc_31, uc_32, uc_33, uc_34, uc_35, uc_36, uc_37, 
      uc_38, uc_39, uc_40, uc_41, uc_42, uc_43, uc_44, uc_45, uc_46, uc_47, 
      n_0_37, n_0_36, n_0_35, n_0_34, n_0_33, n_0_32, n_0_31, n_0_30, n_0_29, 
      n_0_28, n_0_27, n_0_26, n_0_25, n_0_24, n_0_23, uc_48}), .p_0({1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, quotient[15], 
      quotient[14], quotient[13], quotient[12], quotient[11], quotient[10], 
      quotient[9], quotient[8], quotient[7], quotient[6], quotient[5], 
      quotient[4], quotient[3], quotient[2], quotient[1], quotient[0]}));
   DFFR_X1 zero_flag_reg (.D(n_0_41), .RN(n_0_39), .CK(n_0_0), .Q(zero), .QN());
   DFFR_X1 ovfl_flag_reg (.D(n_0_59), .RN(n_0_39), .CK(n_0_0), .Q(ovfl_flag), 
      .QN());
   DFFR_X1 divide_by_zero_error_reg (.D(n_0_58), .RN(n_0_39), .CK(n_0_0), 
      .Q(divide_by_zero_error), .QN());
   DFFR_X1 ready_reg (.D(1'b1), .RN(n_0_39), .CK(n_0_0), .Q(done), .QN());
   DFFR_X1 \out64_reg[63]  (.D(n_0_57), .RN(n_0_39), .CK(n_0_0), .Q(out_c[16]), 
      .QN());
   DFFR_X1 \out64_reg[15]  (.D(n_0_56), .RN(n_0_39), .CK(n_0_0), .Q(out_c[15]), 
      .QN());
   DFFR_X1 \out64_reg[14]  (.D(n_0_55), .RN(n_0_39), .CK(n_0_0), .Q(out_c[14]), 
      .QN());
   DFFR_X1 \out64_reg[13]  (.D(n_0_54), .RN(n_0_39), .CK(n_0_0), .Q(out_c[13]), 
      .QN());
   DFFR_X1 \out64_reg[12]  (.D(n_0_53), .RN(n_0_39), .CK(n_0_0), .Q(out_c[12]), 
      .QN());
   DFFR_X1 \out64_reg[11]  (.D(n_0_52), .RN(n_0_39), .CK(n_0_0), .Q(out_c[11]), 
      .QN());
   DFFR_X1 \out64_reg[10]  (.D(n_0_51), .RN(n_0_39), .CK(n_0_0), .Q(out_c[10]), 
      .QN());
   DFFR_X1 \out64_reg[9]  (.D(n_0_50), .RN(n_0_39), .CK(n_0_0), .Q(out_c[9]), 
      .QN());
   DFFR_X1 \out64_reg[8]  (.D(n_0_49), .RN(n_0_39), .CK(n_0_0), .Q(out_c[8]), 
      .QN());
   DFFR_X1 \out64_reg[7]  (.D(n_0_48), .RN(n_0_39), .CK(n_0_0), .Q(out_c[7]), 
      .QN());
   DFFR_X1 \out64_reg[6]  (.D(n_0_47), .RN(n_0_39), .CK(n_0_0), .Q(out_c[6]), 
      .QN());
   DFFR_X1 \out64_reg[5]  (.D(n_0_46), .RN(n_0_39), .CK(n_0_0), .Q(out_c[5]), 
      .QN());
   DFFR_X1 \out64_reg[4]  (.D(n_0_45), .RN(n_0_39), .CK(n_0_0), .Q(out_c[4]), 
      .QN());
   DFFR_X1 \out64_reg[3]  (.D(n_0_44), .RN(n_0_39), .CK(n_0_0), .Q(out_c[3]), 
      .QN());
   DFFR_X1 \out64_reg[2]  (.D(n_0_43), .RN(n_0_39), .CK(n_0_0), .Q(out_c[2]), 
      .QN());
   DFFR_X1 \out64_reg[1]  (.D(n_0_42), .RN(n_0_39), .CK(n_0_0), .Q(out_c[1]), 
      .QN());
   DFFR_X1 \out64_reg[0]  (.D(quotient[0]), .RN(n_0_39), .CK(n_0_0), .Q(out_c[0]), 
      .QN());
   INV_X1 i_0_0_0 (.A(rst), .ZN(n_0_39));
   CLKGATETST_X1 clk_gate_divide_by_zero_error_reg (.CK(clk), .E(enbl), .SE(1'b0), 
      .GCK(n_0_0));
   AOI22_X1 i_0_2_0 (.A1(n_0_2_778), .A2(n_0_2_774), .B1(n_0_2_775), .B2(
      n_0_2_1421), .ZN(n_0_2_57));
   OAI22_X1 i_0_2_1 (.A1(n_0_2_57), .A2(n_0_2_770), .B1(n_0_2_1044), .B2(
      n_0_2_772), .ZN(n_0_2_58));
   NAND2_X1 i_0_2_2 (.A1(n_0_2_58), .A2(n_0_2_1429), .ZN(n_0_2_59));
   INV_X1 i_0_2_3 (.A(n_0_2_58), .ZN(n_0_2_60));
   AOI22_X1 i_0_2_4 (.A1(n_0_2_59), .A2(n_0_2_769), .B1(n_0_2_60), .B2(
      n_0_2_1190), .ZN(n_0_2_61));
   XNOR2_X1 i_0_2_5 (.A(n_0_2_61), .B(n_0_2_1427), .ZN(n_0_2_62));
   NAND4_X1 i_0_2_6 (.A1(n_0_2_62), .A2(n_0_2_1196), .A3(n_0_2_1197), .A4(
      n_0_2_1431), .ZN(n_0_2_63));
   NAND4_X1 i_0_2_7 (.A1(n_0_2_62), .A2(n_0_2_56), .A3(n_0_2_287), .A4(
      n_0_2_1431), .ZN(n_0_2_64));
   NOR2_X1 i_0_2_8 (.A1(n_0_2_64), .A2(n_0_2_1438), .ZN(n_0_2_65));
   AOI22_X1 i_0_2_9 (.A1(n_0_2_63), .A2(n_0_2_799), .B1(n_0_2_65), .B2(
      n_0_2_1091), .ZN(n_0_2_66));
   OAI21_X1 i_0_2_10 (.A(n_0_2_1255), .B1(n_0_2_66), .B2(n_0_2_766), .ZN(
      n_0_2_67));
   INV_X1 i_0_2_11 (.A(n_0_2_65), .ZN(n_0_2_68));
   INV_X1 i_0_2_12 (.A(n_0_2_63), .ZN(n_0_2_69));
   OAI22_X1 i_0_2_13 (.A1(n_0_2_68), .A2(n_0_2_764), .B1(n_0_2_69), .B2(
      n_0_2_795), .ZN(n_0_2_70));
   OR2_X1 i_0_2_14 (.A1(n_0_2_70), .A2(n_0_2_54), .ZN(n_0_2_71));
   AOI22_X1 i_0_2_15 (.A1(n_0_2_67), .A2(n_0_2_71), .B1(n_0_2_70), .B2(n_0_2_54), 
      .ZN(n_0_2_72));
   AOI22_X1 i_0_2_16 (.A1(n_0_2_63), .A2(n_0_2_800), .B1(n_0_2_65), .B2(
      n_0_2_763), .ZN(n_0_2_73));
   AND2_X1 i_0_2_17 (.A1(n_0_2_73), .A2(n_0_2_1403), .ZN(n_0_2_74));
   OAI22_X1 i_0_2_18 (.A1(n_0_2_72), .A2(n_0_2_74), .B1(n_0_2_1403), .B2(
      n_0_2_73), .ZN(n_0_2_75));
   AOI22_X1 i_0_2_19 (.A1(n_0_2_63), .A2(n_0_2_806), .B1(n_0_2_65), .B2(
      n_0_2_762), .ZN(n_0_2_76));
   NOR2_X1 i_0_2_20 (.A1(n_0_2_76), .A2(n_0_2_1406), .ZN(n_0_2_77));
   INV_X1 i_0_2_21 (.A(n_0_2_76), .ZN(n_0_2_78));
   OAI22_X1 i_0_2_22 (.A1(n_0_2_75), .A2(n_0_2_77), .B1(n_0_2_147), .B2(n_0_2_78), 
      .ZN(n_0_2_79));
   AOI22_X1 i_0_2_23 (.A1(n_0_2_63), .A2(n_0_2_809), .B1(n_0_2_65), .B2(
      n_0_2_761), .ZN(n_0_2_80));
   AND2_X1 i_0_2_24 (.A1(n_0_2_80), .A2(n_0_2_1408), .ZN(n_0_2_81));
   OAI22_X1 i_0_2_25 (.A1(n_0_2_79), .A2(n_0_2_81), .B1(n_0_2_1408), .B2(
      n_0_2_80), .ZN(n_0_2_82));
   AOI22_X1 i_0_2_26 (.A1(n_0_2_63), .A2(n_0_2_812), .B1(n_0_2_65), .B2(
      n_0_2_760), .ZN(n_0_2_83));
   NOR2_X1 i_0_2_27 (.A1(n_0_2_83), .A2(n_0_2_1410), .ZN(n_0_2_84));
   INV_X1 i_0_2_28 (.A(n_0_2_83), .ZN(n_0_2_85));
   OAI22_X1 i_0_2_29 (.A1(n_0_2_82), .A2(n_0_2_84), .B1(n_0_2_281), .B2(n_0_2_85), 
      .ZN(n_0_2_86));
   AOI22_X1 i_0_2_30 (.A1(n_0_2_63), .A2(n_0_2_816), .B1(n_0_2_65), .B2(
      n_0_2_759), .ZN(n_0_2_87));
   AND2_X1 i_0_2_31 (.A1(n_0_2_87), .A2(n_0_2_1413), .ZN(n_0_2_88));
   OAI22_X1 i_0_2_32 (.A1(n_0_2_86), .A2(n_0_2_88), .B1(n_0_2_1413), .B2(
      n_0_2_87), .ZN(n_0_2_89));
   AOI22_X1 i_0_2_33 (.A1(n_0_2_63), .A2(n_0_2_820), .B1(n_0_2_65), .B2(
      n_0_2_758), .ZN(n_0_2_90));
   NOR2_X1 i_0_2_34 (.A1(n_0_2_90), .A2(n_0_2_1415), .ZN(n_0_2_91));
   INV_X1 i_0_2_35 (.A(n_0_2_90), .ZN(n_0_2_92));
   OAI22_X1 i_0_2_36 (.A1(n_0_2_89), .A2(n_0_2_91), .B1(n_0_2_453), .B2(n_0_2_92), 
      .ZN(n_0_2_93));
   AOI22_X1 i_0_2_37 (.A1(n_0_2_63), .A2(n_0_2_823), .B1(n_0_2_65), .B2(
      n_0_2_757), .ZN(n_0_2_94));
   AND2_X1 i_0_2_38 (.A1(n_0_2_94), .A2(n_0_2_1417), .ZN(n_0_2_95));
   OAI22_X1 i_0_2_39 (.A1(n_0_2_93), .A2(n_0_2_95), .B1(n_0_2_1417), .B2(
      n_0_2_94), .ZN(n_0_2_97));
   AOI22_X1 i_0_2_40 (.A1(n_0_2_63), .A2(n_0_2_828), .B1(n_0_2_65), .B2(
      n_0_2_756), .ZN(n_0_2_98));
   NAND2_X1 i_0_2_41 (.A1(n_0_2_98), .A2(n_0_2_1418), .ZN(n_0_2_99));
   INV_X1 i_0_2_42 (.A(n_0_2_98), .ZN(n_0_2_100));
   AOI22_X1 i_0_2_43 (.A1(n_0_2_97), .A2(n_0_2_99), .B1(n_0_2_660), .B2(
      n_0_2_100), .ZN(n_0_2_101));
   AOI22_X1 i_0_2_44 (.A1(n_0_2_63), .A2(n_0_2_831), .B1(n_0_2_65), .B2(
      n_0_2_755), .ZN(n_0_2_102));
   AND2_X1 i_0_2_45 (.A1(n_0_2_102), .A2(n_0_2_1440), .ZN(n_0_2_103));
   OAI22_X1 i_0_2_46 (.A1(n_0_2_101), .A2(n_0_2_103), .B1(n_0_2_1440), .B2(
      n_0_2_102), .ZN(n_0_2_104));
   AOI22_X1 i_0_2_47 (.A1(n_0_2_63), .A2(n_0_2_836), .B1(n_0_2_65), .B2(
      n_0_2_754), .ZN(n_0_2_105));
   NOR2_X1 i_0_2_48 (.A1(n_0_2_105), .A2(n_0_2_1421), .ZN(n_0_2_106));
   INV_X1 i_0_2_49 (.A(n_0_2_105), .ZN(n_0_2_107));
   OAI22_X1 i_0_2_50 (.A1(n_0_2_104), .A2(n_0_2_106), .B1(n_0_2_907), .B2(
      n_0_2_107), .ZN(n_0_2_108));
   XNOR2_X1 i_0_2_51 (.A(n_0_2_778), .B(n_0_2_753), .ZN(n_0_2_109));
   AOI22_X1 i_0_2_52 (.A1(n_0_2_63), .A2(n_0_2_776), .B1(n_0_2_65), .B2(
      n_0_2_109), .ZN(n_0_2_110));
   AND2_X1 i_0_2_53 (.A1(n_0_2_110), .A2(n_0_2_1424), .ZN(n_0_2_111));
   OAI22_X1 i_0_2_54 (.A1(n_0_2_108), .A2(n_0_2_111), .B1(n_0_2_1424), .B2(
      n_0_2_110), .ZN(n_0_2_112));
   XNOR2_X1 i_0_2_55 (.A(n_0_2_57), .B(n_0_2_752), .ZN(n_0_2_113));
   AOI22_X1 i_0_2_56 (.A1(n_0_2_63), .A2(n_0_2_772), .B1(n_0_2_65), .B2(
      n_0_2_113), .ZN(n_0_2_114));
   NOR2_X1 i_0_2_57 (.A1(n_0_2_114), .A2(n_0_2_1429), .ZN(n_0_2_115));
   INV_X1 i_0_2_58 (.A(n_0_2_114), .ZN(n_0_2_116));
   OAI22_X1 i_0_2_59 (.A1(n_0_2_112), .A2(n_0_2_115), .B1(n_0_2_1190), .B2(
      n_0_2_116), .ZN(n_0_2_117));
   XNOR2_X1 i_0_2_60 (.A(n_0_2_58), .B(n_0_2_751), .ZN(n_0_2_118));
   AOI22_X1 i_0_2_61 (.A1(n_0_2_63), .A2(n_0_2_769), .B1(n_0_2_65), .B2(
      n_0_2_118), .ZN(n_0_2_119));
   AND2_X1 i_0_2_62 (.A1(n_0_2_119), .A2(n_0_2_1427), .ZN(n_0_2_120));
   OAI22_X1 i_0_2_63 (.A1(n_0_2_117), .A2(n_0_2_120), .B1(n_0_2_119), .B2(
      n_0_2_1427), .ZN(n_0_2_121));
   XNOR2_X1 i_0_2_64 (.A(n_0_2_121), .B(n_0_2_1428), .ZN(n_0_2_122));
   NOR2_X1 i_0_2_65 (.A1(n_0_2_122), .A2(n_0_2_750), .ZN(n_0_2_123));
   OAI221_X1 i_0_2_66 (.A(n_0_2_123), .B1(n_0_2_767), .B2(n_0_2_1398), .C1(
      n_0_2_1247), .C2(n_0_2_49), .ZN(n_0_2_124));
   XNOR2_X1 i_0_2_67 (.A(n_0_2_124), .B(n_0_2_66), .ZN(n_0_2_125));
   INV_X1 i_0_2_68 (.A(n_0_2_123), .ZN(n_0_2_126));
   AOI22_X1 i_0_2_69 (.A1(in_a[0]), .A2(n_0_2_126), .B1(n_0_2_123), .B2(
      n_0_2_1246), .ZN(n_0_2_127));
   OAI21_X1 i_0_2_70 (.A(n_0_2_1412), .B1(n_0_2_127), .B2(n_0_2_1366), .ZN(
      n_0_2_128));
   NOR2_X1 i_0_2_71 (.A1(n_0_2_128), .A2(n_0_2_54), .ZN(n_0_2_129));
   INV_X1 i_0_2_72 (.A(n_0_2_128), .ZN(n_0_2_130));
   OAI22_X1 i_0_2_73 (.A1(n_0_2_125), .A2(n_0_2_129), .B1(n_0_2_1400), .B2(
      n_0_2_130), .ZN(n_0_2_131));
   INV_X1 i_0_2_74 (.A(n_0_2_67), .ZN(n_0_2_132));
   OAI221_X1 i_0_2_75 (.A(n_0_2_123), .B1(n_0_2_54), .B2(n_0_2_67), .C1(
      n_0_2_1400), .C2(n_0_2_132), .ZN(n_0_2_133));
   XNOR2_X1 i_0_2_76 (.A(n_0_2_133), .B(n_0_2_70), .ZN(n_0_2_134));
   INV_X1 i_0_2_77 (.A(n_0_2_134), .ZN(n_0_2_135));
   NOR2_X1 i_0_2_78 (.A1(n_0_2_135), .A2(n_0_2_1403), .ZN(n_0_2_136));
   OAI22_X1 i_0_2_79 (.A1(n_0_2_131), .A2(n_0_2_136), .B1(n_0_2_96), .B2(
      n_0_2_134), .ZN(n_0_2_137));
   INV_X1 i_0_2_80 (.A(n_0_2_72), .ZN(n_0_2_138));
   OAI221_X1 i_0_2_81 (.A(n_0_2_123), .B1(n_0_2_1403), .B2(n_0_2_72), .C1(
      n_0_2_96), .C2(n_0_2_138), .ZN(n_0_2_139));
   XOR2_X1 i_0_2_82 (.A(n_0_2_139), .B(n_0_2_73), .Z(n_0_2_140));
   NOR2_X1 i_0_2_83 (.A1(n_0_2_140), .A2(n_0_2_147), .ZN(n_0_2_141));
   INV_X1 i_0_2_84 (.A(n_0_2_140), .ZN(n_0_2_142));
   OAI22_X1 i_0_2_85 (.A1(n_0_2_137), .A2(n_0_2_141), .B1(n_0_2_1406), .B2(
      n_0_2_142), .ZN(n_0_2_143));
   INV_X1 i_0_2_86 (.A(n_0_2_75), .ZN(n_0_2_144));
   OAI221_X1 i_0_2_87 (.A(n_0_2_123), .B1(n_0_2_1406), .B2(n_0_2_144), .C1(
      n_0_2_147), .C2(n_0_2_75), .ZN(n_0_2_145));
   XOR2_X1 i_0_2_88 (.A(n_0_2_145), .B(n_0_2_76), .Z(n_0_2_146));
   INV_X1 i_0_2_89 (.A(n_0_2_146), .ZN(n_0_2_148));
   NOR2_X1 i_0_2_90 (.A1(n_0_2_148), .A2(n_0_2_1408), .ZN(n_0_2_149));
   OAI22_X1 i_0_2_91 (.A1(n_0_2_143), .A2(n_0_2_149), .B1(n_0_2_146), .B2(
      n_0_2_209), .ZN(n_0_2_150));
   INV_X1 i_0_2_92 (.A(n_0_2_79), .ZN(n_0_2_151));
   OAI221_X1 i_0_2_93 (.A(n_0_2_123), .B1(n_0_2_1408), .B2(n_0_2_79), .C1(
      n_0_2_209), .C2(n_0_2_151), .ZN(n_0_2_152));
   XOR2_X1 i_0_2_94 (.A(n_0_2_152), .B(n_0_2_80), .Z(n_0_2_153));
   NOR2_X1 i_0_2_95 (.A1(n_0_2_153), .A2(n_0_2_281), .ZN(n_0_2_155));
   INV_X1 i_0_2_96 (.A(n_0_2_153), .ZN(n_0_2_156));
   OAI22_X1 i_0_2_97 (.A1(n_0_2_150), .A2(n_0_2_155), .B1(n_0_2_1410), .B2(
      n_0_2_156), .ZN(n_0_2_157));
   INV_X1 i_0_2_98 (.A(n_0_2_82), .ZN(n_0_2_158));
   OAI221_X1 i_0_2_99 (.A(n_0_2_123), .B1(n_0_2_1410), .B2(n_0_2_158), .C1(
      n_0_2_281), .C2(n_0_2_82), .ZN(n_0_2_159));
   XOR2_X1 i_0_2_100 (.A(n_0_2_159), .B(n_0_2_83), .Z(n_0_2_160));
   INV_X1 i_0_2_101 (.A(n_0_2_160), .ZN(n_0_2_161));
   NAND2_X1 i_0_2_102 (.A1(n_0_2_161), .A2(n_0_2_1413), .ZN(n_0_2_162));
   AOI22_X1 i_0_2_103 (.A1(n_0_2_157), .A2(n_0_2_162), .B1(n_0_2_160), .B2(
      n_0_2_363), .ZN(n_0_2_163));
   INV_X1 i_0_2_104 (.A(n_0_2_86), .ZN(n_0_2_164));
   OAI221_X1 i_0_2_105 (.A(n_0_2_123), .B1(n_0_2_1413), .B2(n_0_2_86), .C1(
      n_0_2_363), .C2(n_0_2_164), .ZN(n_0_2_165));
   XOR2_X1 i_0_2_106 (.A(n_0_2_165), .B(n_0_2_87), .Z(n_0_2_166));
   NOR2_X1 i_0_2_107 (.A1(n_0_2_166), .A2(n_0_2_453), .ZN(n_0_2_167));
   INV_X1 i_0_2_108 (.A(n_0_2_166), .ZN(n_0_2_168));
   OAI22_X1 i_0_2_109 (.A1(n_0_2_163), .A2(n_0_2_167), .B1(n_0_2_1415), .B2(
      n_0_2_168), .ZN(n_0_2_169));
   INV_X1 i_0_2_110 (.A(n_0_2_89), .ZN(n_0_2_170));
   OAI221_X1 i_0_2_111 (.A(n_0_2_123), .B1(n_0_2_1415), .B2(n_0_2_170), .C1(
      n_0_2_453), .C2(n_0_2_89), .ZN(n_0_2_171));
   XOR2_X1 i_0_2_112 (.A(n_0_2_171), .B(n_0_2_90), .Z(n_0_2_172));
   INV_X1 i_0_2_113 (.A(n_0_2_172), .ZN(n_0_2_173));
   NOR2_X1 i_0_2_114 (.A1(n_0_2_173), .A2(n_0_2_1417), .ZN(n_0_2_174));
   OAI22_X1 i_0_2_115 (.A1(n_0_2_169), .A2(n_0_2_174), .B1(n_0_2_172), .B2(
      n_0_2_458), .ZN(n_0_2_175));
   INV_X1 i_0_2_116 (.A(n_0_2_93), .ZN(n_0_2_176));
   OAI221_X1 i_0_2_117 (.A(n_0_2_123), .B1(n_0_2_1417), .B2(n_0_2_93), .C1(
      n_0_2_458), .C2(n_0_2_176), .ZN(n_0_2_177));
   XOR2_X1 i_0_2_118 (.A(n_0_2_177), .B(n_0_2_94), .Z(n_0_2_178));
   NOR2_X1 i_0_2_119 (.A1(n_0_2_178), .A2(n_0_2_660), .ZN(n_0_2_179));
   INV_X1 i_0_2_120 (.A(n_0_2_178), .ZN(n_0_2_180));
   OAI22_X1 i_0_2_121 (.A1(n_0_2_175), .A2(n_0_2_179), .B1(n_0_2_1418), .B2(
      n_0_2_180), .ZN(n_0_2_181));
   INV_X1 i_0_2_122 (.A(n_0_2_97), .ZN(n_0_2_182));
   OAI221_X1 i_0_2_123 (.A(n_0_2_123), .B1(n_0_2_1418), .B2(n_0_2_182), .C1(
      n_0_2_660), .C2(n_0_2_97), .ZN(n_0_2_183));
   XOR2_X1 i_0_2_124 (.A(n_0_2_183), .B(n_0_2_98), .Z(n_0_2_184));
   INV_X1 i_0_2_125 (.A(n_0_2_184), .ZN(n_0_2_185));
   NOR2_X1 i_0_2_126 (.A1(n_0_2_185), .A2(n_0_2_1440), .ZN(n_0_2_186));
   OAI22_X1 i_0_2_127 (.A1(n_0_2_181), .A2(n_0_2_186), .B1(n_0_2_780), .B2(
      n_0_2_184), .ZN(n_0_2_187));
   INV_X1 i_0_2_128 (.A(n_0_2_101), .ZN(n_0_2_188));
   OAI221_X1 i_0_2_129 (.A(n_0_2_123), .B1(n_0_2_1440), .B2(n_0_2_101), .C1(
      n_0_2_780), .C2(n_0_2_188), .ZN(n_0_2_189));
   XOR2_X1 i_0_2_130 (.A(n_0_2_189), .B(n_0_2_102), .Z(n_0_2_190));
   NOR2_X1 i_0_2_131 (.A1(n_0_2_190), .A2(n_0_2_907), .ZN(n_0_2_191));
   INV_X1 i_0_2_132 (.A(n_0_2_190), .ZN(n_0_2_192));
   OAI22_X1 i_0_2_133 (.A1(n_0_2_187), .A2(n_0_2_191), .B1(n_0_2_1421), .B2(
      n_0_2_192), .ZN(n_0_2_193));
   INV_X1 i_0_2_134 (.A(n_0_2_104), .ZN(n_0_2_194));
   OAI221_X1 i_0_2_135 (.A(n_0_2_123), .B1(n_0_2_1421), .B2(n_0_2_194), .C1(
      n_0_2_907), .C2(n_0_2_104), .ZN(n_0_2_195));
   XOR2_X1 i_0_2_136 (.A(n_0_2_195), .B(n_0_2_105), .Z(n_0_2_196));
   OR2_X1 i_0_2_137 (.A1(n_0_2_196), .A2(n_0_2_1044), .ZN(n_0_2_197));
   AOI22_X1 i_0_2_138 (.A1(n_0_2_193), .A2(n_0_2_197), .B1(n_0_2_196), .B2(
      n_0_2_1044), .ZN(n_0_2_198));
   INV_X1 i_0_2_139 (.A(n_0_2_108), .ZN(n_0_2_199));
   OAI221_X1 i_0_2_140 (.A(n_0_2_123), .B1(n_0_2_108), .B2(n_0_2_1424), .C1(
      n_0_2_1044), .C2(n_0_2_199), .ZN(n_0_2_200));
   XOR2_X1 i_0_2_141 (.A(n_0_2_200), .B(n_0_2_110), .Z(n_0_2_201));
   NAND2_X1 i_0_2_142 (.A1(n_0_2_201), .A2(n_0_2_1190), .ZN(n_0_2_202));
   INV_X1 i_0_2_143 (.A(n_0_2_201), .ZN(n_0_2_203));
   AOI22_X1 i_0_2_144 (.A1(n_0_2_198), .A2(n_0_2_202), .B1(n_0_2_203), .B2(
      n_0_2_1429), .ZN(n_0_2_204));
   INV_X1 i_0_2_145 (.A(n_0_2_112), .ZN(n_0_2_205));
   OAI221_X1 i_0_2_146 (.A(n_0_2_123), .B1(n_0_2_1429), .B2(n_0_2_205), .C1(
      n_0_2_1190), .C2(n_0_2_112), .ZN(n_0_2_206));
   XOR2_X1 i_0_2_147 (.A(n_0_2_206), .B(n_0_2_114), .Z(n_0_2_207));
   INV_X1 i_0_2_148 (.A(n_0_2_207), .ZN(n_0_2_208));
   NOR2_X1 i_0_2_149 (.A1(n_0_2_208), .A2(n_0_2_1427), .ZN(n_0_2_210));
   OAI22_X1 i_0_2_150 (.A1(n_0_2_204), .A2(n_0_2_210), .B1(n_0_2_1352), .B2(
      n_0_2_207), .ZN(n_0_2_211));
   INV_X1 i_0_2_151 (.A(n_0_2_117), .ZN(n_0_2_212));
   OAI221_X1 i_0_2_152 (.A(n_0_2_123), .B1(n_0_2_1427), .B2(n_0_2_117), .C1(
      n_0_2_1352), .C2(n_0_2_212), .ZN(n_0_2_213));
   XNOR2_X1 i_0_2_153 (.A(n_0_2_213), .B(n_0_2_119), .ZN(n_0_2_214));
   AND2_X1 i_0_2_154 (.A1(n_0_2_214), .A2(n_0_2_1428), .ZN(n_0_2_215));
   OAI22_X1 i_0_2_155 (.A1(n_0_2_211), .A2(n_0_2_215), .B1(n_0_2_1428), .B2(
      n_0_2_214), .ZN(n_0_2_216));
   OAI21_X1 i_0_2_156 (.A(n_0_2_1431), .B1(n_0_2_216), .B2(n_0_2_1434), .ZN(
      n_0_2_217));
   AOI21_X1 i_0_2_157 (.A(n_0_2_217), .B1(n_0_2_1434), .B2(n_0_2_216), .ZN(
      n_0_2_218));
   INV_X1 i_0_2_158 (.A(n_0_2_218), .ZN(n_0_2_219));
   NOR2_X1 i_0_2_159 (.A1(n_0_2_219), .A2(n_0_2_51), .ZN(n_0_2_220));
   NAND2_X1 i_0_2_160 (.A1(n_0_2_220), .A2(in_b[0]), .ZN(n_0_2_221));
   INV_X1 i_0_2_161 (.A(n_0_2_221), .ZN(n_0_2_1522));
   INV_X1 i_0_2_162 (.A(n_0_2_220), .ZN(n_0_2_222));
   NAND2_X1 i_0_2_163 (.A1(n_0_2_127), .A2(n_0_2_749), .ZN(n_0_2_223));
   OAI21_X1 i_0_2_164 (.A(n_0_2_223), .B1(n_0_2_127), .B2(n_0_2_749), .ZN(
      n_0_2_224));
   NAND2_X1 i_0_2_165 (.A1(n_0_2_218), .A2(n_0_2_154), .ZN(n_0_2_225));
   INV_X1 i_0_2_166 (.A(n_0_2_225), .ZN(n_0_2_226));
   OAI22_X1 i_0_2_167 (.A1(n_0_2_222), .A2(n_0_2_224), .B1(n_0_2_226), .B2(
      n_0_2_127), .ZN(n_0_2_1525));
   INV_X1 i_0_2_168 (.A(n_0_2_1525), .ZN(n_0_2_227));
   AOI22_X1 i_0_2_169 (.A1(n_0_2_1525), .A2(n_0_2_54), .B1(n_0_2_227), .B2(
      n_0_2_1400), .ZN(n_0_2_228));
   AOI21_X1 i_0_2_170 (.A(n_0_2_1397), .B1(n_0_2_1522), .B2(n_0_2_1367), 
      .ZN(n_0_2_229));
   XNOR2_X1 i_0_2_171 (.A(n_0_2_228), .B(n_0_2_229), .ZN(n_0_2_1579));
   OAI22_X1 i_0_2_172 (.A1(n_0_2_1522), .A2(n_0_2_749), .B1(n_0_2_221), .B2(
      n_0_2_748), .ZN(n_0_2_1573));
   XNOR2_X1 i_0_2_173 (.A(n_0_2_214), .B(n_0_2_1428), .ZN(n_0_2_230));
   XNOR2_X1 i_0_2_174 (.A(n_0_2_211), .B(n_0_2_230), .ZN(n_0_2_231));
   OAI22_X1 i_0_2_175 (.A1(n_0_2_222), .A2(n_0_2_231), .B1(n_0_2_226), .B2(
      n_0_2_214), .ZN(n_0_2_1570));
   NAND2_X1 i_0_2_176 (.A1(n_0_2_1570), .A2(n_0_2_52), .ZN(n_0_2_0));
   XNOR2_X1 i_0_2_177 (.A(n_0_2_1570), .B(n_0_2_1434), .ZN(n_0_2_1));
   OAI22_X1 i_0_2_178 (.A1(n_0_2_208), .A2(n_0_2_1352), .B1(n_0_2_207), .B2(
      n_0_2_1427), .ZN(n_0_2_232));
   XNOR2_X1 i_0_2_179 (.A(n_0_2_204), .B(n_0_2_232), .ZN(n_0_2_233));
   OAI22_X1 i_0_2_180 (.A1(n_0_2_222), .A2(n_0_2_233), .B1(n_0_2_226), .B2(
      n_0_2_208), .ZN(n_0_2_1567));
   NAND2_X1 i_0_2_181 (.A1(n_0_2_1567), .A2(n_0_2_1516), .ZN(n_0_2_2));
   XNOR2_X1 i_0_2_182 (.A(n_0_2_1567), .B(n_0_2_1428), .ZN(n_0_2_3));
   AOI22_X1 i_0_2_183 (.A1(n_0_2_201), .A2(n_0_2_1190), .B1(n_0_2_203), .B2(
      n_0_2_1429), .ZN(n_0_2_234));
   XNOR2_X1 i_0_2_184 (.A(n_0_2_198), .B(n_0_2_234), .ZN(n_0_2_235));
   AOI22_X1 i_0_2_185 (.A1(n_0_2_220), .A2(n_0_2_235), .B1(n_0_2_225), .B2(
      n_0_2_201), .ZN(n_0_2_236));
   INV_X1 i_0_2_186 (.A(n_0_2_236), .ZN(n_0_2_1564));
   NAND2_X1 i_0_2_187 (.A1(n_0_2_1564), .A2(n_0_2_1352), .ZN(n_0_2_4));
   OAI22_X1 i_0_2_188 (.A1(n_0_2_1564), .A2(n_0_2_1427), .B1(n_0_2_236), 
      .B2(n_0_2_1352), .ZN(n_0_2_5));
   XOR2_X1 i_0_2_189 (.A(n_0_2_196), .B(n_0_2_1424), .Z(n_0_2_237));
   XNOR2_X1 i_0_2_190 (.A(n_0_2_193), .B(n_0_2_237), .ZN(n_0_2_238));
   AOI22_X1 i_0_2_191 (.A1(n_0_2_220), .A2(n_0_2_238), .B1(n_0_2_225), .B2(
      n_0_2_196), .ZN(n_0_2_239));
   INV_X1 i_0_2_192 (.A(n_0_2_239), .ZN(n_0_2_1561));
   NAND2_X1 i_0_2_193 (.A1(n_0_2_1561), .A2(n_0_2_1190), .ZN(n_0_2_6));
   OAI22_X1 i_0_2_194 (.A1(n_0_2_1561), .A2(n_0_2_1429), .B1(n_0_2_239), 
      .B2(n_0_2_1190), .ZN(n_0_2_7));
   OAI22_X1 i_0_2_195 (.A1(n_0_2_192), .A2(n_0_2_1421), .B1(n_0_2_190), .B2(
      n_0_2_907), .ZN(n_0_2_240));
   XNOR2_X1 i_0_2_196 (.A(n_0_2_187), .B(n_0_2_240), .ZN(n_0_2_241));
   OAI22_X1 i_0_2_197 (.A1(n_0_2_222), .A2(n_0_2_241), .B1(n_0_2_226), .B2(
      n_0_2_192), .ZN(n_0_2_1558));
   NAND2_X1 i_0_2_198 (.A1(n_0_2_1558), .A2(n_0_2_1044), .ZN(n_0_2_8));
   XNOR2_X1 i_0_2_199 (.A(n_0_2_1558), .B(n_0_2_1424), .ZN(n_0_2_9));
   AOI22_X1 i_0_2_200 (.A1(n_0_2_184), .A2(n_0_2_1440), .B1(n_0_2_185), .B2(
      n_0_2_780), .ZN(n_0_2_242));
   XNOR2_X1 i_0_2_201 (.A(n_0_2_181), .B(n_0_2_242), .ZN(n_0_2_243));
   AOI22_X1 i_0_2_202 (.A1(n_0_2_220), .A2(n_0_2_243), .B1(n_0_2_225), .B2(
      n_0_2_184), .ZN(n_0_2_244));
   INV_X1 i_0_2_203 (.A(n_0_2_244), .ZN(n_0_2_1555));
   NAND2_X1 i_0_2_204 (.A1(n_0_2_1555), .A2(n_0_2_907), .ZN(n_0_2_10));
   OAI22_X1 i_0_2_205 (.A1(n_0_2_1555), .A2(n_0_2_1421), .B1(n_0_2_244), 
      .B2(n_0_2_907), .ZN(n_0_2_11));
   XNOR2_X1 i_0_2_206 (.A(n_0_2_178), .B(n_0_2_1418), .ZN(n_0_2_245));
   XNOR2_X1 i_0_2_207 (.A(n_0_2_175), .B(n_0_2_245), .ZN(n_0_2_246));
   AOI22_X1 i_0_2_208 (.A1(n_0_2_220), .A2(n_0_2_246), .B1(n_0_2_225), .B2(
      n_0_2_178), .ZN(n_0_2_247));
   INV_X1 i_0_2_209 (.A(n_0_2_247), .ZN(n_0_2_1552));
   NAND2_X1 i_0_2_210 (.A1(n_0_2_1552), .A2(n_0_2_780), .ZN(n_0_2_12));
   OAI22_X1 i_0_2_211 (.A1(n_0_2_1552), .A2(n_0_2_1440), .B1(n_0_2_247), 
      .B2(n_0_2_780), .ZN(n_0_2_13));
   OAI22_X1 i_0_2_212 (.A1(n_0_2_173), .A2(n_0_2_458), .B1(n_0_2_172), .B2(
      n_0_2_1417), .ZN(n_0_2_248));
   XNOR2_X1 i_0_2_213 (.A(n_0_2_169), .B(n_0_2_248), .ZN(n_0_2_249));
   OAI22_X1 i_0_2_214 (.A1(n_0_2_222), .A2(n_0_2_249), .B1(n_0_2_226), .B2(
      n_0_2_173), .ZN(n_0_2_1549));
   NAND2_X1 i_0_2_215 (.A1(n_0_2_1549), .A2(n_0_2_660), .ZN(n_0_2_14));
   XNOR2_X1 i_0_2_216 (.A(n_0_2_1549), .B(n_0_2_1418), .ZN(n_0_2_15));
   XNOR2_X1 i_0_2_217 (.A(n_0_2_166), .B(n_0_2_1415), .ZN(n_0_2_250));
   XNOR2_X1 i_0_2_218 (.A(n_0_2_163), .B(n_0_2_250), .ZN(n_0_2_251));
   AOI22_X1 i_0_2_219 (.A1(n_0_2_220), .A2(n_0_2_251), .B1(n_0_2_225), .B2(
      n_0_2_166), .ZN(n_0_2_252));
   INV_X1 i_0_2_220 (.A(n_0_2_252), .ZN(n_0_2_1546));
   NAND2_X1 i_0_2_221 (.A1(n_0_2_1546), .A2(n_0_2_458), .ZN(n_0_2_16));
   OAI22_X1 i_0_2_222 (.A1(n_0_2_1546), .A2(n_0_2_1417), .B1(n_0_2_252), 
      .B2(n_0_2_458), .ZN(n_0_2_17));
   OAI22_X1 i_0_2_223 (.A1(n_0_2_161), .A2(n_0_2_363), .B1(n_0_2_160), .B2(
      n_0_2_1413), .ZN(n_0_2_253));
   XNOR2_X1 i_0_2_224 (.A(n_0_2_157), .B(n_0_2_253), .ZN(n_0_2_254));
   OAI22_X1 i_0_2_225 (.A1(n_0_2_222), .A2(n_0_2_254), .B1(n_0_2_226), .B2(
      n_0_2_161), .ZN(n_0_2_1543));
   NAND2_X1 i_0_2_226 (.A1(n_0_2_1543), .A2(n_0_2_453), .ZN(n_0_2_18));
   XNOR2_X1 i_0_2_227 (.A(n_0_2_1543), .B(n_0_2_1415), .ZN(n_0_2_19));
   AOI22_X1 i_0_2_228 (.A1(n_0_2_153), .A2(n_0_2_281), .B1(n_0_2_156), .B2(
      n_0_2_1410), .ZN(n_0_2_255));
   XNOR2_X1 i_0_2_229 (.A(n_0_2_150), .B(n_0_2_255), .ZN(n_0_2_256));
   AOI22_X1 i_0_2_230 (.A1(n_0_2_220), .A2(n_0_2_256), .B1(n_0_2_225), .B2(
      n_0_2_153), .ZN(n_0_2_257));
   INV_X1 i_0_2_231 (.A(n_0_2_257), .ZN(n_0_2_1540));
   NAND2_X1 i_0_2_232 (.A1(n_0_2_1540), .A2(n_0_2_363), .ZN(n_0_2_20));
   OAI22_X1 i_0_2_233 (.A1(n_0_2_1540), .A2(n_0_2_1413), .B1(n_0_2_257), 
      .B2(n_0_2_363), .ZN(n_0_2_21));
   AOI22_X1 i_0_2_234 (.A1(n_0_2_146), .A2(n_0_2_1408), .B1(n_0_2_148), .B2(
      n_0_2_209), .ZN(n_0_2_258));
   XNOR2_X1 i_0_2_235 (.A(n_0_2_143), .B(n_0_2_258), .ZN(n_0_2_259));
   AOI22_X1 i_0_2_236 (.A1(n_0_2_220), .A2(n_0_2_259), .B1(n_0_2_225), .B2(
      n_0_2_146), .ZN(n_0_2_260));
   INV_X1 i_0_2_237 (.A(n_0_2_260), .ZN(n_0_2_1537));
   NAND2_X1 i_0_2_238 (.A1(n_0_2_1537), .A2(n_0_2_281), .ZN(n_0_2_22));
   OAI22_X1 i_0_2_239 (.A1(n_0_2_1537), .A2(n_0_2_1410), .B1(n_0_2_260), 
      .B2(n_0_2_281), .ZN(n_0_2_23));
   AOI22_X1 i_0_2_240 (.A1(n_0_2_140), .A2(n_0_2_147), .B1(n_0_2_142), .B2(
      n_0_2_1406), .ZN(n_0_2_261));
   XNOR2_X1 i_0_2_241 (.A(n_0_2_137), .B(n_0_2_261), .ZN(n_0_2_262));
   AOI22_X1 i_0_2_242 (.A1(n_0_2_220), .A2(n_0_2_262), .B1(n_0_2_225), .B2(
      n_0_2_140), .ZN(n_0_2_263));
   INV_X1 i_0_2_243 (.A(n_0_2_263), .ZN(n_0_2_1534));
   NAND2_X1 i_0_2_244 (.A1(n_0_2_1534), .A2(n_0_2_209), .ZN(n_0_2_1602));
   OAI22_X1 i_0_2_245 (.A1(n_0_2_1534), .A2(n_0_2_1408), .B1(n_0_2_263), 
      .B2(n_0_2_209), .ZN(n_0_2_1598));
   AOI22_X1 i_0_2_246 (.A1(n_0_2_134), .A2(n_0_2_1403), .B1(n_0_2_135), .B2(
      n_0_2_96), .ZN(n_0_2_264));
   XNOR2_X1 i_0_2_247 (.A(n_0_2_264), .B(n_0_2_131), .ZN(n_0_2_265));
   AOI22_X1 i_0_2_248 (.A1(n_0_2_220), .A2(n_0_2_265), .B1(n_0_2_225), .B2(
      n_0_2_134), .ZN(n_0_2_266));
   INV_X1 i_0_2_249 (.A(n_0_2_266), .ZN(n_0_2_1531));
   NAND2_X1 i_0_2_250 (.A1(n_0_2_1531), .A2(n_0_2_147), .ZN(n_0_2_1595));
   OAI22_X1 i_0_2_251 (.A1(n_0_2_1531), .A2(n_0_2_1406), .B1(n_0_2_266), 
      .B2(n_0_2_147), .ZN(n_0_2_1591));
   NAND2_X1 i_0_2_252 (.A1(n_0_2_1525), .A2(n_0_2_54), .ZN(n_0_2_267));
   AOI22_X1 i_0_2_253 (.A1(n_0_2_267), .A2(n_0_2_229), .B1(n_0_2_1400), .B2(
      n_0_2_227), .ZN(n_0_2_268));
   NAND2_X1 i_0_2_254 (.A1(n_0_2_268), .A2(n_0_2_96), .ZN(n_0_2_1590));
   INV_X1 i_0_2_255 (.A(n_0_2_125), .ZN(n_0_2_269));
   AOI22_X1 i_0_2_256 (.A1(n_0_2_269), .A2(n_0_2_1400), .B1(n_0_2_125), .B2(
      n_0_2_54), .ZN(n_0_2_270));
   XOR2_X1 i_0_2_257 (.A(n_0_2_270), .B(n_0_2_128), .Z(n_0_2_271));
   OAI22_X1 i_0_2_258 (.A1(n_0_2_222), .A2(n_0_2_271), .B1(n_0_2_226), .B2(
      n_0_2_125), .ZN(n_0_2_1528));
   NAND2_X1 i_0_2_259 (.A1(n_0_2_1528), .A2(n_0_2_96), .ZN(n_0_2_1588));
   NAND2_X1 i_0_2_260 (.A1(n_0_2_268), .A2(n_0_2_1528), .ZN(n_0_2_1589));
   OAI21_X1 i_0_2_261 (.A(n_0_2_1589), .B1(n_0_2_268), .B2(n_0_2_1528), .ZN(
      n_0_2_272));
   XNOR2_X1 i_0_2_262 (.A(n_0_2_272), .B(n_0_2_1403), .ZN(n_0_2_1585));
   NAND2_X1 i_0_2_263 (.A1(n_0_2_65), .A2(n_0_2_1394), .ZN(n_0_2_273));
   INV_X1 i_0_2_264 (.A(n_0_2_273), .ZN(quotient[8]));
   AOI22_X1 i_0_2_265 (.A1(n_0_2_273), .A2(n_0_2_846), .B1(n_0_2_1443), .B2(
      n_0_2_847), .ZN(n_0_49));
   NAND2_X1 i_0_2_266 (.A1(n_0_2_123), .A2(n_0_2_1394), .ZN(n_0_2_274));
   INV_X1 i_0_2_267 (.A(n_0_2_274), .ZN(quotient[7]));
   AOI22_X1 i_0_2_268 (.A1(n_0_2_274), .A2(n_0_2_846), .B1(n_0_2_847), .B2(
      n_0_2_1442), .ZN(n_0_48));
   NOR4_X1 i_0_2_269 (.A1(n_0_48), .A2(n_0_55), .A3(n_0_57), .A4(n_0_56), 
      .ZN(n_0_2_275));
   NAND3_X1 i_0_2_270 (.A1(n_0_2_275), .A2(n_0_2_747), .A3(n_0_2_746), .ZN(
      n_0_2_276));
   NOR3_X1 i_0_2_271 (.A1(n_0_2_276), .A2(n_0_50), .A3(n_0_49), .ZN(n_0_41));
   NOR3_X1 i_0_2_272 (.A1(n_0_41), .A2(n_0_56), .A3(n_0_2_48), .ZN(n_0_40));
   NAND2_X1 i_0_2_273 (.A1(n_0_2_220), .A2(n_0_2_1394), .ZN(n_0_2_277));
   AOI22_X1 i_0_2_274 (.A1(n_0_2_277), .A2(n_0_2_846), .B1(n_0_2_1441), .B2(
      n_0_2_847), .ZN(n_0_47));
   INV_X1 i_0_2_275 (.A(n_0_2_277), .ZN(quotient[6]));
   XNOR2_X1 i_0_2_276 (.A(n_0_2_1433), .B(n_0_2_24), .ZN(n_0_2_278));
   XOR2_X1 i_0_2_277 (.A(n_0_2_1439), .B(n_0_2_44), .Z(n_0_2_279));
   XNOR2_X1 i_0_2_278 (.A(n_0_2_1438), .B(n_0_2_43), .ZN(n_0_2_280));
   XOR2_X1 i_0_2_279 (.A(n_0_2_1436), .B(n_0_2_42), .Z(n_0_2_282));
   XNOR2_X1 i_0_2_280 (.A(n_0_2_1434), .B(n_0_2_41), .ZN(n_0_2_283));
   XOR2_X1 i_0_2_281 (.A(n_0_2_1428), .B(n_0_2_40), .Z(n_0_2_284));
   XNOR2_X1 i_0_2_282 (.A(n_0_2_1427), .B(n_0_2_39), .ZN(n_0_2_285));
   XOR2_X1 i_0_2_283 (.A(n_0_2_1429), .B(n_0_2_38), .Z(n_0_2_286));
   XNOR2_X1 i_0_2_284 (.A(n_0_2_1424), .B(n_0_2_37), .ZN(n_0_2_288));
   XOR2_X1 i_0_2_285 (.A(n_0_2_1421), .B(n_0_2_36), .Z(n_0_2_289));
   XNOR2_X1 i_0_2_286 (.A(n_0_2_1440), .B(n_0_2_35), .ZN(n_0_2_290));
   XOR2_X1 i_0_2_287 (.A(n_0_2_1418), .B(n_0_2_34), .Z(n_0_2_291));
   XNOR2_X1 i_0_2_288 (.A(n_0_2_1417), .B(n_0_2_33), .ZN(n_0_2_292));
   XOR2_X1 i_0_2_289 (.A(n_0_2_1415), .B(n_0_2_32), .Z(n_0_2_293));
   XNOR2_X1 i_0_2_290 (.A(n_0_2_1413), .B(n_0_2_31), .ZN(n_0_2_294));
   XOR2_X1 i_0_2_291 (.A(n_0_2_1410), .B(n_0_2_30), .Z(n_0_2_295));
   XNOR2_X1 i_0_2_292 (.A(n_0_2_318), .B(n_0_2_297), .ZN(n_0_2_296));
   XNOR2_X1 i_0_2_293 (.A(n_0_2_1408), .B(n_0_2_29), .ZN(n_0_2_297));
   XNOR2_X1 i_0_2_294 (.A(n_0_2_321), .B(n_0_2_299), .ZN(n_0_2_298));
   XOR2_X1 i_0_2_295 (.A(n_0_2_1406), .B(n_0_2_28), .Z(n_0_2_299));
   XNOR2_X1 i_0_2_296 (.A(n_0_2_323), .B(n_0_2_301), .ZN(n_0_2_300));
   XNOR2_X1 i_0_2_297 (.A(n_0_2_1403), .B(n_0_2_27), .ZN(n_0_2_301));
   XNOR2_X1 i_0_2_298 (.A(n_0_2_26), .B(n_0_2_303), .ZN(n_0_2_302));
   XOR2_X1 i_0_2_299 (.A(n_0_2_1400), .B(n_0_2_326), .Z(n_0_2_303));
   XNOR2_X1 i_0_2_300 (.A(n_0_2_748), .B(n_0_2_327), .ZN(n_0_2_304));
   MUX2_X1 i_0_2_301 (.A(quotient[2]), .B(n_0_24), .S(n_0_2_847), .Z(n_0_43));
   MUX2_X1 i_0_2_302 (.A(quotient[3]), .B(n_0_25), .S(n_0_2_847), .Z(n_0_44));
   MUX2_X1 i_0_2_303 (.A(quotient[4]), .B(n_0_26), .S(n_0_2_847), .Z(n_0_45));
   MUX2_X1 i_0_2_304 (.A(quotient[5]), .B(n_0_27), .S(n_0_2_847), .Z(n_0_46));
   NOR2_X1 i_0_2_305 (.A1(n_0_2_24), .A2(n_0_2_50), .ZN(n_0_2_305));
   NAND2_X1 i_0_2_306 (.A1(n_0_2_24), .A2(n_0_2_50), .ZN(n_0_2_306));
   XNOR2_X1 i_0_2_307 (.A(n_0_2_490), .B(n_0_2_307), .ZN(n_0_2_24));
   NAND2_X1 i_0_2_308 (.A1(n_0_2_376), .A2(n_0_2_308), .ZN(n_0_2_307));
   XNOR2_X1 i_0_2_309 (.A(n_0_2_1439), .B(n_0_2_379), .ZN(n_0_2_308));
   NOR2_X1 i_0_2_310 (.A1(n_0_2_43), .A2(n_0_2_55), .ZN(n_0_2_309));
   NOR2_X1 i_0_2_311 (.A1(n_0_2_41), .A2(n_0_2_52), .ZN(n_0_2_310));
   NOR2_X1 i_0_2_312 (.A1(n_0_2_39), .A2(n_0_2_1352), .ZN(n_0_2_311));
   NOR2_X1 i_0_2_313 (.A1(n_0_2_37), .A2(n_0_2_1044), .ZN(n_0_2_312));
   NOR2_X1 i_0_2_314 (.A1(n_0_2_35), .A2(n_0_2_780), .ZN(n_0_2_313));
   NOR2_X1 i_0_2_315 (.A1(n_0_2_33), .A2(n_0_2_458), .ZN(n_0_2_314));
   NOR2_X1 i_0_2_316 (.A1(n_0_2_31), .A2(n_0_2_363), .ZN(n_0_2_315));
   AOI21_X1 i_0_2_317 (.A(n_0_2_317), .B1(n_0_2_318), .B2(n_0_2_335), .ZN(
      n_0_2_316));
   NOR2_X1 i_0_2_318 (.A1(n_0_2_29), .A2(n_0_2_209), .ZN(n_0_2_317));
   AOI21_X1 i_0_2_319 (.A(n_0_2_319), .B1(n_0_2_28), .B2(n_0_2_147), .ZN(
      n_0_2_318));
   INV_X1 i_0_2_320 (.A(n_0_2_320), .ZN(n_0_2_319));
   OAI21_X1 i_0_2_321 (.A(n_0_2_321), .B1(n_0_2_28), .B2(n_0_2_147), .ZN(
      n_0_2_320));
   AOI21_X1 i_0_2_322 (.A(n_0_2_322), .B1(n_0_2_323), .B2(n_0_2_330), .ZN(
      n_0_2_321));
   NOR2_X1 i_0_2_323 (.A1(n_0_2_27), .A2(n_0_2_96), .ZN(n_0_2_322));
   OAI21_X1 i_0_2_324 (.A(n_0_2_324), .B1(n_0_2_26), .B2(n_0_2_54), .ZN(
      n_0_2_323));
   INV_X1 i_0_2_325 (.A(n_0_2_325), .ZN(n_0_2_324));
   AOI21_X1 i_0_2_326 (.A(n_0_2_326), .B1(n_0_2_26), .B2(n_0_2_54), .ZN(
      n_0_2_325));
   OAI21_X1 i_0_2_327 (.A(n_0_2_1412), .B1(n_0_2_327), .B2(n_0_2_1366), .ZN(
      n_0_2_326));
   INV_X1 i_0_2_328 (.A(n_0_2_327), .ZN(n_0_2_25));
   NAND2_X1 i_0_2_329 (.A1(in_b[0]), .A2(n_0_2_376), .ZN(n_0_2_327));
   XOR2_X1 i_0_2_330 (.A(n_0_2_329), .B(n_0_2_328), .Z(n_0_2_26));
   NAND2_X1 i_0_2_331 (.A1(n_0_2_376), .A2(n_0_2_748), .ZN(n_0_2_328));
   NAND2_X1 i_0_2_332 (.A1(in_b[0]), .A2(n_0_2_494), .ZN(n_0_2_329));
   NAND2_X1 i_0_2_333 (.A1(n_0_2_27), .A2(n_0_2_96), .ZN(n_0_2_330));
   XNOR2_X1 i_0_2_334 (.A(n_0_2_424), .B(n_0_2_331), .ZN(n_0_2_27));
   NAND2_X1 i_0_2_335 (.A1(n_0_2_376), .A2(n_0_2_332), .ZN(n_0_2_331));
   XNOR2_X1 i_0_2_336 (.A(n_0_2_1400), .B(n_0_2_427), .ZN(n_0_2_332));
   XNOR2_X1 i_0_2_337 (.A(n_0_2_429), .B(n_0_2_333), .ZN(n_0_2_28));
   NAND2_X1 i_0_2_338 (.A1(n_0_2_376), .A2(n_0_2_334), .ZN(n_0_2_333));
   XOR2_X1 i_0_2_339 (.A(n_0_2_1403), .B(n_0_2_421), .Z(n_0_2_334));
   NAND2_X1 i_0_2_340 (.A1(n_0_2_29), .A2(n_0_2_209), .ZN(n_0_2_335));
   XNOR2_X1 i_0_2_341 (.A(n_0_2_432), .B(n_0_2_336), .ZN(n_0_2_29));
   NAND2_X1 i_0_2_342 (.A1(n_0_2_376), .A2(n_0_2_337), .ZN(n_0_2_336));
   XNOR2_X1 i_0_2_343 (.A(n_0_2_1406), .B(n_0_2_419), .ZN(n_0_2_337));
   XNOR2_X1 i_0_2_344 (.A(n_0_2_436), .B(n_0_2_338), .ZN(n_0_2_30));
   NAND2_X1 i_0_2_345 (.A1(n_0_2_376), .A2(n_0_2_339), .ZN(n_0_2_338));
   XOR2_X1 i_0_2_346 (.A(n_0_2_1408), .B(n_0_2_416), .Z(n_0_2_339));
   NAND2_X1 i_0_2_347 (.A1(n_0_2_31), .A2(n_0_2_363), .ZN(n_0_2_340));
   XNOR2_X1 i_0_2_348 (.A(n_0_2_439), .B(n_0_2_341), .ZN(n_0_2_31));
   NAND2_X1 i_0_2_349 (.A1(n_0_2_376), .A2(n_0_2_342), .ZN(n_0_2_341));
   XNOR2_X1 i_0_2_350 (.A(n_0_2_1410), .B(n_0_2_414), .ZN(n_0_2_342));
   XNOR2_X1 i_0_2_351 (.A(n_0_2_443), .B(n_0_2_343), .ZN(n_0_2_32));
   NAND2_X1 i_0_2_352 (.A1(n_0_2_376), .A2(n_0_2_344), .ZN(n_0_2_343));
   XOR2_X1 i_0_2_353 (.A(n_0_2_1413), .B(n_0_2_411), .Z(n_0_2_344));
   NAND2_X1 i_0_2_354 (.A1(n_0_2_33), .A2(n_0_2_458), .ZN(n_0_2_345));
   XNOR2_X1 i_0_2_355 (.A(n_0_2_446), .B(n_0_2_346), .ZN(n_0_2_33));
   NAND2_X1 i_0_2_356 (.A1(n_0_2_376), .A2(n_0_2_347), .ZN(n_0_2_346));
   XNOR2_X1 i_0_2_357 (.A(n_0_2_1415), .B(n_0_2_409), .ZN(n_0_2_347));
   XNOR2_X1 i_0_2_358 (.A(n_0_2_450), .B(n_0_2_348), .ZN(n_0_2_34));
   NAND2_X1 i_0_2_359 (.A1(n_0_2_376), .A2(n_0_2_349), .ZN(n_0_2_348));
   XOR2_X1 i_0_2_360 (.A(n_0_2_1417), .B(n_0_2_406), .Z(n_0_2_349));
   NAND2_X1 i_0_2_361 (.A1(n_0_2_35), .A2(n_0_2_780), .ZN(n_0_2_350));
   XNOR2_X1 i_0_2_362 (.A(n_0_2_454), .B(n_0_2_351), .ZN(n_0_2_35));
   NAND2_X1 i_0_2_363 (.A1(n_0_2_376), .A2(n_0_2_352), .ZN(n_0_2_351));
   XNOR2_X1 i_0_2_364 (.A(n_0_2_1418), .B(n_0_2_404), .ZN(n_0_2_352));
   XNOR2_X1 i_0_2_365 (.A(n_0_2_459), .B(n_0_2_353), .ZN(n_0_2_36));
   NAND2_X1 i_0_2_366 (.A1(n_0_2_376), .A2(n_0_2_354), .ZN(n_0_2_353));
   XOR2_X1 i_0_2_367 (.A(n_0_2_1440), .B(n_0_2_401), .Z(n_0_2_354));
   NAND2_X1 i_0_2_368 (.A1(n_0_2_37), .A2(n_0_2_1044), .ZN(n_0_2_355));
   XNOR2_X1 i_0_2_369 (.A(n_0_2_462), .B(n_0_2_356), .ZN(n_0_2_37));
   NAND2_X1 i_0_2_370 (.A1(n_0_2_376), .A2(n_0_2_357), .ZN(n_0_2_356));
   XNOR2_X1 i_0_2_371 (.A(n_0_2_1421), .B(n_0_2_399), .ZN(n_0_2_357));
   XNOR2_X1 i_0_2_372 (.A(n_0_2_466), .B(n_0_2_358), .ZN(n_0_2_38));
   NAND2_X1 i_0_2_373 (.A1(n_0_2_376), .A2(n_0_2_359), .ZN(n_0_2_358));
   XOR2_X1 i_0_2_374 (.A(n_0_2_1424), .B(n_0_2_396), .Z(n_0_2_359));
   NAND2_X1 i_0_2_375 (.A1(n_0_2_39), .A2(n_0_2_1352), .ZN(n_0_2_360));
   XNOR2_X1 i_0_2_376 (.A(n_0_2_469), .B(n_0_2_361), .ZN(n_0_2_39));
   NAND2_X1 i_0_2_377 (.A1(n_0_2_376), .A2(n_0_2_362), .ZN(n_0_2_361));
   XNOR2_X1 i_0_2_378 (.A(n_0_2_1429), .B(n_0_2_394), .ZN(n_0_2_362));
   XNOR2_X1 i_0_2_379 (.A(n_0_2_473), .B(n_0_2_364), .ZN(n_0_2_40));
   NAND2_X1 i_0_2_380 (.A1(n_0_2_376), .A2(n_0_2_365), .ZN(n_0_2_364));
   XOR2_X1 i_0_2_381 (.A(n_0_2_1427), .B(n_0_2_391), .Z(n_0_2_365));
   NAND2_X1 i_0_2_382 (.A1(n_0_2_41), .A2(n_0_2_52), .ZN(n_0_2_366));
   XNOR2_X1 i_0_2_383 (.A(n_0_2_476), .B(n_0_2_367), .ZN(n_0_2_41));
   NAND2_X1 i_0_2_384 (.A1(n_0_2_376), .A2(n_0_2_368), .ZN(n_0_2_367));
   XNOR2_X1 i_0_2_385 (.A(n_0_2_1428), .B(n_0_2_389), .ZN(n_0_2_368));
   XNOR2_X1 i_0_2_386 (.A(n_0_2_480), .B(n_0_2_369), .ZN(n_0_2_42));
   NAND2_X1 i_0_2_387 (.A1(n_0_2_376), .A2(n_0_2_370), .ZN(n_0_2_369));
   XOR2_X1 i_0_2_388 (.A(n_0_2_1434), .B(n_0_2_386), .Z(n_0_2_370));
   NAND2_X1 i_0_2_389 (.A1(n_0_2_43), .A2(n_0_2_55), .ZN(n_0_2_371));
   XNOR2_X1 i_0_2_390 (.A(n_0_2_483), .B(n_0_2_372), .ZN(n_0_2_43));
   NAND2_X1 i_0_2_391 (.A1(n_0_2_376), .A2(n_0_2_373), .ZN(n_0_2_372));
   XNOR2_X1 i_0_2_392 (.A(n_0_2_1436), .B(n_0_2_384), .ZN(n_0_2_373));
   XNOR2_X1 i_0_2_393 (.A(n_0_2_487), .B(n_0_2_374), .ZN(n_0_2_44));
   NAND2_X1 i_0_2_394 (.A1(n_0_2_376), .A2(n_0_2_375), .ZN(n_0_2_374));
   XOR2_X1 i_0_2_395 (.A(n_0_2_1438), .B(n_0_2_381), .Z(n_0_2_375));
   AND2_X1 i_0_2_396 (.A1(n_0_2_1394), .A2(n_0_2_376), .ZN(quotient[2]));
   NOR4_X1 i_0_2_397 (.A1(n_0_2_1432), .A2(n_0_2_1433), .A3(n_0_2_378), .A4(
      n_0_2_377), .ZN(n_0_2_376));
   NOR2_X1 i_0_2_398 (.A1(n_0_2_490), .A2(n_0_2_56), .ZN(n_0_2_377));
   AOI21_X1 i_0_2_399 (.A(n_0_2_379), .B1(n_0_2_490), .B2(n_0_2_56), .ZN(
      n_0_2_378));
   AOI21_X1 i_0_2_400 (.A(n_0_2_380), .B1(n_0_2_381), .B2(n_0_2_486), .ZN(
      n_0_2_379));
   NOR2_X1 i_0_2_401 (.A1(n_0_2_487), .A2(n_0_2_55), .ZN(n_0_2_380));
   AOI21_X1 i_0_2_402 (.A(n_0_2_382), .B1(n_0_2_483), .B2(n_0_2_53), .ZN(
      n_0_2_381));
   INV_X1 i_0_2_403 (.A(n_0_2_383), .ZN(n_0_2_382));
   OAI21_X1 i_0_2_404 (.A(n_0_2_384), .B1(n_0_2_483), .B2(n_0_2_53), .ZN(
      n_0_2_383));
   AOI21_X1 i_0_2_405 (.A(n_0_2_385), .B1(n_0_2_386), .B2(n_0_2_479), .ZN(
      n_0_2_384));
   NOR2_X1 i_0_2_406 (.A1(n_0_2_480), .A2(n_0_2_52), .ZN(n_0_2_385));
   AOI21_X1 i_0_2_407 (.A(n_0_2_387), .B1(n_0_2_476), .B2(n_0_2_1516), .ZN(
      n_0_2_386));
   INV_X1 i_0_2_408 (.A(n_0_2_388), .ZN(n_0_2_387));
   OAI21_X1 i_0_2_409 (.A(n_0_2_389), .B1(n_0_2_476), .B2(n_0_2_1516), .ZN(
      n_0_2_388));
   AOI21_X1 i_0_2_410 (.A(n_0_2_390), .B1(n_0_2_391), .B2(n_0_2_472), .ZN(
      n_0_2_389));
   NOR2_X1 i_0_2_411 (.A1(n_0_2_473), .A2(n_0_2_1352), .ZN(n_0_2_390));
   AOI21_X1 i_0_2_412 (.A(n_0_2_392), .B1(n_0_2_469), .B2(n_0_2_1190), .ZN(
      n_0_2_391));
   INV_X1 i_0_2_413 (.A(n_0_2_393), .ZN(n_0_2_392));
   OAI21_X1 i_0_2_414 (.A(n_0_2_394), .B1(n_0_2_469), .B2(n_0_2_1190), .ZN(
      n_0_2_393));
   AOI21_X1 i_0_2_415 (.A(n_0_2_395), .B1(n_0_2_396), .B2(n_0_2_465), .ZN(
      n_0_2_394));
   NOR2_X1 i_0_2_416 (.A1(n_0_2_466), .A2(n_0_2_1044), .ZN(n_0_2_395));
   AOI21_X1 i_0_2_417 (.A(n_0_2_397), .B1(n_0_2_462), .B2(n_0_2_907), .ZN(
      n_0_2_396));
   INV_X1 i_0_2_418 (.A(n_0_2_398), .ZN(n_0_2_397));
   OAI21_X1 i_0_2_419 (.A(n_0_2_399), .B1(n_0_2_462), .B2(n_0_2_907), .ZN(
      n_0_2_398));
   AOI21_X1 i_0_2_420 (.A(n_0_2_400), .B1(n_0_2_401), .B2(n_0_2_457), .ZN(
      n_0_2_399));
   NOR2_X1 i_0_2_421 (.A1(n_0_2_459), .A2(n_0_2_780), .ZN(n_0_2_400));
   AOI21_X1 i_0_2_422 (.A(n_0_2_402), .B1(n_0_2_454), .B2(n_0_2_660), .ZN(
      n_0_2_401));
   INV_X1 i_0_2_423 (.A(n_0_2_403), .ZN(n_0_2_402));
   OAI21_X1 i_0_2_424 (.A(n_0_2_404), .B1(n_0_2_454), .B2(n_0_2_660), .ZN(
      n_0_2_403));
   AOI21_X1 i_0_2_425 (.A(n_0_2_405), .B1(n_0_2_406), .B2(n_0_2_449), .ZN(
      n_0_2_404));
   NOR2_X1 i_0_2_426 (.A1(n_0_2_450), .A2(n_0_2_458), .ZN(n_0_2_405));
   AOI21_X1 i_0_2_427 (.A(n_0_2_407), .B1(n_0_2_446), .B2(n_0_2_453), .ZN(
      n_0_2_406));
   INV_X1 i_0_2_428 (.A(n_0_2_408), .ZN(n_0_2_407));
   OAI21_X1 i_0_2_429 (.A(n_0_2_409), .B1(n_0_2_446), .B2(n_0_2_453), .ZN(
      n_0_2_408));
   AOI21_X1 i_0_2_430 (.A(n_0_2_410), .B1(n_0_2_411), .B2(n_0_2_442), .ZN(
      n_0_2_409));
   NOR2_X1 i_0_2_431 (.A1(n_0_2_443), .A2(n_0_2_363), .ZN(n_0_2_410));
   AOI21_X1 i_0_2_432 (.A(n_0_2_412), .B1(n_0_2_439), .B2(n_0_2_281), .ZN(
      n_0_2_411));
   INV_X1 i_0_2_433 (.A(n_0_2_413), .ZN(n_0_2_412));
   OAI21_X1 i_0_2_434 (.A(n_0_2_414), .B1(n_0_2_439), .B2(n_0_2_281), .ZN(
      n_0_2_413));
   AOI21_X1 i_0_2_435 (.A(n_0_2_415), .B1(n_0_2_416), .B2(n_0_2_435), .ZN(
      n_0_2_414));
   NOR2_X1 i_0_2_436 (.A1(n_0_2_436), .A2(n_0_2_209), .ZN(n_0_2_415));
   AOI21_X1 i_0_2_437 (.A(n_0_2_417), .B1(n_0_2_432), .B2(n_0_2_147), .ZN(
      n_0_2_416));
   INV_X1 i_0_2_438 (.A(n_0_2_418), .ZN(n_0_2_417));
   OAI21_X1 i_0_2_439 (.A(n_0_2_419), .B1(n_0_2_432), .B2(n_0_2_147), .ZN(
      n_0_2_418));
   AOI21_X1 i_0_2_440 (.A(n_0_2_420), .B1(n_0_2_421), .B2(n_0_2_428), .ZN(
      n_0_2_419));
   NOR2_X1 i_0_2_441 (.A1(n_0_2_429), .A2(n_0_2_96), .ZN(n_0_2_420));
   AOI21_X1 i_0_2_442 (.A(n_0_2_422), .B1(n_0_2_427), .B2(n_0_2_54), .ZN(
      n_0_2_421));
   INV_X1 i_0_2_443 (.A(n_0_2_423), .ZN(n_0_2_422));
   OAI21_X1 i_0_2_444 (.A(n_0_2_424), .B1(n_0_2_427), .B2(n_0_2_54), .ZN(
      n_0_2_423));
   XOR2_X1 i_0_2_445 (.A(n_0_2_426), .B(n_0_2_425), .Z(n_0_2_424));
   NAND2_X1 i_0_2_446 (.A1(n_0_2_494), .A2(n_0_2_748), .ZN(n_0_2_425));
   NAND2_X1 i_0_2_447 (.A1(in_b[0]), .A2(n_0_2_615), .ZN(n_0_2_426));
   OAI21_X1 i_0_2_448 (.A(n_0_2_1412), .B1(n_0_2_745), .B2(n_0_2_493), .ZN(
      n_0_2_427));
   NAND2_X1 i_0_2_449 (.A1(n_0_2_429), .A2(n_0_2_96), .ZN(n_0_2_428));
   XOR2_X1 i_0_2_450 (.A(n_0_2_540), .B(n_0_2_430), .Z(n_0_2_429));
   NAND2_X1 i_0_2_451 (.A1(n_0_2_494), .A2(n_0_2_431), .ZN(n_0_2_430));
   XNOR2_X1 i_0_2_452 (.A(n_0_2_1400), .B(n_0_2_539), .ZN(n_0_2_431));
   XNOR2_X1 i_0_2_453 (.A(n_0_2_545), .B(n_0_2_433), .ZN(n_0_2_432));
   NAND2_X1 i_0_2_454 (.A1(n_0_2_494), .A2(n_0_2_434), .ZN(n_0_2_433));
   XOR2_X1 i_0_2_455 (.A(n_0_2_1403), .B(n_0_2_536), .Z(n_0_2_434));
   NAND2_X1 i_0_2_456 (.A1(n_0_2_436), .A2(n_0_2_209), .ZN(n_0_2_435));
   XOR2_X1 i_0_2_457 (.A(n_0_2_549), .B(n_0_2_437), .Z(n_0_2_436));
   NAND2_X1 i_0_2_458 (.A1(n_0_2_494), .A2(n_0_2_438), .ZN(n_0_2_437));
   XNOR2_X1 i_0_2_459 (.A(n_0_2_1406), .B(n_0_2_534), .ZN(n_0_2_438));
   XNOR2_X1 i_0_2_460 (.A(n_0_2_553), .B(n_0_2_440), .ZN(n_0_2_439));
   NAND2_X1 i_0_2_461 (.A1(n_0_2_494), .A2(n_0_2_441), .ZN(n_0_2_440));
   XOR2_X1 i_0_2_462 (.A(n_0_2_1408), .B(n_0_2_531), .Z(n_0_2_441));
   NAND2_X1 i_0_2_463 (.A1(n_0_2_443), .A2(n_0_2_363), .ZN(n_0_2_442));
   XOR2_X1 i_0_2_464 (.A(n_0_2_557), .B(n_0_2_444), .Z(n_0_2_443));
   NAND2_X1 i_0_2_465 (.A1(n_0_2_494), .A2(n_0_2_445), .ZN(n_0_2_444));
   XNOR2_X1 i_0_2_466 (.A(n_0_2_1410), .B(n_0_2_529), .ZN(n_0_2_445));
   XNOR2_X1 i_0_2_467 (.A(n_0_2_561), .B(n_0_2_447), .ZN(n_0_2_446));
   NAND2_X1 i_0_2_468 (.A1(n_0_2_494), .A2(n_0_2_448), .ZN(n_0_2_447));
   XOR2_X1 i_0_2_469 (.A(n_0_2_1413), .B(n_0_2_526), .Z(n_0_2_448));
   NAND2_X1 i_0_2_470 (.A1(n_0_2_450), .A2(n_0_2_458), .ZN(n_0_2_449));
   XOR2_X1 i_0_2_471 (.A(n_0_2_566), .B(n_0_2_451), .Z(n_0_2_450));
   NAND2_X1 i_0_2_472 (.A1(n_0_2_494), .A2(n_0_2_452), .ZN(n_0_2_451));
   XNOR2_X1 i_0_2_473 (.A(n_0_2_1415), .B(n_0_2_524), .ZN(n_0_2_452));
   XNOR2_X1 i_0_2_474 (.A(n_0_2_570), .B(n_0_2_455), .ZN(n_0_2_454));
   NAND2_X1 i_0_2_475 (.A1(n_0_2_494), .A2(n_0_2_456), .ZN(n_0_2_455));
   XOR2_X1 i_0_2_476 (.A(n_0_2_1417), .B(n_0_2_522), .Z(n_0_2_456));
   NAND2_X1 i_0_2_477 (.A1(n_0_2_459), .A2(n_0_2_780), .ZN(n_0_2_457));
   XOR2_X1 i_0_2_478 (.A(n_0_2_575), .B(n_0_2_460), .Z(n_0_2_459));
   NAND2_X1 i_0_2_479 (.A1(n_0_2_494), .A2(n_0_2_461), .ZN(n_0_2_460));
   XNOR2_X1 i_0_2_480 (.A(n_0_2_1418), .B(n_0_2_520), .ZN(n_0_2_461));
   XNOR2_X1 i_0_2_481 (.A(n_0_2_579), .B(n_0_2_463), .ZN(n_0_2_462));
   NAND2_X1 i_0_2_482 (.A1(n_0_2_494), .A2(n_0_2_464), .ZN(n_0_2_463));
   XOR2_X1 i_0_2_483 (.A(n_0_2_1440), .B(n_0_2_518), .Z(n_0_2_464));
   NAND2_X1 i_0_2_484 (.A1(n_0_2_466), .A2(n_0_2_1044), .ZN(n_0_2_465));
   XOR2_X1 i_0_2_485 (.A(n_0_2_584), .B(n_0_2_467), .Z(n_0_2_466));
   NAND2_X1 i_0_2_486 (.A1(n_0_2_494), .A2(n_0_2_468), .ZN(n_0_2_467));
   XNOR2_X1 i_0_2_487 (.A(n_0_2_1421), .B(n_0_2_516), .ZN(n_0_2_468));
   XNOR2_X1 i_0_2_488 (.A(n_0_2_588), .B(n_0_2_470), .ZN(n_0_2_469));
   NAND2_X1 i_0_2_489 (.A1(n_0_2_494), .A2(n_0_2_471), .ZN(n_0_2_470));
   XOR2_X1 i_0_2_490 (.A(n_0_2_1424), .B(n_0_2_514), .Z(n_0_2_471));
   NAND2_X1 i_0_2_491 (.A1(n_0_2_473), .A2(n_0_2_1352), .ZN(n_0_2_472));
   XOR2_X1 i_0_2_492 (.A(n_0_2_593), .B(n_0_2_474), .Z(n_0_2_473));
   NAND2_X1 i_0_2_493 (.A1(n_0_2_494), .A2(n_0_2_475), .ZN(n_0_2_474));
   XNOR2_X1 i_0_2_494 (.A(n_0_2_1429), .B(n_0_2_512), .ZN(n_0_2_475));
   XNOR2_X1 i_0_2_495 (.A(n_0_2_597), .B(n_0_2_477), .ZN(n_0_2_476));
   NAND2_X1 i_0_2_496 (.A1(n_0_2_494), .A2(n_0_2_478), .ZN(n_0_2_477));
   XOR2_X1 i_0_2_497 (.A(n_0_2_1427), .B(n_0_2_510), .Z(n_0_2_478));
   NAND2_X1 i_0_2_498 (.A1(n_0_2_480), .A2(n_0_2_52), .ZN(n_0_2_479));
   XOR2_X1 i_0_2_499 (.A(n_0_2_601), .B(n_0_2_481), .Z(n_0_2_480));
   NAND2_X1 i_0_2_500 (.A1(n_0_2_494), .A2(n_0_2_482), .ZN(n_0_2_481));
   XNOR2_X1 i_0_2_501 (.A(n_0_2_1428), .B(n_0_2_508), .ZN(n_0_2_482));
   XNOR2_X1 i_0_2_502 (.A(n_0_2_605), .B(n_0_2_484), .ZN(n_0_2_483));
   NAND2_X1 i_0_2_503 (.A1(n_0_2_494), .A2(n_0_2_485), .ZN(n_0_2_484));
   XOR2_X1 i_0_2_504 (.A(n_0_2_1434), .B(n_0_2_505), .Z(n_0_2_485));
   NAND2_X1 i_0_2_505 (.A1(n_0_2_487), .A2(n_0_2_55), .ZN(n_0_2_486));
   XOR2_X1 i_0_2_506 (.A(n_0_2_610), .B(n_0_2_488), .Z(n_0_2_487));
   NAND2_X1 i_0_2_507 (.A1(n_0_2_494), .A2(n_0_2_489), .ZN(n_0_2_488));
   XNOR2_X1 i_0_2_508 (.A(n_0_2_1436), .B(n_0_2_503), .ZN(n_0_2_489));
   XNOR2_X1 i_0_2_509 (.A(n_0_2_497), .B(n_0_2_491), .ZN(n_0_2_490));
   NAND2_X1 i_0_2_510 (.A1(n_0_2_494), .A2(n_0_2_492), .ZN(n_0_2_491));
   XOR2_X1 i_0_2_511 (.A(n_0_2_1438), .B(n_0_2_501), .Z(n_0_2_492));
   NOR2_X1 i_0_2_512 (.A1(n_0_2_1395), .A2(n_0_2_493), .ZN(quotient[3]));
   INV_X1 i_0_2_513 (.A(n_0_2_494), .ZN(n_0_2_493));
   AOI21_X1 i_0_2_514 (.A(n_0_2_495), .B1(n_0_2_496), .B2(n_0_2_501), .ZN(
      n_0_2_494));
   OAI21_X1 i_0_2_515 (.A(n_0_2_744), .B1(n_0_2_497), .B2(n_0_2_55), .ZN(
      n_0_2_495));
   NAND2_X1 i_0_2_516 (.A1(n_0_2_497), .A2(n_0_2_55), .ZN(n_0_2_496));
   INV_X1 i_0_2_517 (.A(n_0_2_498), .ZN(n_0_2_497));
   AOI22_X1 i_0_2_518 (.A1(n_0_2_615), .A2(n_0_2_499), .B1(n_0_2_613), .B2(
      n_0_2_701), .ZN(n_0_2_498));
   XNOR2_X1 i_0_2_519 (.A(n_0_2_620), .B(n_0_2_500), .ZN(n_0_2_499));
   XNOR2_X1 i_0_2_520 (.A(n_0_2_1436), .B(n_0_2_700), .ZN(n_0_2_500));
   AOI21_X1 i_0_2_521 (.A(n_0_2_502), .B1(n_0_2_503), .B2(n_0_2_609), .ZN(
      n_0_2_501));
   NOR2_X1 i_0_2_522 (.A1(n_0_2_610), .A2(n_0_2_1436), .ZN(n_0_2_502));
   OAI21_X1 i_0_2_523 (.A(n_0_2_504), .B1(n_0_2_505), .B2(n_0_2_604), .ZN(
      n_0_2_503));
   NAND2_X1 i_0_2_524 (.A1(n_0_2_605), .A2(n_0_2_52), .ZN(n_0_2_504));
   AOI21_X1 i_0_2_525 (.A(n_0_2_506), .B1(n_0_2_508), .B2(n_0_2_1516), .ZN(
      n_0_2_505));
   NOR2_X1 i_0_2_526 (.A1(n_0_2_601), .A2(n_0_2_507), .ZN(n_0_2_506));
   NOR2_X1 i_0_2_527 (.A1(n_0_2_1516), .A2(n_0_2_508), .ZN(n_0_2_507));
   OAI21_X1 i_0_2_528 (.A(n_0_2_509), .B1(n_0_2_510), .B2(n_0_2_596), .ZN(
      n_0_2_508));
   NAND2_X1 i_0_2_529 (.A1(n_0_2_597), .A2(n_0_2_1352), .ZN(n_0_2_509));
   AOI21_X1 i_0_2_530 (.A(n_0_2_511), .B1(n_0_2_512), .B2(n_0_2_592), .ZN(
      n_0_2_510));
   NOR2_X1 i_0_2_531 (.A1(n_0_2_593), .A2(n_0_2_1429), .ZN(n_0_2_511));
   OAI21_X1 i_0_2_532 (.A(n_0_2_513), .B1(n_0_2_514), .B2(n_0_2_587), .ZN(
      n_0_2_512));
   NAND2_X1 i_0_2_533 (.A1(n_0_2_588), .A2(n_0_2_1044), .ZN(n_0_2_513));
   AOI21_X1 i_0_2_534 (.A(n_0_2_515), .B1(n_0_2_516), .B2(n_0_2_583), .ZN(
      n_0_2_514));
   NOR2_X1 i_0_2_535 (.A1(n_0_2_584), .A2(n_0_2_1421), .ZN(n_0_2_515));
   OAI21_X1 i_0_2_536 (.A(n_0_2_517), .B1(n_0_2_518), .B2(n_0_2_578), .ZN(
      n_0_2_516));
   NAND2_X1 i_0_2_537 (.A1(n_0_2_579), .A2(n_0_2_780), .ZN(n_0_2_517));
   AOI21_X1 i_0_2_538 (.A(n_0_2_519), .B1(n_0_2_520), .B2(n_0_2_574), .ZN(
      n_0_2_518));
   NOR2_X1 i_0_2_539 (.A1(n_0_2_575), .A2(n_0_2_1418), .ZN(n_0_2_519));
   OAI21_X1 i_0_2_540 (.A(n_0_2_521), .B1(n_0_2_522), .B2(n_0_2_569), .ZN(
      n_0_2_520));
   NAND2_X1 i_0_2_541 (.A1(n_0_2_570), .A2(n_0_2_458), .ZN(n_0_2_521));
   AOI21_X1 i_0_2_542 (.A(n_0_2_523), .B1(n_0_2_524), .B2(n_0_2_565), .ZN(
      n_0_2_522));
   NOR2_X1 i_0_2_543 (.A1(n_0_2_566), .A2(n_0_2_1415), .ZN(n_0_2_523));
   OAI21_X1 i_0_2_544 (.A(n_0_2_525), .B1(n_0_2_526), .B2(n_0_2_560), .ZN(
      n_0_2_524));
   NAND2_X1 i_0_2_545 (.A1(n_0_2_561), .A2(n_0_2_363), .ZN(n_0_2_525));
   AOI21_X1 i_0_2_546 (.A(n_0_2_527), .B1(n_0_2_529), .B2(n_0_2_281), .ZN(
      n_0_2_526));
   NOR2_X1 i_0_2_547 (.A1(n_0_2_557), .A2(n_0_2_528), .ZN(n_0_2_527));
   NOR2_X1 i_0_2_548 (.A1(n_0_2_281), .A2(n_0_2_529), .ZN(n_0_2_528));
   OAI21_X1 i_0_2_549 (.A(n_0_2_530), .B1(n_0_2_531), .B2(n_0_2_552), .ZN(
      n_0_2_529));
   NAND2_X1 i_0_2_550 (.A1(n_0_2_553), .A2(n_0_2_209), .ZN(n_0_2_530));
   AOI21_X1 i_0_2_551 (.A(n_0_2_532), .B1(n_0_2_534), .B2(n_0_2_147), .ZN(
      n_0_2_531));
   NOR2_X1 i_0_2_552 (.A1(n_0_2_549), .A2(n_0_2_533), .ZN(n_0_2_532));
   NOR2_X1 i_0_2_553 (.A1(n_0_2_147), .A2(n_0_2_534), .ZN(n_0_2_533));
   OAI21_X1 i_0_2_554 (.A(n_0_2_535), .B1(n_0_2_536), .B2(n_0_2_544), .ZN(
      n_0_2_534));
   NAND2_X1 i_0_2_555 (.A1(n_0_2_545), .A2(n_0_2_96), .ZN(n_0_2_535));
   AOI21_X1 i_0_2_556 (.A(n_0_2_537), .B1(n_0_2_539), .B2(n_0_2_54), .ZN(
      n_0_2_536));
   NOR2_X1 i_0_2_557 (.A1(n_0_2_540), .A2(n_0_2_538), .ZN(n_0_2_537));
   NOR2_X1 i_0_2_558 (.A1(n_0_2_539), .A2(n_0_2_54), .ZN(n_0_2_538));
   OAI21_X1 i_0_2_559 (.A(n_0_2_1412), .B1(n_0_2_745), .B2(n_0_2_614), .ZN(
      n_0_2_539));
   AOI22_X1 i_0_2_560 (.A1(n_0_2_542), .A2(n_0_2_613), .B1(n_0_2_615), .B2(
      n_0_2_541), .ZN(n_0_2_540));
   XNOR2_X1 i_0_2_561 (.A(n_0_2_543), .B(n_0_2_748), .ZN(n_0_2_541));
   INV_X1 i_0_2_562 (.A(n_0_2_543), .ZN(n_0_2_542));
   NAND2_X1 i_0_2_563 (.A1(in_b[0]), .A2(n_0_2_704), .ZN(n_0_2_543));
   NOR2_X1 i_0_2_564 (.A1(n_0_2_545), .A2(n_0_2_96), .ZN(n_0_2_544));
   INV_X1 i_0_2_565 (.A(n_0_2_546), .ZN(n_0_2_545));
   AOI22_X1 i_0_2_566 (.A1(n_0_2_615), .A2(n_0_2_547), .B1(n_0_2_613), .B2(
      n_0_2_661), .ZN(n_0_2_546));
   XNOR2_X1 i_0_2_567 (.A(n_0_2_661), .B(n_0_2_548), .ZN(n_0_2_547));
   XOR2_X1 i_0_2_568 (.A(n_0_2_1400), .B(n_0_2_662), .Z(n_0_2_548));
   AOI22_X1 i_0_2_569 (.A1(n_0_2_615), .A2(n_0_2_550), .B1(n_0_2_613), .B2(
      n_0_2_664), .ZN(n_0_2_549));
   XNOR2_X1 i_0_2_570 (.A(n_0_2_657), .B(n_0_2_551), .ZN(n_0_2_550));
   XNOR2_X1 i_0_2_571 (.A(n_0_2_1403), .B(n_0_2_664), .ZN(n_0_2_551));
   NOR2_X1 i_0_2_572 (.A1(n_0_2_553), .A2(n_0_2_209), .ZN(n_0_2_552));
   INV_X1 i_0_2_573 (.A(n_0_2_554), .ZN(n_0_2_553));
   AOI22_X1 i_0_2_574 (.A1(n_0_2_615), .A2(n_0_2_555), .B1(n_0_2_613), .B2(
      n_0_2_665), .ZN(n_0_2_554));
   XNOR2_X1 i_0_2_575 (.A(n_0_2_655), .B(n_0_2_556), .ZN(n_0_2_555));
   XOR2_X1 i_0_2_576 (.A(n_0_2_1406), .B(n_0_2_665), .Z(n_0_2_556));
   AOI22_X1 i_0_2_577 (.A1(n_0_2_615), .A2(n_0_2_558), .B1(n_0_2_613), .B2(
      n_0_2_668), .ZN(n_0_2_557));
   XNOR2_X1 i_0_2_578 (.A(n_0_2_652), .B(n_0_2_559), .ZN(n_0_2_558));
   XNOR2_X1 i_0_2_579 (.A(n_0_2_1408), .B(n_0_2_668), .ZN(n_0_2_559));
   NOR2_X1 i_0_2_580 (.A1(n_0_2_561), .A2(n_0_2_363), .ZN(n_0_2_560));
   INV_X1 i_0_2_581 (.A(n_0_2_562), .ZN(n_0_2_561));
   AOI22_X1 i_0_2_582 (.A1(n_0_2_615), .A2(n_0_2_563), .B1(n_0_2_613), .B2(
      n_0_2_670), .ZN(n_0_2_562));
   XNOR2_X1 i_0_2_583 (.A(n_0_2_650), .B(n_0_2_564), .ZN(n_0_2_563));
   XOR2_X1 i_0_2_584 (.A(n_0_2_1410), .B(n_0_2_670), .Z(n_0_2_564));
   NAND2_X1 i_0_2_585 (.A1(n_0_2_566), .A2(n_0_2_1415), .ZN(n_0_2_565));
   AOI22_X1 i_0_2_586 (.A1(n_0_2_615), .A2(n_0_2_567), .B1(n_0_2_613), .B2(
      n_0_2_673), .ZN(n_0_2_566));
   XNOR2_X1 i_0_2_587 (.A(n_0_2_647), .B(n_0_2_568), .ZN(n_0_2_567));
   XNOR2_X1 i_0_2_588 (.A(n_0_2_1413), .B(n_0_2_673), .ZN(n_0_2_568));
   NOR2_X1 i_0_2_589 (.A1(n_0_2_570), .A2(n_0_2_458), .ZN(n_0_2_569));
   INV_X1 i_0_2_590 (.A(n_0_2_571), .ZN(n_0_2_570));
   AOI22_X1 i_0_2_591 (.A1(n_0_2_615), .A2(n_0_2_572), .B1(n_0_2_613), .B2(
      n_0_2_675), .ZN(n_0_2_571));
   XNOR2_X1 i_0_2_592 (.A(n_0_2_645), .B(n_0_2_573), .ZN(n_0_2_572));
   XOR2_X1 i_0_2_593 (.A(n_0_2_1415), .B(n_0_2_675), .Z(n_0_2_573));
   NAND2_X1 i_0_2_594 (.A1(n_0_2_575), .A2(n_0_2_1418), .ZN(n_0_2_574));
   AOI22_X1 i_0_2_595 (.A1(n_0_2_615), .A2(n_0_2_576), .B1(n_0_2_613), .B2(
      n_0_2_678), .ZN(n_0_2_575));
   XNOR2_X1 i_0_2_596 (.A(n_0_2_642), .B(n_0_2_577), .ZN(n_0_2_576));
   XNOR2_X1 i_0_2_597 (.A(n_0_2_1417), .B(n_0_2_678), .ZN(n_0_2_577));
   NOR2_X1 i_0_2_598 (.A1(n_0_2_579), .A2(n_0_2_780), .ZN(n_0_2_578));
   INV_X1 i_0_2_599 (.A(n_0_2_580), .ZN(n_0_2_579));
   AOI22_X1 i_0_2_600 (.A1(n_0_2_680), .A2(n_0_2_613), .B1(n_0_2_615), .B2(
      n_0_2_581), .ZN(n_0_2_580));
   XNOR2_X1 i_0_2_601 (.A(n_0_2_640), .B(n_0_2_582), .ZN(n_0_2_581));
   XOR2_X1 i_0_2_602 (.A(n_0_2_1418), .B(n_0_2_680), .Z(n_0_2_582));
   NAND2_X1 i_0_2_603 (.A1(n_0_2_584), .A2(n_0_2_1421), .ZN(n_0_2_583));
   AOI22_X1 i_0_2_604 (.A1(n_0_2_683), .A2(n_0_2_613), .B1(n_0_2_615), .B2(
      n_0_2_585), .ZN(n_0_2_584));
   XNOR2_X1 i_0_2_605 (.A(n_0_2_637), .B(n_0_2_586), .ZN(n_0_2_585));
   XNOR2_X1 i_0_2_606 (.A(n_0_2_1440), .B(n_0_2_683), .ZN(n_0_2_586));
   NOR2_X1 i_0_2_607 (.A1(n_0_2_588), .A2(n_0_2_1044), .ZN(n_0_2_587));
   INV_X1 i_0_2_608 (.A(n_0_2_589), .ZN(n_0_2_588));
   AOI22_X1 i_0_2_609 (.A1(n_0_2_685), .A2(n_0_2_613), .B1(n_0_2_615), .B2(
      n_0_2_590), .ZN(n_0_2_589));
   XNOR2_X1 i_0_2_610 (.A(n_0_2_635), .B(n_0_2_591), .ZN(n_0_2_590));
   XOR2_X1 i_0_2_611 (.A(n_0_2_1421), .B(n_0_2_685), .Z(n_0_2_591));
   NAND2_X1 i_0_2_612 (.A1(n_0_2_593), .A2(n_0_2_1429), .ZN(n_0_2_592));
   AOI22_X1 i_0_2_613 (.A1(n_0_2_615), .A2(n_0_2_594), .B1(n_0_2_613), .B2(
      n_0_2_688), .ZN(n_0_2_593));
   XNOR2_X1 i_0_2_614 (.A(n_0_2_632), .B(n_0_2_595), .ZN(n_0_2_594));
   XNOR2_X1 i_0_2_615 (.A(n_0_2_1424), .B(n_0_2_688), .ZN(n_0_2_595));
   NOR2_X1 i_0_2_616 (.A1(n_0_2_597), .A2(n_0_2_1352), .ZN(n_0_2_596));
   INV_X1 i_0_2_617 (.A(n_0_2_598), .ZN(n_0_2_597));
   AOI22_X1 i_0_2_618 (.A1(n_0_2_690), .A2(n_0_2_613), .B1(n_0_2_615), .B2(
      n_0_2_599), .ZN(n_0_2_598));
   XNOR2_X1 i_0_2_619 (.A(n_0_2_630), .B(n_0_2_600), .ZN(n_0_2_599));
   XOR2_X1 i_0_2_620 (.A(n_0_2_1429), .B(n_0_2_690), .Z(n_0_2_600));
   AOI22_X1 i_0_2_621 (.A1(n_0_2_693), .A2(n_0_2_613), .B1(n_0_2_615), .B2(
      n_0_2_602), .ZN(n_0_2_601));
   XNOR2_X1 i_0_2_622 (.A(n_0_2_627), .B(n_0_2_603), .ZN(n_0_2_602));
   XNOR2_X1 i_0_2_623 (.A(n_0_2_1427), .B(n_0_2_693), .ZN(n_0_2_603));
   NOR2_X1 i_0_2_624 (.A1(n_0_2_605), .A2(n_0_2_52), .ZN(n_0_2_604));
   INV_X1 i_0_2_625 (.A(n_0_2_606), .ZN(n_0_2_605));
   AOI22_X1 i_0_2_626 (.A1(n_0_2_695), .A2(n_0_2_613), .B1(n_0_2_615), .B2(
      n_0_2_607), .ZN(n_0_2_606));
   XNOR2_X1 i_0_2_627 (.A(n_0_2_625), .B(n_0_2_608), .ZN(n_0_2_607));
   XOR2_X1 i_0_2_628 (.A(n_0_2_1428), .B(n_0_2_695), .Z(n_0_2_608));
   NAND2_X1 i_0_2_629 (.A1(n_0_2_610), .A2(n_0_2_1436), .ZN(n_0_2_609));
   AOI22_X1 i_0_2_630 (.A1(n_0_2_615), .A2(n_0_2_611), .B1(n_0_2_613), .B2(
      n_0_2_698), .ZN(n_0_2_610));
   XNOR2_X1 i_0_2_631 (.A(n_0_2_622), .B(n_0_2_612), .ZN(n_0_2_611));
   XNOR2_X1 i_0_2_632 (.A(n_0_2_1434), .B(n_0_2_698), .ZN(n_0_2_612));
   NAND2_X1 i_0_2_633 (.A1(n_0_2_46), .A2(n_0_2_616), .ZN(n_0_2_613));
   NOR2_X1 i_0_2_634 (.A1(n_0_2_1395), .A2(n_0_2_614), .ZN(quotient[4]));
   INV_X1 i_0_2_635 (.A(n_0_2_615), .ZN(n_0_2_614));
   NOR3_X1 i_0_2_636 (.A1(n_0_2_1432), .A2(n_0_2_47), .A3(n_0_2_617), .ZN(
      n_0_2_615));
   NOR2_X1 i_0_2_637 (.A1(n_0_2_1432), .A2(n_0_2_617), .ZN(n_0_2_616));
   XNOR2_X1 i_0_2_638 (.A(n_0_2_1438), .B(n_0_2_618), .ZN(n_0_2_617));
   OAI21_X1 i_0_2_639 (.A(n_0_2_619), .B1(n_0_2_700), .B2(n_0_2_1436), .ZN(
      n_0_2_618));
   OAI21_X1 i_0_2_640 (.A(n_0_2_620), .B1(n_0_2_701), .B2(n_0_2_53), .ZN(
      n_0_2_619));
   AOI21_X1 i_0_2_641 (.A(n_0_2_621), .B1(n_0_2_622), .B2(n_0_2_697), .ZN(
      n_0_2_620));
   NOR2_X1 i_0_2_642 (.A1(n_0_2_698), .A2(n_0_2_52), .ZN(n_0_2_621));
   AOI21_X1 i_0_2_643 (.A(n_0_2_623), .B1(n_0_2_695), .B2(n_0_2_1516), .ZN(
      n_0_2_622));
   INV_X1 i_0_2_644 (.A(n_0_2_624), .ZN(n_0_2_623));
   OAI21_X1 i_0_2_645 (.A(n_0_2_625), .B1(n_0_2_695), .B2(n_0_2_1516), .ZN(
      n_0_2_624));
   AOI21_X1 i_0_2_646 (.A(n_0_2_626), .B1(n_0_2_627), .B2(n_0_2_692), .ZN(
      n_0_2_625));
   NOR2_X1 i_0_2_647 (.A1(n_0_2_693), .A2(n_0_2_1352), .ZN(n_0_2_626));
   AOI21_X1 i_0_2_648 (.A(n_0_2_628), .B1(n_0_2_690), .B2(n_0_2_1190), .ZN(
      n_0_2_627));
   INV_X1 i_0_2_649 (.A(n_0_2_629), .ZN(n_0_2_628));
   OAI21_X1 i_0_2_650 (.A(n_0_2_630), .B1(n_0_2_690), .B2(n_0_2_1190), .ZN(
      n_0_2_629));
   AOI21_X1 i_0_2_651 (.A(n_0_2_631), .B1(n_0_2_632), .B2(n_0_2_687), .ZN(
      n_0_2_630));
   NOR2_X1 i_0_2_652 (.A1(n_0_2_688), .A2(n_0_2_1044), .ZN(n_0_2_631));
   AOI21_X1 i_0_2_653 (.A(n_0_2_633), .B1(n_0_2_685), .B2(n_0_2_907), .ZN(
      n_0_2_632));
   INV_X1 i_0_2_654 (.A(n_0_2_634), .ZN(n_0_2_633));
   OAI21_X1 i_0_2_655 (.A(n_0_2_635), .B1(n_0_2_685), .B2(n_0_2_907), .ZN(
      n_0_2_634));
   AOI21_X1 i_0_2_656 (.A(n_0_2_636), .B1(n_0_2_637), .B2(n_0_2_682), .ZN(
      n_0_2_635));
   NOR2_X1 i_0_2_657 (.A1(n_0_2_683), .A2(n_0_2_780), .ZN(n_0_2_636));
   AOI21_X1 i_0_2_658 (.A(n_0_2_638), .B1(n_0_2_680), .B2(n_0_2_660), .ZN(
      n_0_2_637));
   INV_X1 i_0_2_659 (.A(n_0_2_639), .ZN(n_0_2_638));
   OAI21_X1 i_0_2_660 (.A(n_0_2_640), .B1(n_0_2_680), .B2(n_0_2_660), .ZN(
      n_0_2_639));
   AOI21_X1 i_0_2_661 (.A(n_0_2_641), .B1(n_0_2_642), .B2(n_0_2_677), .ZN(
      n_0_2_640));
   NOR2_X1 i_0_2_662 (.A1(n_0_2_678), .A2(n_0_2_458), .ZN(n_0_2_641));
   AOI21_X1 i_0_2_663 (.A(n_0_2_643), .B1(n_0_2_675), .B2(n_0_2_453), .ZN(
      n_0_2_642));
   INV_X1 i_0_2_664 (.A(n_0_2_644), .ZN(n_0_2_643));
   OAI21_X1 i_0_2_665 (.A(n_0_2_645), .B1(n_0_2_675), .B2(n_0_2_453), .ZN(
      n_0_2_644));
   AOI21_X1 i_0_2_666 (.A(n_0_2_646), .B1(n_0_2_647), .B2(n_0_2_672), .ZN(
      n_0_2_645));
   NOR2_X1 i_0_2_667 (.A1(n_0_2_673), .A2(n_0_2_363), .ZN(n_0_2_646));
   AOI21_X1 i_0_2_668 (.A(n_0_2_648), .B1(n_0_2_670), .B2(n_0_2_281), .ZN(
      n_0_2_647));
   INV_X1 i_0_2_669 (.A(n_0_2_649), .ZN(n_0_2_648));
   OAI21_X1 i_0_2_670 (.A(n_0_2_650), .B1(n_0_2_670), .B2(n_0_2_281), .ZN(
      n_0_2_649));
   AOI21_X1 i_0_2_671 (.A(n_0_2_651), .B1(n_0_2_652), .B2(n_0_2_666), .ZN(
      n_0_2_650));
   NOR2_X1 i_0_2_672 (.A1(n_0_2_668), .A2(n_0_2_209), .ZN(n_0_2_651));
   AOI21_X1 i_0_2_673 (.A(n_0_2_653), .B1(n_0_2_665), .B2(n_0_2_147), .ZN(
      n_0_2_652));
   INV_X1 i_0_2_674 (.A(n_0_2_654), .ZN(n_0_2_653));
   OAI21_X1 i_0_2_675 (.A(n_0_2_655), .B1(n_0_2_665), .B2(n_0_2_147), .ZN(
      n_0_2_654));
   AOI21_X1 i_0_2_676 (.A(n_0_2_656), .B1(n_0_2_657), .B2(n_0_2_663), .ZN(
      n_0_2_655));
   NOR2_X1 i_0_2_677 (.A1(n_0_2_664), .A2(n_0_2_96), .ZN(n_0_2_656));
   AOI21_X1 i_0_2_678 (.A(n_0_2_658), .B1(n_0_2_662), .B2(n_0_2_54), .ZN(
      n_0_2_657));
   INV_X1 i_0_2_679 (.A(n_0_2_659), .ZN(n_0_2_658));
   OAI21_X1 i_0_2_680 (.A(n_0_2_661), .B1(n_0_2_662), .B2(n_0_2_54), .ZN(
      n_0_2_659));
   OAI22_X1 i_0_2_681 (.A1(n_0_2_738), .A2(n_0_2_705), .B1(n_0_2_703), .B2(
      n_0_2_221), .ZN(n_0_2_661));
   OAI21_X1 i_0_2_682 (.A(n_0_2_1412), .B1(n_0_2_705), .B2(n_0_2_745), .ZN(
      n_0_2_662));
   NAND2_X1 i_0_2_683 (.A1(n_0_2_664), .A2(n_0_2_96), .ZN(n_0_2_663));
   OAI22_X1 i_0_2_684 (.A1(n_0_2_737), .A2(n_0_2_705), .B1(n_0_2_703), .B2(
      n_0_2_227), .ZN(n_0_2_664));
   OAI22_X1 i_0_2_685 (.A1(n_0_2_1585), .A2(n_0_2_705), .B1(n_0_2_703), .B2(
      n_0_2_736), .ZN(n_0_2_665));
   NAND2_X1 i_0_2_686 (.A1(n_0_2_668), .A2(n_0_2_209), .ZN(n_0_2_666));
   OAI22_X1 i_0_2_687 (.A1(n_0_2_669), .A2(n_0_2_705), .B1(n_0_2_703), .B2(
      n_0_2_266), .ZN(n_0_2_668));
   XNOR2_X1 i_0_2_688 (.A(n_0_2_1591), .B(n_0_2_735), .ZN(n_0_2_669));
   OAI22_X1 i_0_2_689 (.A1(n_0_2_705), .A2(n_0_2_671), .B1(n_0_2_703), .B2(
      n_0_2_263), .ZN(n_0_2_670));
   XNOR2_X1 i_0_2_690 (.A(n_0_2_1598), .B(n_0_2_733), .ZN(n_0_2_671));
   NAND2_X1 i_0_2_691 (.A1(n_0_2_673), .A2(n_0_2_363), .ZN(n_0_2_672));
   OAI22_X1 i_0_2_692 (.A1(n_0_2_705), .A2(n_0_2_674), .B1(n_0_2_703), .B2(
      n_0_2_260), .ZN(n_0_2_673));
   XNOR2_X1 i_0_2_693 (.A(n_0_2_23), .B(n_0_2_731), .ZN(n_0_2_674));
   OAI22_X1 i_0_2_694 (.A1(n_0_2_705), .A2(n_0_2_676), .B1(n_0_2_703), .B2(
      n_0_2_257), .ZN(n_0_2_675));
   XNOR2_X1 i_0_2_695 (.A(n_0_2_21), .B(n_0_2_729), .ZN(n_0_2_676));
   NAND2_X1 i_0_2_696 (.A1(n_0_2_678), .A2(n_0_2_458), .ZN(n_0_2_677));
   OAI22_X1 i_0_2_697 (.A1(n_0_2_705), .A2(n_0_2_679), .B1(n_0_2_703), .B2(
      n_0_2_743), .ZN(n_0_2_678));
   XNOR2_X1 i_0_2_698 (.A(n_0_2_19), .B(n_0_2_727), .ZN(n_0_2_679));
   OAI22_X1 i_0_2_699 (.A1(n_0_2_705), .A2(n_0_2_681), .B1(n_0_2_703), .B2(
      n_0_2_252), .ZN(n_0_2_680));
   XNOR2_X1 i_0_2_700 (.A(n_0_2_17), .B(n_0_2_725), .ZN(n_0_2_681));
   NAND2_X1 i_0_2_701 (.A1(n_0_2_683), .A2(n_0_2_780), .ZN(n_0_2_682));
   OAI22_X1 i_0_2_702 (.A1(n_0_2_705), .A2(n_0_2_684), .B1(n_0_2_703), .B2(
      n_0_2_742), .ZN(n_0_2_683));
   XNOR2_X1 i_0_2_703 (.A(n_0_2_15), .B(n_0_2_723), .ZN(n_0_2_684));
   OAI22_X1 i_0_2_704 (.A1(n_0_2_705), .A2(n_0_2_686), .B1(n_0_2_703), .B2(
      n_0_2_247), .ZN(n_0_2_685));
   XNOR2_X1 i_0_2_705 (.A(n_0_2_13), .B(n_0_2_721), .ZN(n_0_2_686));
   NAND2_X1 i_0_2_706 (.A1(n_0_2_688), .A2(n_0_2_1044), .ZN(n_0_2_687));
   OAI22_X1 i_0_2_707 (.A1(n_0_2_705), .A2(n_0_2_689), .B1(n_0_2_703), .B2(
      n_0_2_244), .ZN(n_0_2_688));
   XNOR2_X1 i_0_2_708 (.A(n_0_2_11), .B(n_0_2_719), .ZN(n_0_2_689));
   OAI22_X1 i_0_2_709 (.A1(n_0_2_705), .A2(n_0_2_691), .B1(n_0_2_703), .B2(
      n_0_2_741), .ZN(n_0_2_690));
   XNOR2_X1 i_0_2_710 (.A(n_0_2_9), .B(n_0_2_717), .ZN(n_0_2_691));
   NAND2_X1 i_0_2_711 (.A1(n_0_2_693), .A2(n_0_2_1352), .ZN(n_0_2_692));
   OAI22_X1 i_0_2_712 (.A1(n_0_2_705), .A2(n_0_2_694), .B1(n_0_2_703), .B2(
      n_0_2_239), .ZN(n_0_2_693));
   XNOR2_X1 i_0_2_713 (.A(n_0_2_7), .B(n_0_2_715), .ZN(n_0_2_694));
   OAI22_X1 i_0_2_714 (.A1(n_0_2_705), .A2(n_0_2_696), .B1(n_0_2_703), .B2(
      n_0_2_236), .ZN(n_0_2_695));
   XNOR2_X1 i_0_2_715 (.A(n_0_2_5), .B(n_0_2_713), .ZN(n_0_2_696));
   NAND2_X1 i_0_2_716 (.A1(n_0_2_698), .A2(n_0_2_52), .ZN(n_0_2_697));
   OAI22_X1 i_0_2_717 (.A1(n_0_2_705), .A2(n_0_2_699), .B1(n_0_2_703), .B2(
      n_0_2_740), .ZN(n_0_2_698));
   XNOR2_X1 i_0_2_718 (.A(n_0_2_3), .B(n_0_2_711), .ZN(n_0_2_699));
   INV_X1 i_0_2_719 (.A(n_0_2_701), .ZN(n_0_2_700));
   OAI22_X1 i_0_2_720 (.A1(n_0_2_705), .A2(n_0_2_702), .B1(n_0_2_703), .B2(
      n_0_2_739), .ZN(n_0_2_701));
   XNOR2_X1 i_0_2_721 (.A(n_0_2_1), .B(n_0_2_709), .ZN(n_0_2_702));
   NOR4_X1 i_0_2_722 (.A1(n_0_2_706), .A2(n_0_2_1433), .A3(n_0_2_1432), .A4(
      n_0_2_1435), .ZN(n_0_2_703));
   NOR2_X1 i_0_2_723 (.A1(n_0_2_1395), .A2(n_0_2_705), .ZN(quotient[5]));
   INV_X1 i_0_2_724 (.A(n_0_2_705), .ZN(n_0_2_704));
   OR3_X1 i_0_2_725 (.A1(n_0_2_706), .A2(n_0_2_1432), .A3(n_0_2_45), .ZN(
      n_0_2_705));
   XNOR2_X1 i_0_2_726 (.A(n_0_2_1436), .B(n_0_2_707), .ZN(n_0_2_706));
   NAND2_X1 i_0_2_727 (.A1(n_0_2_708), .A2(n_0_2_0), .ZN(n_0_2_707));
   OAI21_X1 i_0_2_728 (.A(n_0_2_709), .B1(n_0_2_52), .B2(n_0_2_1570), .ZN(
      n_0_2_708));
   NAND2_X1 i_0_2_729 (.A1(n_0_2_710), .A2(n_0_2_2), .ZN(n_0_2_709));
   OAI21_X1 i_0_2_730 (.A(n_0_2_711), .B1(n_0_2_1516), .B2(n_0_2_1567), .ZN(
      n_0_2_710));
   NAND2_X1 i_0_2_731 (.A1(n_0_2_712), .A2(n_0_2_4), .ZN(n_0_2_711));
   OAI21_X1 i_0_2_732 (.A(n_0_2_713), .B1(n_0_2_1352), .B2(n_0_2_1564), .ZN(
      n_0_2_712));
   NAND2_X1 i_0_2_733 (.A1(n_0_2_714), .A2(n_0_2_6), .ZN(n_0_2_713));
   OAI21_X1 i_0_2_734 (.A(n_0_2_715), .B1(n_0_2_1190), .B2(n_0_2_1561), .ZN(
      n_0_2_714));
   NAND2_X1 i_0_2_735 (.A1(n_0_2_716), .A2(n_0_2_8), .ZN(n_0_2_715));
   OAI21_X1 i_0_2_736 (.A(n_0_2_717), .B1(n_0_2_1044), .B2(n_0_2_1558), .ZN(
      n_0_2_716));
   NAND2_X1 i_0_2_737 (.A1(n_0_2_718), .A2(n_0_2_10), .ZN(n_0_2_717));
   OAI21_X1 i_0_2_738 (.A(n_0_2_719), .B1(n_0_2_907), .B2(n_0_2_1555), .ZN(
      n_0_2_718));
   NAND2_X1 i_0_2_739 (.A1(n_0_2_720), .A2(n_0_2_12), .ZN(n_0_2_719));
   OAI21_X1 i_0_2_740 (.A(n_0_2_721), .B1(n_0_2_780), .B2(n_0_2_1552), .ZN(
      n_0_2_720));
   NAND2_X1 i_0_2_741 (.A1(n_0_2_722), .A2(n_0_2_14), .ZN(n_0_2_721));
   OAI21_X1 i_0_2_742 (.A(n_0_2_723), .B1(n_0_2_660), .B2(n_0_2_1549), .ZN(
      n_0_2_722));
   NAND2_X1 i_0_2_743 (.A1(n_0_2_724), .A2(n_0_2_16), .ZN(n_0_2_723));
   OAI21_X1 i_0_2_744 (.A(n_0_2_725), .B1(n_0_2_458), .B2(n_0_2_1546), .ZN(
      n_0_2_724));
   NAND2_X1 i_0_2_745 (.A1(n_0_2_726), .A2(n_0_2_18), .ZN(n_0_2_725));
   OAI21_X1 i_0_2_746 (.A(n_0_2_727), .B1(n_0_2_453), .B2(n_0_2_1543), .ZN(
      n_0_2_726));
   NAND2_X1 i_0_2_747 (.A1(n_0_2_728), .A2(n_0_2_20), .ZN(n_0_2_727));
   OAI21_X1 i_0_2_748 (.A(n_0_2_729), .B1(n_0_2_363), .B2(n_0_2_1540), .ZN(
      n_0_2_728));
   NAND2_X1 i_0_2_749 (.A1(n_0_2_730), .A2(n_0_2_22), .ZN(n_0_2_729));
   OAI21_X1 i_0_2_750 (.A(n_0_2_731), .B1(n_0_2_281), .B2(n_0_2_1537), .ZN(
      n_0_2_730));
   NAND2_X1 i_0_2_751 (.A1(n_0_2_732), .A2(n_0_2_1602), .ZN(n_0_2_731));
   OAI21_X1 i_0_2_752 (.A(n_0_2_733), .B1(n_0_2_209), .B2(n_0_2_1534), .ZN(
      n_0_2_732));
   NAND2_X1 i_0_2_753 (.A1(n_0_2_734), .A2(n_0_2_1595), .ZN(n_0_2_733));
   OAI21_X1 i_0_2_754 (.A(n_0_2_735), .B1(n_0_2_147), .B2(n_0_2_1531), .ZN(
      n_0_2_734));
   NAND3_X1 i_0_2_755 (.A1(n_0_2_1588), .A2(n_0_2_1589), .A3(n_0_2_1590), 
      .ZN(n_0_2_735));
   INV_X1 i_0_2_756 (.A(n_0_2_1528), .ZN(n_0_2_736));
   INV_X1 i_0_2_757 (.A(n_0_2_1579), .ZN(n_0_2_737));
   INV_X1 i_0_2_758 (.A(n_0_2_1573), .ZN(n_0_2_738));
   INV_X1 i_0_2_759 (.A(n_0_2_1570), .ZN(n_0_2_739));
   INV_X1 i_0_2_760 (.A(n_0_2_1567), .ZN(n_0_2_740));
   INV_X1 i_0_2_761 (.A(n_0_2_1558), .ZN(n_0_2_741));
   INV_X1 i_0_2_762 (.A(n_0_2_1549), .ZN(n_0_2_742));
   INV_X1 i_0_2_763 (.A(n_0_2_1543), .ZN(n_0_2_743));
   NAND2_X1 i_0_2_764 (.A1(n_0_2_53), .A2(n_0_2_46), .ZN(n_0_2_45));
   INV_X1 i_0_2_765 (.A(n_0_2_47), .ZN(n_0_2_46));
   NAND2_X1 i_0_2_766 (.A1(n_0_2_1437), .A2(n_0_2_50), .ZN(n_0_2_47));
   AND2_X1 i_0_2_767 (.A1(n_0_2_56), .A2(n_0_2_1431), .ZN(n_0_2_744));
   NAND2_X1 i_0_2_768 (.A1(in_b[0]), .A2(n_0_2_49), .ZN(n_0_2_745));
   NOR4_X1 i_0_2_769 (.A1(n_0_53), .A2(n_0_52), .A3(n_0_54), .A4(n_0_51), 
      .ZN(n_0_2_746));
   INV_X1 i_0_2_770 (.A(n_0_2_747), .ZN(n_0_2_48));
   NOR2_X1 i_0_2_771 (.A1(n_0_59), .A2(n_0_58), .ZN(n_0_2_747));
   INV_X1 i_0_2_772 (.A(n_0_2_749), .ZN(n_0_2_748));
   NAND2_X1 i_0_2_773 (.A1(n_0_2_1412), .A2(n_0_2_1367), .ZN(n_0_2_749));
   OAI21_X1 i_0_2_774 (.A(n_0_2_1247), .B1(in_b[0]), .B2(n_0_2_1444), .ZN(
      n_0_2_1246));
   NAND2_X1 i_0_2_775 (.A1(n_0_2_1430), .A2(n_0_2_1516), .ZN(n_0_2_750));
   XOR2_X1 i_0_2_776 (.A(n_0_2_1190), .B(n_0_2_769), .Z(n_0_2_751));
   OAI21_X1 i_0_2_777 (.A(n_0_2_771), .B1(n_0_2_1044), .B2(n_0_2_772), .ZN(
      n_0_2_752));
   AOI22_X1 i_0_2_778 (.A1(n_0_2_907), .A2(n_0_2_776), .B1(n_0_2_1421), .B2(
      n_0_2_775), .ZN(n_0_2_753));
   XOR2_X1 i_0_2_779 (.A(n_0_2_835), .B(n_0_2_779), .Z(n_0_2_754));
   XNOR2_X1 i_0_2_780 (.A(n_0_2_830), .B(n_0_2_781), .ZN(n_0_2_755));
   XOR2_X1 i_0_2_781 (.A(n_0_2_827), .B(n_0_2_782), .Z(n_0_2_756));
   XNOR2_X1 i_0_2_782 (.A(n_0_2_822), .B(n_0_2_783), .ZN(n_0_2_757));
   XOR2_X1 i_0_2_783 (.A(n_0_2_819), .B(n_0_2_784), .Z(n_0_2_758));
   XNOR2_X1 i_0_2_784 (.A(n_0_2_814), .B(n_0_2_785), .ZN(n_0_2_759));
   XOR2_X1 i_0_2_785 (.A(n_0_2_788), .B(n_0_2_787), .Z(n_0_2_760));
   XOR2_X1 i_0_2_786 (.A(n_0_2_808), .B(n_0_2_790), .Z(n_0_2_761));
   XNOR2_X1 i_0_2_787 (.A(n_0_2_804), .B(n_0_2_791), .ZN(n_0_2_762));
   XOR2_X1 i_0_2_788 (.A(n_0_2_794), .B(n_0_2_793), .Z(n_0_2_763));
   XNOR2_X1 i_0_2_789 (.A(n_0_2_795), .B(n_0_2_765), .ZN(n_0_2_764));
   OAI22_X1 i_0_2_790 (.A1(n_0_2_1367), .A2(n_0_2_799), .B1(n_0_2_1398), 
      .B2(n_0_2_798), .ZN(n_0_2_765));
   NOR2_X1 i_0_2_791 (.A1(n_0_2_49), .A2(n_0_2_1247), .ZN(n_0_2_766));
   NAND2_X1 i_0_2_792 (.A1(n_0_2_49), .A2(n_0_2_1247), .ZN(n_0_2_1255));
   INV_X1 i_0_2_793 (.A(n_0_2_1247), .ZN(n_0_2_767));
   NAND2_X1 i_0_2_794 (.A1(in_b[0]), .A2(n_0_2_1444), .ZN(n_0_2_1247));
   INV_X1 i_0_2_795 (.A(n_0_2_768), .ZN(n_0_2_1091));
   AOI21_X1 i_0_2_796 (.A(n_0_2_798), .B1(n_0_2_1405), .B2(n_0_2_799), .ZN(
      n_0_2_768));
   AND2_X1 i_0_2_797 (.A1(n_0_2_53), .A2(n_0_2_1196), .ZN(n_0_2_287));
   AND2_X1 i_0_2_798 (.A1(n_0_2_52), .A2(n_0_2_1426), .ZN(n_0_2_1196));
   AOI21_X1 i_0_2_799 (.A(n_0_2_876), .B1(n_0_2_878), .B2(n_0_2_875), .ZN(
      n_0_2_769));
   INV_X1 i_0_2_800 (.A(n_0_2_771), .ZN(n_0_2_770));
   NAND2_X1 i_0_2_801 (.A1(n_0_2_1044), .A2(n_0_2_772), .ZN(n_0_2_771));
   XNOR2_X1 i_0_2_802 (.A(n_0_2_880), .B(n_0_2_773), .ZN(n_0_2_772));
   OAI211_X1 i_0_2_803 (.A(n_0_2_882), .B(n_0_2_875), .C1(n_0_2_1421), .C2(
      n_0_2_884), .ZN(n_0_2_773));
   NAND2_X1 i_0_2_804 (.A1(n_0_2_907), .A2(n_0_2_776), .ZN(n_0_2_774));
   INV_X1 i_0_2_805 (.A(n_0_2_776), .ZN(n_0_2_775));
   XNOR2_X1 i_0_2_806 (.A(n_0_2_885), .B(n_0_2_777), .ZN(n_0_2_776));
   OAI211_X1 i_0_2_807 (.A(n_0_2_887), .B(n_0_2_875), .C1(n_0_2_1440), .C2(
      n_0_2_889), .ZN(n_0_2_777));
   OAI22_X1 i_0_2_808 (.A1(n_0_2_780), .A2(n_0_2_836), .B1(n_0_2_834), .B2(
      n_0_2_779), .ZN(n_0_2_778));
   AOI22_X1 i_0_2_809 (.A1(n_0_2_1418), .A2(n_0_2_832), .B1(n_0_2_830), .B2(
      n_0_2_781), .ZN(n_0_2_779));
   OAI22_X1 i_0_2_810 (.A1(n_0_2_458), .A2(n_0_2_828), .B1(n_0_2_826), .B2(
      n_0_2_782), .ZN(n_0_2_781));
   AOI22_X1 i_0_2_811 (.A1(n_0_2_1415), .A2(n_0_2_824), .B1(n_0_2_822), .B2(
      n_0_2_783), .ZN(n_0_2_782));
   OAI22_X1 i_0_2_812 (.A1(n_0_2_363), .A2(n_0_2_820), .B1(n_0_2_818), .B2(
      n_0_2_784), .ZN(n_0_2_783));
   AOI22_X1 i_0_2_813 (.A1(n_0_2_1410), .A2(n_0_2_815), .B1(n_0_2_814), .B2(
      n_0_2_785), .ZN(n_0_2_784));
   OAI22_X1 i_0_2_814 (.A1(n_0_2_209), .A2(n_0_2_812), .B1(n_0_2_788), .B2(
      n_0_2_786), .ZN(n_0_2_785));
   INV_X1 i_0_2_815 (.A(n_0_2_787), .ZN(n_0_2_786));
   XNOR2_X1 i_0_2_816 (.A(n_0_2_1408), .B(n_0_2_812), .ZN(n_0_2_787));
   AOI22_X1 i_0_2_817 (.A1(n_0_2_1406), .A2(n_0_2_810), .B1(n_0_2_808), .B2(
      n_0_2_789), .ZN(n_0_2_788));
   INV_X1 i_0_2_818 (.A(n_0_2_790), .ZN(n_0_2_789));
   AOI22_X1 i_0_2_819 (.A1(n_0_2_1403), .A2(n_0_2_805), .B1(n_0_2_804), .B2(
      n_0_2_791), .ZN(n_0_2_790));
   OAI22_X1 i_0_2_820 (.A1(n_0_2_54), .A2(n_0_2_800), .B1(n_0_2_794), .B2(
      n_0_2_792), .ZN(n_0_2_791));
   INV_X1 i_0_2_821 (.A(n_0_2_793), .ZN(n_0_2_792));
   AOI22_X1 i_0_2_822 (.A1(n_0_2_1400), .A2(n_0_2_801), .B1(n_0_2_54), .B2(
      n_0_2_800), .ZN(n_0_2_793));
   OAI22_X1 i_0_2_823 (.A1(n_0_2_797), .A2(n_0_2_795), .B1(n_0_2_1398), .B2(
      n_0_2_798), .ZN(n_0_2_794));
   XNOR2_X1 i_0_2_824 (.A(n_0_2_939), .B(n_0_2_796), .ZN(n_0_2_795));
   NAND2_X1 i_0_2_825 (.A1(in_b[0]), .A2(n_0_2_875), .ZN(n_0_2_796));
   NOR2_X1 i_0_2_826 (.A1(n_0_2_1367), .A2(n_0_2_799), .ZN(n_0_2_797));
   NOR2_X1 i_0_2_827 (.A1(n_0_2_1405), .A2(n_0_2_799), .ZN(n_0_2_798));
   AOI21_X1 i_0_2_828 (.A(n_0_2_1392), .B1(in_a[1]), .B2(n_0_2_1393), .ZN(
      n_0_2_799));
   INV_X1 i_0_2_829 (.A(n_0_2_801), .ZN(n_0_2_800));
   XNOR2_X1 i_0_2_830 (.A(n_0_2_937), .B(n_0_2_802), .ZN(n_0_2_801));
   NAND2_X1 i_0_2_831 (.A1(n_0_2_875), .A2(n_0_2_803), .ZN(n_0_2_802));
   AOI21_X1 i_0_2_832 (.A(n_0_2_935), .B1(n_0_2_1366), .B2(n_0_2_939), .ZN(
      n_0_2_803));
   AOI22_X1 i_0_2_833 (.A1(n_0_2_1403), .A2(n_0_2_805), .B1(n_0_2_96), .B2(
      n_0_2_806), .ZN(n_0_2_804));
   INV_X1 i_0_2_834 (.A(n_0_2_806), .ZN(n_0_2_805));
   XNOR2_X1 i_0_2_835 (.A(n_0_2_930), .B(n_0_2_807), .ZN(n_0_2_806));
   NOR3_X1 i_0_2_836 (.A1(n_0_2_933), .A2(n_0_2_932), .A3(n_0_2_874), .ZN(
      n_0_2_807));
   AOI22_X1 i_0_2_837 (.A1(n_0_2_1406), .A2(n_0_2_810), .B1(n_0_2_147), .B2(
      n_0_2_809), .ZN(n_0_2_808));
   INV_X1 i_0_2_838 (.A(n_0_2_810), .ZN(n_0_2_809));
   XNOR2_X1 i_0_2_839 (.A(n_0_2_925), .B(n_0_2_811), .ZN(n_0_2_810));
   OAI211_X1 i_0_2_840 (.A(n_0_2_928), .B(n_0_2_875), .C1(n_0_2_96), .C2(
      n_0_2_929), .ZN(n_0_2_811));
   XNOR2_X1 i_0_2_841 (.A(n_0_2_920), .B(n_0_2_813), .ZN(n_0_2_812));
   AOI211_X1 i_0_2_842 (.A(n_0_2_922), .B(n_0_2_874), .C1(n_0_2_147), .C2(
      n_0_2_924), .ZN(n_0_2_813));
   AOI22_X1 i_0_2_843 (.A1(n_0_2_1410), .A2(n_0_2_815), .B1(n_0_2_281), .B2(
      n_0_2_816), .ZN(n_0_2_814));
   INV_X1 i_0_2_844 (.A(n_0_2_816), .ZN(n_0_2_815));
   XNOR2_X1 i_0_2_845 (.A(n_0_2_915), .B(n_0_2_817), .ZN(n_0_2_816));
   AOI211_X1 i_0_2_846 (.A(n_0_2_917), .B(n_0_2_874), .C1(n_0_2_209), .C2(
      n_0_2_919), .ZN(n_0_2_817));
   INV_X1 i_0_2_847 (.A(n_0_2_819), .ZN(n_0_2_818));
   XNOR2_X1 i_0_2_848 (.A(n_0_2_1413), .B(n_0_2_820), .ZN(n_0_2_819));
   XNOR2_X1 i_0_2_849 (.A(n_0_2_910), .B(n_0_2_821), .ZN(n_0_2_820));
   AOI211_X1 i_0_2_850 (.A(n_0_2_912), .B(n_0_2_874), .C1(n_0_2_281), .C2(
      n_0_2_914), .ZN(n_0_2_821));
   AOI22_X1 i_0_2_851 (.A1(n_0_2_1415), .A2(n_0_2_824), .B1(n_0_2_453), .B2(
      n_0_2_823), .ZN(n_0_2_822));
   INV_X1 i_0_2_852 (.A(n_0_2_824), .ZN(n_0_2_823));
   XNOR2_X1 i_0_2_853 (.A(n_0_2_904), .B(n_0_2_825), .ZN(n_0_2_824));
   AOI221_X1 i_0_2_854 (.A(n_0_2_874), .B1(n_0_2_363), .B2(n_0_2_909), .C1(
      n_0_2_1413), .C2(n_0_2_908), .ZN(n_0_2_825));
   INV_X1 i_0_2_855 (.A(n_0_2_827), .ZN(n_0_2_826));
   XNOR2_X1 i_0_2_856 (.A(n_0_2_1417), .B(n_0_2_828), .ZN(n_0_2_827));
   XNOR2_X1 i_0_2_857 (.A(n_0_2_940), .B(n_0_2_829), .ZN(n_0_2_828));
   AOI221_X1 i_0_2_858 (.A(n_0_2_874), .B1(n_0_2_1415), .B2(n_0_2_901), .C1(
      n_0_2_453), .C2(n_0_2_902), .ZN(n_0_2_829));
   AOI22_X1 i_0_2_859 (.A1(n_0_2_1418), .A2(n_0_2_832), .B1(n_0_2_660), .B2(
      n_0_2_831), .ZN(n_0_2_830));
   INV_X1 i_0_2_860 (.A(n_0_2_832), .ZN(n_0_2_831));
   XNOR2_X1 i_0_2_861 (.A(n_0_2_895), .B(n_0_2_833), .ZN(n_0_2_832));
   OAI211_X1 i_0_2_862 (.A(n_0_2_898), .B(n_0_2_875), .C1(n_0_2_458), .C2(
      n_0_2_899), .ZN(n_0_2_833));
   INV_X1 i_0_2_863 (.A(n_0_2_835), .ZN(n_0_2_834));
   AOI22_X1 i_0_2_864 (.A1(n_0_2_1440), .A2(n_0_2_837), .B1(n_0_2_780), .B2(
      n_0_2_836), .ZN(n_0_2_835));
   INV_X1 i_0_2_865 (.A(n_0_2_837), .ZN(n_0_2_836));
   XNOR2_X1 i_0_2_866 (.A(n_0_2_890), .B(n_0_2_838), .ZN(n_0_2_837));
   AOI211_X1 i_0_2_867 (.A(n_0_2_893), .B(n_0_2_874), .C1(n_0_2_660), .C2(
      n_0_2_894), .ZN(n_0_2_838));
   INV_X1 i_0_2_868 (.A(n_0_2_839), .ZN(n_0_50));
   AOI22_X1 i_0_2_869 (.A1(quotient[9]), .A2(n_0_2_846), .B1(n_0_31), .B2(
      n_0_2_847), .ZN(n_0_2_839));
   INV_X1 i_0_2_870 (.A(n_0_2_840), .ZN(n_0_51));
   AOI22_X1 i_0_2_871 (.A1(quotient[10]), .A2(n_0_2_846), .B1(n_0_32), .B2(
      n_0_2_847), .ZN(n_0_2_840));
   INV_X1 i_0_2_872 (.A(n_0_2_841), .ZN(n_0_52));
   AOI22_X1 i_0_2_873 (.A1(quotient[11]), .A2(n_0_2_846), .B1(n_0_33), .B2(
      n_0_2_847), .ZN(n_0_2_841));
   INV_X1 i_0_2_874 (.A(n_0_2_842), .ZN(n_0_53));
   AOI22_X1 i_0_2_875 (.A1(quotient[12]), .A2(n_0_2_846), .B1(n_0_34), .B2(
      n_0_2_847), .ZN(n_0_2_842));
   INV_X1 i_0_2_876 (.A(n_0_2_843), .ZN(n_0_54));
   AOI22_X1 i_0_2_877 (.A1(quotient[13]), .A2(n_0_2_846), .B1(n_0_35), .B2(
      n_0_2_847), .ZN(n_0_2_843));
   INV_X1 i_0_2_878 (.A(n_0_2_844), .ZN(n_0_55));
   AOI22_X1 i_0_2_879 (.A1(quotient[14]), .A2(n_0_2_846), .B1(n_0_36), .B2(
      n_0_2_847), .ZN(n_0_2_844));
   INV_X1 i_0_2_880 (.A(n_0_2_845), .ZN(n_0_56));
   AOI22_X1 i_0_2_881 (.A1(quotient[15]), .A2(n_0_2_846), .B1(n_0_37), .B2(
      n_0_2_847), .ZN(n_0_2_845));
   AND2_X1 i_0_2_882 (.A1(n_0_38), .A2(n_0_2_847), .ZN(n_0_57));
   INV_X1 i_0_2_883 (.A(n_0_2_847), .ZN(n_0_2_846));
   XNOR2_X1 i_0_2_884 (.A(in_b[15]), .B(n_0_2_1451), .ZN(n_0_2_847));
   INV_X1 i_0_2_885 (.A(n_0_2_848), .ZN(n_0_58));
   AOI21_X1 i_0_2_886 (.A(divide_by_zero_error), .B1(n_0_2_856), .B2(n_0_2_849), 
      .ZN(n_0_2_848));
   NOR4_X1 i_0_2_887 (.A1(n_0_2_866), .A2(n_0_2_862), .A3(n_0_2_853), .A4(
      n_0_2_850), .ZN(n_0_2_849));
   NAND3_X1 i_0_2_888 (.A1(n_0_2_1405), .A2(n_0_2_851), .A3(n_0_2_852), .ZN(
      n_0_2_850));
   NOR3_X1 i_0_2_889 (.A1(in_b[3]), .A2(in_b[2]), .A3(in_b[1]), .ZN(n_0_2_851));
   NOR4_X1 i_0_2_890 (.A1(in_b[7]), .A2(in_b[6]), .A3(in_b[5]), .A4(in_b[4]), 
      .ZN(n_0_2_852));
   NAND3_X1 i_0_2_891 (.A1(n_0_2_1453), .A2(n_0_2_855), .A3(n_0_2_854), .ZN(
      n_0_2_853));
   NOR4_X1 i_0_2_892 (.A1(in_b[16]), .A2(in_b[15]), .A3(in_b[14]), .A4(in_b[13]), 
      .ZN(n_0_2_854));
   NOR3_X1 i_0_2_893 (.A1(in_b[12]), .A2(in_b[10]), .A3(in_b[9]), .ZN(n_0_2_855));
   NOR2_X1 i_0_2_894 (.A1(in_b[21]), .A2(n_0_2_857), .ZN(n_0_2_856));
   NAND3_X1 i_0_2_895 (.A1(n_0_2_861), .A2(n_0_2_860), .A3(n_0_2_858), .ZN(
      n_0_2_857));
   NOR4_X1 i_0_2_896 (.A1(in_b[24]), .A2(in_b[23]), .A3(in_b[22]), .A4(n_0_2_859), 
      .ZN(n_0_2_858));
   OR4_X1 i_0_2_897 (.A1(in_b[20]), .A2(in_b[19]), .A3(in_b[18]), .A4(in_b[17]), 
      .ZN(n_0_2_859));
   NOR4_X1 i_0_2_898 (.A1(in_b[27]), .A2(in_b[26]), .A3(in_b[32]), .A4(in_b[29]), 
      .ZN(n_0_2_860));
   NOR4_X1 i_0_2_899 (.A1(in_b[28]), .A2(in_b[25]), .A3(in_b[31]), .A4(in_b[30]), 
      .ZN(n_0_2_861));
   NAND4_X1 i_0_2_900 (.A1(n_0_2_865), .A2(n_0_2_864), .A3(n_0_2_870), .A4(
      n_0_2_863), .ZN(n_0_2_862));
   NOR4_X1 i_0_2_901 (.A1(in_b[51]), .A2(in_b[50]), .A3(in_b[56]), .A4(in_b[53]), 
      .ZN(n_0_2_863));
   NOR4_X1 i_0_2_902 (.A1(in_b[36]), .A2(in_b[33]), .A3(in_b[39]), .A4(in_b[38]), 
      .ZN(n_0_2_864));
   NOR4_X1 i_0_2_903 (.A1(in_b[43]), .A2(in_b[42]), .A3(in_b[48]), .A4(in_b[45]), 
      .ZN(n_0_2_865));
   NAND4_X1 i_0_2_904 (.A1(n_0_2_869), .A2(n_0_2_868), .A3(n_0_2_871), .A4(
      n_0_2_867), .ZN(n_0_2_866));
   NOR4_X1 i_0_2_905 (.A1(in_b[52]), .A2(in_b[49]), .A3(in_b[55]), .A4(in_b[54]), 
      .ZN(n_0_2_867));
   NOR4_X1 i_0_2_906 (.A1(in_b[35]), .A2(in_b[34]), .A3(in_b[40]), .A4(in_b[37]), 
      .ZN(n_0_2_868));
   NOR4_X1 i_0_2_907 (.A1(in_b[44]), .A2(in_b[41]), .A3(in_b[47]), .A4(in_b[46]), 
      .ZN(n_0_2_869));
   NOR4_X1 i_0_2_908 (.A1(in_b[60]), .A2(in_b[59]), .A3(in_b[58]), .A4(in_b[57]), 
      .ZN(n_0_2_870));
   NOR4_X1 i_0_2_909 (.A1(in_b[63]), .A2(in_b[11]), .A3(in_b[62]), .A4(in_b[61]), 
      .ZN(n_0_2_871));
   AOI21_X1 i_0_2_910 (.A(n_0_2_1395), .B1(n_0_2_873), .B2(n_0_2_872), .ZN(
      n_0_59));
   AOI211_X1 i_0_2_911 (.A(n_0_2_1360), .B(n_0_2_1254), .C1(n_0_2_1396), 
      .C2(n_0_2_1371), .ZN(n_0_2_872));
   NOR4_X1 i_0_2_912 (.A1(n_0_2_1343), .A2(n_0_2_1331), .A3(n_0_2_1309), 
      .A4(n_0_2_1282), .ZN(n_0_2_873));
   NOR2_X1 i_0_2_913 (.A1(n_0_2_1395), .A2(n_0_2_874), .ZN(quotient[9]));
   INV_X1 i_0_2_914 (.A(n_0_2_875), .ZN(n_0_2_874));
   AOI221_X1 i_0_2_915 (.A(n_0_2_1425), .B1(n_0_2_1424), .B2(n_0_2_879), 
      .C1(n_0_2_878), .C2(n_0_2_876), .ZN(n_0_2_875));
   INV_X1 i_0_2_916 (.A(n_0_2_877), .ZN(n_0_2_876));
   AOI21_X1 i_0_2_917 (.A(n_0_2_1007), .B1(n_0_2_944), .B2(n_0_2_943), .ZN(
      n_0_2_877));
   OR2_X1 i_0_2_918 (.A1(n_0_2_1424), .A2(n_0_2_879), .ZN(n_0_2_878));
   OAI21_X1 i_0_2_919 (.A(n_0_2_882), .B1(n_0_2_883), .B2(n_0_2_880), .ZN(
      n_0_2_879));
   XNOR2_X1 i_0_2_920 (.A(n_0_2_946), .B(n_0_2_881), .ZN(n_0_2_880));
   OAI211_X1 i_0_2_921 (.A(n_0_2_949), .B(n_0_2_943), .C1(n_0_2_1440), .C2(
      n_0_2_950), .ZN(n_0_2_881));
   NAND2_X1 i_0_2_922 (.A1(n_0_2_1421), .A2(n_0_2_884), .ZN(n_0_2_882));
   NOR2_X1 i_0_2_923 (.A1(n_0_2_1421), .A2(n_0_2_884), .ZN(n_0_2_883));
   OAI21_X1 i_0_2_924 (.A(n_0_2_887), .B1(n_0_2_888), .B2(n_0_2_885), .ZN(
      n_0_2_884));
   XNOR2_X1 i_0_2_925 (.A(n_0_2_951), .B(n_0_2_886), .ZN(n_0_2_885));
   OAI211_X1 i_0_2_926 (.A(n_0_2_954), .B(n_0_2_943), .C1(n_0_2_1418), .C2(
      n_0_2_955), .ZN(n_0_2_886));
   NAND2_X1 i_0_2_927 (.A1(n_0_2_1440), .A2(n_0_2_889), .ZN(n_0_2_887));
   NOR2_X1 i_0_2_928 (.A1(n_0_2_1440), .A2(n_0_2_889), .ZN(n_0_2_888));
   AOI22_X1 i_0_2_929 (.A1(n_0_2_660), .A2(n_0_2_894), .B1(n_0_2_892), .B2(
      n_0_2_890), .ZN(n_0_2_889));
   XNOR2_X1 i_0_2_930 (.A(n_0_2_956), .B(n_0_2_891), .ZN(n_0_2_890));
   OAI211_X1 i_0_2_931 (.A(n_0_2_959), .B(n_0_2_943), .C1(n_0_2_1417), .C2(
      n_0_2_960), .ZN(n_0_2_891));
   INV_X1 i_0_2_932 (.A(n_0_2_893), .ZN(n_0_2_892));
   NOR2_X1 i_0_2_933 (.A1(n_0_2_660), .A2(n_0_2_894), .ZN(n_0_2_893));
   AOI21_X1 i_0_2_934 (.A(n_0_2_897), .B1(n_0_2_898), .B2(n_0_2_895), .ZN(
      n_0_2_894));
   XNOR2_X1 i_0_2_935 (.A(n_0_2_961), .B(n_0_2_896), .ZN(n_0_2_895));
   AND3_X1 i_0_2_936 (.A1(n_0_2_965), .A2(n_0_2_963), .A3(n_0_2_943), .ZN(
      n_0_2_896));
   NOR2_X1 i_0_2_937 (.A1(n_0_2_458), .A2(n_0_2_899), .ZN(n_0_2_897));
   NAND2_X1 i_0_2_938 (.A1(n_0_2_458), .A2(n_0_2_899), .ZN(n_0_2_898));
   AOI21_X1 i_0_2_939 (.A(n_0_2_900), .B1(n_0_2_1415), .B2(n_0_2_940), .ZN(
      n_0_2_899));
   AOI21_X1 i_0_2_940 (.A(n_0_2_902), .B1(n_0_2_453), .B2(n_0_2_941), .ZN(
      n_0_2_900));
   INV_X1 i_0_2_941 (.A(n_0_2_902), .ZN(n_0_2_901));
   AOI21_X1 i_0_2_942 (.A(n_0_2_903), .B1(n_0_2_908), .B2(n_0_2_905), .ZN(
      n_0_2_902));
   AOI21_X1 i_0_2_943 (.A(n_0_2_363), .B1(n_0_2_909), .B2(n_0_2_904), .ZN(
      n_0_2_903));
   INV_X1 i_0_2_944 (.A(n_0_2_905), .ZN(n_0_2_904));
   XNOR2_X1 i_0_2_945 (.A(n_0_2_972), .B(n_0_2_906), .ZN(n_0_2_905));
   AND3_X1 i_0_2_946 (.A1(n_0_2_976), .A2(n_0_2_974), .A3(n_0_2_943), .ZN(
      n_0_2_906));
   INV_X1 i_0_2_947 (.A(n_0_2_909), .ZN(n_0_2_908));
   AOI21_X1 i_0_2_948 (.A(n_0_2_912), .B1(n_0_2_913), .B2(n_0_2_910), .ZN(
      n_0_2_909));
   XNOR2_X1 i_0_2_949 (.A(n_0_2_978), .B(n_0_2_911), .ZN(n_0_2_910));
   AND3_X1 i_0_2_950 (.A1(n_0_2_982), .A2(n_0_2_980), .A3(n_0_2_943), .ZN(
      n_0_2_911));
   NOR2_X1 i_0_2_951 (.A1(n_0_2_281), .A2(n_0_2_914), .ZN(n_0_2_912));
   NAND2_X1 i_0_2_952 (.A1(n_0_2_281), .A2(n_0_2_914), .ZN(n_0_2_913));
   AOI21_X1 i_0_2_953 (.A(n_0_2_917), .B1(n_0_2_918), .B2(n_0_2_915), .ZN(
      n_0_2_914));
   XOR2_X1 i_0_2_954 (.A(n_0_2_984), .B(n_0_2_916), .Z(n_0_2_915));
   OAI211_X1 i_0_2_955 (.A(n_0_2_987), .B(n_0_2_943), .C1(n_0_2_1406), .C2(
      n_0_2_988), .ZN(n_0_2_916));
   NOR2_X1 i_0_2_956 (.A1(n_0_2_209), .A2(n_0_2_919), .ZN(n_0_2_917));
   NAND2_X1 i_0_2_957 (.A1(n_0_2_209), .A2(n_0_2_919), .ZN(n_0_2_918));
   AOI21_X1 i_0_2_958 (.A(n_0_2_922), .B1(n_0_2_923), .B2(n_0_2_920), .ZN(
      n_0_2_919));
   XNOR2_X1 i_0_2_959 (.A(n_0_2_989), .B(n_0_2_921), .ZN(n_0_2_920));
   AND3_X1 i_0_2_960 (.A1(n_0_2_993), .A2(n_0_2_991), .A3(n_0_2_943), .ZN(
      n_0_2_921));
   NOR2_X1 i_0_2_961 (.A1(n_0_2_147), .A2(n_0_2_924), .ZN(n_0_2_922));
   NAND2_X1 i_0_2_962 (.A1(n_0_2_147), .A2(n_0_2_924), .ZN(n_0_2_923));
   AOI21_X1 i_0_2_963 (.A(n_0_2_927), .B1(n_0_2_928), .B2(n_0_2_925), .ZN(
      n_0_2_924));
   XOR2_X1 i_0_2_964 (.A(n_0_2_995), .B(n_0_2_926), .Z(n_0_2_925));
   NAND3_X1 i_0_2_965 (.A1(n_0_2_998), .A2(n_0_2_997), .A3(n_0_2_943), .ZN(
      n_0_2_926));
   NOR2_X1 i_0_2_966 (.A1(n_0_2_96), .A2(n_0_2_929), .ZN(n_0_2_927));
   NAND2_X1 i_0_2_967 (.A1(n_0_2_96), .A2(n_0_2_929), .ZN(n_0_2_928));
   AOI21_X1 i_0_2_968 (.A(n_0_2_932), .B1(n_0_2_934), .B2(n_0_2_930), .ZN(
      n_0_2_929));
   XNOR2_X1 i_0_2_969 (.A(n_0_2_1000), .B(n_0_2_931), .ZN(n_0_2_930));
   OAI211_X1 i_0_2_970 (.A(n_0_2_1003), .B(n_0_2_943), .C1(n_0_2_1367), .C2(
      n_0_2_1004), .ZN(n_0_2_931));
   NOR3_X1 i_0_2_971 (.A1(n_0_2_936), .A2(n_0_2_935), .A3(n_0_2_54), .ZN(
      n_0_2_932));
   INV_X1 i_0_2_972 (.A(n_0_2_934), .ZN(n_0_2_933));
   OAI21_X1 i_0_2_973 (.A(n_0_2_54), .B1(n_0_2_936), .B2(n_0_2_935), .ZN(
      n_0_2_934));
   OAI21_X1 i_0_2_974 (.A(n_0_2_1412), .B1(n_0_2_1398), .B2(n_0_2_939), .ZN(
      n_0_2_935));
   AOI21_X1 i_0_2_975 (.A(n_0_2_937), .B1(n_0_2_1366), .B2(n_0_2_939), .ZN(
      n_0_2_936));
   XOR2_X1 i_0_2_976 (.A(n_0_2_1004), .B(n_0_2_938), .Z(n_0_2_937));
   NAND2_X1 i_0_2_977 (.A1(in_b[0]), .A2(n_0_2_943), .ZN(n_0_2_938));
   XOR2_X1 i_0_2_978 (.A(in_a[2]), .B(n_0_2_1006), .Z(n_0_2_939));
   INV_X1 i_0_2_979 (.A(n_0_2_941), .ZN(n_0_2_940));
   XNOR2_X1 i_0_2_980 (.A(n_0_2_967), .B(n_0_2_942), .ZN(n_0_2_941));
   OAI211_X1 i_0_2_981 (.A(n_0_2_970), .B(n_0_2_943), .C1(n_0_2_1413), .C2(
      n_0_2_971), .ZN(n_0_2_942));
   AND2_X1 i_0_2_982 (.A1(n_0_2_1394), .A2(n_0_2_943), .ZN(quotient[10]));
   AOI221_X1 i_0_2_983 (.A(n_0_2_1422), .B1(n_0_2_1421), .B2(n_0_2_945), 
      .C1(n_0_2_1007), .C2(n_0_2_944), .ZN(n_0_2_943));
   OR2_X1 i_0_2_984 (.A1(n_0_2_1421), .A2(n_0_2_945), .ZN(n_0_2_944));
   AOI21_X1 i_0_2_985 (.A(n_0_2_948), .B1(n_0_2_949), .B2(n_0_2_946), .ZN(
      n_0_2_945));
   XNOR2_X1 i_0_2_986 (.A(n_0_2_1015), .B(n_0_2_947), .ZN(n_0_2_946));
   OAI211_X1 i_0_2_987 (.A(n_0_2_1018), .B(n_0_2_1010), .C1(n_0_2_1418), 
      .C2(n_0_2_1019), .ZN(n_0_2_947));
   NOR2_X1 i_0_2_988 (.A1(n_0_2_1440), .A2(n_0_2_950), .ZN(n_0_2_948));
   NAND2_X1 i_0_2_989 (.A1(n_0_2_1440), .A2(n_0_2_950), .ZN(n_0_2_949));
   AOI21_X1 i_0_2_990 (.A(n_0_2_953), .B1(n_0_2_954), .B2(n_0_2_951), .ZN(
      n_0_2_950));
   XOR2_X1 i_0_2_991 (.A(n_0_2_1020), .B(n_0_2_952), .Z(n_0_2_951));
   AOI211_X1 i_0_2_992 (.A(n_0_2_1022), .B(n_0_2_1009), .C1(n_0_2_1417), 
      .C2(n_0_2_1024), .ZN(n_0_2_952));
   NOR2_X1 i_0_2_993 (.A1(n_0_2_1418), .A2(n_0_2_955), .ZN(n_0_2_953));
   NAND2_X1 i_0_2_994 (.A1(n_0_2_1418), .A2(n_0_2_955), .ZN(n_0_2_954));
   AOI21_X1 i_0_2_995 (.A(n_0_2_958), .B1(n_0_2_959), .B2(n_0_2_956), .ZN(
      n_0_2_955));
   XOR2_X1 i_0_2_996 (.A(n_0_2_1025), .B(n_0_2_957), .Z(n_0_2_956));
   AOI211_X1 i_0_2_997 (.A(n_0_2_1030), .B(n_0_2_1009), .C1(n_0_2_453), .C2(
      n_0_2_1031), .ZN(n_0_2_957));
   NOR2_X1 i_0_2_998 (.A1(n_0_2_1417), .A2(n_0_2_960), .ZN(n_0_2_958));
   NAND2_X1 i_0_2_999 (.A1(n_0_2_1417), .A2(n_0_2_960), .ZN(n_0_2_959));
   AOI21_X1 i_0_2_1000 (.A(n_0_2_964), .B1(n_0_2_965), .B2(n_0_2_961), .ZN(
      n_0_2_960));
   XOR2_X1 i_0_2_1001 (.A(n_0_2_1032), .B(n_0_2_962), .Z(n_0_2_961));
   NAND3_X1 i_0_2_1002 (.A1(n_0_2_1035), .A2(n_0_2_1034), .A3(n_0_2_1010), 
      .ZN(n_0_2_962));
   INV_X1 i_0_2_1003 (.A(n_0_2_964), .ZN(n_0_2_963));
   NOR2_X1 i_0_2_1004 (.A1(n_0_2_1415), .A2(n_0_2_966), .ZN(n_0_2_964));
   NAND2_X1 i_0_2_1005 (.A1(n_0_2_1415), .A2(n_0_2_966), .ZN(n_0_2_965));
   AOI21_X1 i_0_2_1006 (.A(n_0_2_969), .B1(n_0_2_970), .B2(n_0_2_967), .ZN(
      n_0_2_966));
   XNOR2_X1 i_0_2_1007 (.A(n_0_2_1037), .B(n_0_2_968), .ZN(n_0_2_967));
   NAND3_X1 i_0_2_1008 (.A1(n_0_2_1040), .A2(n_0_2_1039), .A3(n_0_2_1010), 
      .ZN(n_0_2_968));
   NOR2_X1 i_0_2_1009 (.A1(n_0_2_1413), .A2(n_0_2_971), .ZN(n_0_2_969));
   NAND2_X1 i_0_2_1010 (.A1(n_0_2_1413), .A2(n_0_2_971), .ZN(n_0_2_970));
   AOI21_X1 i_0_2_1011 (.A(n_0_2_975), .B1(n_0_2_976), .B2(n_0_2_972), .ZN(
      n_0_2_971));
   XOR2_X1 i_0_2_1012 (.A(n_0_2_1042), .B(n_0_2_973), .Z(n_0_2_972));
   OAI211_X1 i_0_2_1013 (.A(n_0_2_1046), .B(n_0_2_1010), .C1(n_0_2_209), 
      .C2(n_0_2_1047), .ZN(n_0_2_973));
   INV_X1 i_0_2_1014 (.A(n_0_2_975), .ZN(n_0_2_974));
   NOR2_X1 i_0_2_1015 (.A1(n_0_2_1410), .A2(n_0_2_977), .ZN(n_0_2_975));
   NAND2_X1 i_0_2_1016 (.A1(n_0_2_1410), .A2(n_0_2_977), .ZN(n_0_2_976));
   AOI21_X1 i_0_2_1017 (.A(n_0_2_981), .B1(n_0_2_982), .B2(n_0_2_978), .ZN(
      n_0_2_977));
   XOR2_X1 i_0_2_1018 (.A(n_0_2_1048), .B(n_0_2_979), .Z(n_0_2_978));
   NAND3_X1 i_0_2_1019 (.A1(n_0_2_1051), .A2(n_0_2_1050), .A3(n_0_2_1010), 
      .ZN(n_0_2_979));
   INV_X1 i_0_2_1020 (.A(n_0_2_981), .ZN(n_0_2_980));
   NOR2_X1 i_0_2_1021 (.A1(n_0_2_1408), .A2(n_0_2_983), .ZN(n_0_2_981));
   NAND2_X1 i_0_2_1022 (.A1(n_0_2_1408), .A2(n_0_2_983), .ZN(n_0_2_982));
   AOI21_X1 i_0_2_1023 (.A(n_0_2_986), .B1(n_0_2_987), .B2(n_0_2_984), .ZN(
      n_0_2_983));
   XNOR2_X1 i_0_2_1024 (.A(n_0_2_1053), .B(n_0_2_985), .ZN(n_0_2_984));
   OAI211_X1 i_0_2_1025 (.A(n_0_2_1056), .B(n_0_2_1010), .C1(n_0_2_1403), 
      .C2(n_0_2_1057), .ZN(n_0_2_985));
   NOR2_X1 i_0_2_1026 (.A1(n_0_2_1406), .A2(n_0_2_988), .ZN(n_0_2_986));
   NAND2_X1 i_0_2_1027 (.A1(n_0_2_1406), .A2(n_0_2_988), .ZN(n_0_2_987));
   AOI21_X1 i_0_2_1028 (.A(n_0_2_992), .B1(n_0_2_993), .B2(n_0_2_989), .ZN(
      n_0_2_988));
   XOR2_X1 i_0_2_1029 (.A(n_0_2_1058), .B(n_0_2_990), .Z(n_0_2_989));
   AOI211_X1 i_0_2_1030 (.A(n_0_2_1061), .B(n_0_2_1009), .C1(n_0_2_54), .C2(
      n_0_2_1062), .ZN(n_0_2_990));
   INV_X1 i_0_2_1031 (.A(n_0_2_992), .ZN(n_0_2_991));
   NOR2_X1 i_0_2_1032 (.A1(n_0_2_1403), .A2(n_0_2_994), .ZN(n_0_2_992));
   NAND2_X1 i_0_2_1033 (.A1(n_0_2_1403), .A2(n_0_2_994), .ZN(n_0_2_993));
   AOI22_X1 i_0_2_1034 (.A1(n_0_2_54), .A2(n_0_2_999), .B1(n_0_2_998), .B2(
      n_0_2_995), .ZN(n_0_2_994));
   XOR2_X1 i_0_2_1035 (.A(n_0_2_1063), .B(n_0_2_996), .Z(n_0_2_995));
   NAND3_X1 i_0_2_1036 (.A1(n_0_2_1066), .A2(n_0_2_1065), .A3(n_0_2_1010), 
      .ZN(n_0_2_996));
   NAND2_X1 i_0_2_1037 (.A1(n_0_2_54), .A2(n_0_2_999), .ZN(n_0_2_997));
   OR2_X1 i_0_2_1038 (.A1(n_0_2_54), .A2(n_0_2_999), .ZN(n_0_2_998));
   AOI21_X1 i_0_2_1039 (.A(n_0_2_1002), .B1(n_0_2_1003), .B2(n_0_2_1000), 
      .ZN(n_0_2_999));
   XNOR2_X1 i_0_2_1040 (.A(n_0_2_1068), .B(n_0_2_1001), .ZN(n_0_2_1000));
   NAND2_X1 i_0_2_1041 (.A1(in_b[0]), .A2(n_0_2_1010), .ZN(n_0_2_1001));
   NOR2_X1 i_0_2_1042 (.A1(n_0_2_1367), .A2(n_0_2_1004), .ZN(n_0_2_1002));
   OAI21_X1 i_0_2_1043 (.A(n_0_2_49), .B1(n_0_2_1405), .B2(n_0_2_1004), .ZN(
      n_0_2_1003));
   XNOR2_X1 i_0_2_1044 (.A(n_0_2_1446), .B(n_0_2_1005), .ZN(n_0_2_1004));
   AOI21_X1 i_0_2_1045 (.A(n_0_2_1452), .B1(n_0_2_1445), .B2(n_0_2_1006), 
      .ZN(n_0_2_1005));
   OAI21_X1 i_0_2_1046 (.A(in_a[63]), .B1(in_a[1]), .B2(n_0_2_1393), .ZN(
      n_0_2_1006));
   INV_X1 i_0_2_1047 (.A(n_0_2_1008), .ZN(n_0_2_1007));
   AOI21_X1 i_0_2_1048 (.A(n_0_2_1011), .B1(n_0_2_1013), .B2(n_0_2_1010), 
      .ZN(n_0_2_1008));
   NOR2_X1 i_0_2_1049 (.A1(n_0_2_1395), .A2(n_0_2_1009), .ZN(quotient[11]));
   INV_X1 i_0_2_1050 (.A(n_0_2_1010), .ZN(n_0_2_1009));
   AOI221_X1 i_0_2_1051 (.A(n_0_2_1420), .B1(n_0_2_1440), .B2(n_0_2_1014), 
      .C1(n_0_2_1013), .C2(n_0_2_1011), .ZN(n_0_2_1010));
   INV_X1 i_0_2_1052 (.A(n_0_2_1012), .ZN(n_0_2_1011));
   AOI21_X1 i_0_2_1053 (.A(n_0_2_1074), .B1(n_0_2_1370), .B2(n_0_2_1072), 
      .ZN(n_0_2_1012));
   OR2_X1 i_0_2_1054 (.A1(n_0_2_1440), .A2(n_0_2_1014), .ZN(n_0_2_1013));
   AOI21_X1 i_0_2_1055 (.A(n_0_2_1017), .B1(n_0_2_1018), .B2(n_0_2_1015), 
      .ZN(n_0_2_1014));
   XNOR2_X1 i_0_2_1056 (.A(n_0_2_1077), .B(n_0_2_1016), .ZN(n_0_2_1015));
   NAND3_X1 i_0_2_1057 (.A1(n_0_2_1080), .A2(n_0_2_1079), .A3(n_0_2_1070), 
      .ZN(n_0_2_1016));
   NOR2_X1 i_0_2_1058 (.A1(n_0_2_1418), .A2(n_0_2_1019), .ZN(n_0_2_1017));
   NAND2_X1 i_0_2_1059 (.A1(n_0_2_1418), .A2(n_0_2_1019), .ZN(n_0_2_1018));
   AOI21_X1 i_0_2_1060 (.A(n_0_2_1022), .B1(n_0_2_1023), .B2(n_0_2_1020), 
      .ZN(n_0_2_1019));
   AOI22_X1 i_0_2_1061 (.A1(n_0_2_1121), .A2(n_0_2_1071), .B1(n_0_2_1070), 
      .B2(n_0_2_1021), .ZN(n_0_2_1020));
   XOR2_X1 i_0_2_1062 (.A(n_0_2_1120), .B(n_0_2_1082), .Z(n_0_2_1021));
   NOR2_X1 i_0_2_1063 (.A1(n_0_2_1417), .A2(n_0_2_1024), .ZN(n_0_2_1022));
   NAND2_X1 i_0_2_1064 (.A1(n_0_2_1417), .A2(n_0_2_1024), .ZN(n_0_2_1023));
   AOI22_X1 i_0_2_1065 (.A1(n_0_2_453), .A2(n_0_2_1031), .B1(n_0_2_1029), 
      .B2(n_0_2_1025), .ZN(n_0_2_1024));
   OAI21_X1 i_0_2_1066 (.A(n_0_2_1026), .B1(n_0_2_1118), .B2(n_0_2_1070), 
      .ZN(n_0_2_1025));
   NAND2_X1 i_0_2_1067 (.A1(n_0_2_1070), .A2(n_0_2_1027), .ZN(n_0_2_1026));
   XNOR2_X1 i_0_2_1068 (.A(n_0_2_1083), .B(n_0_2_1028), .ZN(n_0_2_1027));
   OAI21_X1 i_0_2_1069 (.A(n_0_2_1116), .B1(n_0_2_1413), .B2(n_0_2_1118), 
      .ZN(n_0_2_1028));
   INV_X1 i_0_2_1070 (.A(n_0_2_1030), .ZN(n_0_2_1029));
   NOR2_X1 i_0_2_1071 (.A1(n_0_2_453), .A2(n_0_2_1031), .ZN(n_0_2_1030));
   AOI22_X1 i_0_2_1072 (.A1(n_0_2_1413), .A2(n_0_2_1036), .B1(n_0_2_1034), 
      .B2(n_0_2_1032), .ZN(n_0_2_1031));
   AOI22_X1 i_0_2_1073 (.A1(n_0_2_1114), .A2(n_0_2_1071), .B1(n_0_2_1070), 
      .B2(n_0_2_1033), .ZN(n_0_2_1032));
   XOR2_X1 i_0_2_1074 (.A(n_0_2_1112), .B(n_0_2_1085), .Z(n_0_2_1033));
   OR2_X1 i_0_2_1075 (.A1(n_0_2_1413), .A2(n_0_2_1036), .ZN(n_0_2_1034));
   NAND2_X1 i_0_2_1076 (.A1(n_0_2_1413), .A2(n_0_2_1036), .ZN(n_0_2_1035));
   AOI22_X1 i_0_2_1077 (.A1(n_0_2_281), .A2(n_0_2_1041), .B1(n_0_2_1040), 
      .B2(n_0_2_1037), .ZN(n_0_2_1036));
   AOI22_X1 i_0_2_1078 (.A1(n_0_2_1110), .A2(n_0_2_1071), .B1(n_0_2_1070), 
      .B2(n_0_2_1038), .ZN(n_0_2_1037));
   XOR2_X1 i_0_2_1079 (.A(n_0_2_1109), .B(n_0_2_1086), .Z(n_0_2_1038));
   NAND2_X1 i_0_2_1080 (.A1(n_0_2_281), .A2(n_0_2_1041), .ZN(n_0_2_1039));
   OR2_X1 i_0_2_1081 (.A1(n_0_2_281), .A2(n_0_2_1041), .ZN(n_0_2_1040));
   AOI21_X1 i_0_2_1082 (.A(n_0_2_1045), .B1(n_0_2_1046), .B2(n_0_2_1042), 
      .ZN(n_0_2_1041));
   AOI22_X1 i_0_2_1083 (.A1(n_0_2_1107), .A2(n_0_2_1071), .B1(n_0_2_1070), 
      .B2(n_0_2_1043), .ZN(n_0_2_1042));
   XOR2_X1 i_0_2_1084 (.A(n_0_2_1088), .B(n_0_2_1087), .Z(n_0_2_1043));
   NOR2_X1 i_0_2_1085 (.A1(n_0_2_209), .A2(n_0_2_1047), .ZN(n_0_2_1045));
   NAND2_X1 i_0_2_1086 (.A1(n_0_2_209), .A2(n_0_2_1047), .ZN(n_0_2_1046));
   AOI22_X1 i_0_2_1087 (.A1(n_0_2_1406), .A2(n_0_2_1052), .B1(n_0_2_1051), 
      .B2(n_0_2_1048), .ZN(n_0_2_1047));
   AOI22_X1 i_0_2_1088 (.A1(n_0_2_1105), .A2(n_0_2_1071), .B1(n_0_2_1070), 
      .B2(n_0_2_1049), .ZN(n_0_2_1048));
   XNOR2_X1 i_0_2_1089 (.A(n_0_2_1103), .B(n_0_2_1089), .ZN(n_0_2_1049));
   NAND2_X1 i_0_2_1090 (.A1(n_0_2_1406), .A2(n_0_2_1052), .ZN(n_0_2_1050));
   OR2_X1 i_0_2_1091 (.A1(n_0_2_1406), .A2(n_0_2_1052), .ZN(n_0_2_1051));
   AOI21_X1 i_0_2_1092 (.A(n_0_2_1055), .B1(n_0_2_1056), .B2(n_0_2_1053), 
      .ZN(n_0_2_1052));
   XNOR2_X1 i_0_2_1093 (.A(n_0_2_1090), .B(n_0_2_1054), .ZN(n_0_2_1053));
   OAI211_X1 i_0_2_1094 (.A(n_0_2_1094), .B(n_0_2_1070), .C1(n_0_2_1400), 
      .C2(n_0_2_1095), .ZN(n_0_2_1054));
   NOR2_X1 i_0_2_1095 (.A1(n_0_2_1403), .A2(n_0_2_1057), .ZN(n_0_2_1055));
   NAND2_X1 i_0_2_1096 (.A1(n_0_2_1403), .A2(n_0_2_1057), .ZN(n_0_2_1056));
   AOI22_X1 i_0_2_1097 (.A1(n_0_2_54), .A2(n_0_2_1062), .B1(n_0_2_1060), 
      .B2(n_0_2_1058), .ZN(n_0_2_1057));
   XNOR2_X1 i_0_2_1098 (.A(n_0_2_1098), .B(n_0_2_1059), .ZN(n_0_2_1058));
   NAND3_X1 i_0_2_1099 (.A1(n_0_2_1100), .A2(n_0_2_1097), .A3(n_0_2_1070), 
      .ZN(n_0_2_1059));
   INV_X1 i_0_2_1100 (.A(n_0_2_1061), .ZN(n_0_2_1060));
   NOR2_X1 i_0_2_1101 (.A1(n_0_2_54), .A2(n_0_2_1062), .ZN(n_0_2_1061));
   AOI22_X1 i_0_2_1102 (.A1(n_0_2_1366), .A2(n_0_2_1068), .B1(n_0_2_1066), 
      .B2(n_0_2_1063), .ZN(n_0_2_1062));
   XOR2_X1 i_0_2_1103 (.A(n_0_2_1101), .B(n_0_2_1064), .Z(n_0_2_1063));
   NAND2_X1 i_0_2_1104 (.A1(in_b[0]), .A2(n_0_2_1070), .ZN(n_0_2_1064));
   NAND2_X1 i_0_2_1105 (.A1(n_0_2_1366), .A2(n_0_2_1068), .ZN(n_0_2_1065));
   INV_X1 i_0_2_1106 (.A(n_0_2_1067), .ZN(n_0_2_1066));
   AOI21_X1 i_0_2_1107 (.A(n_0_2_1398), .B1(in_b[0]), .B2(n_0_2_1068), .ZN(
      n_0_2_1067));
   XNOR2_X1 i_0_2_1108 (.A(in_a[4]), .B(n_0_2_1069), .ZN(n_0_2_1068));
   AND2_X1 i_0_2_1109 (.A1(in_a[63]), .A2(n_0_2_1391), .ZN(n_0_2_1069));
   NOR2_X1 i_0_2_1110 (.A1(n_0_2_1395), .A2(n_0_2_1071), .ZN(quotient[12]));
   INV_X1 i_0_2_1111 (.A(n_0_2_1071), .ZN(n_0_2_1070));
   NAND2_X1 i_0_2_1112 (.A1(n_0_2_1073), .A2(n_0_2_1072), .ZN(n_0_2_1071));
   AOI21_X1 i_0_2_1113 (.A(n_0_2_1419), .B1(n_0_2_1418), .B2(n_0_2_1076), 
      .ZN(n_0_2_1072));
   OAI21_X1 i_0_2_1114 (.A(n_0_2_1074), .B1(n_0_2_1418), .B2(n_0_2_1076), 
      .ZN(n_0_2_1073));
   INV_X1 i_0_2_1115 (.A(n_0_2_1075), .ZN(n_0_2_1074));
   AOI22_X1 i_0_2_1116 (.A1(n_0_2_1370), .A2(n_0_2_1129), .B1(n_0_2_1370), 
      .B2(n_0_2_1125), .ZN(n_0_2_1075));
   AOI22_X1 i_0_2_1117 (.A1(n_0_2_458), .A2(n_0_2_1081), .B1(n_0_2_1079), 
      .B2(n_0_2_1077), .ZN(n_0_2_1076));
   XNOR2_X1 i_0_2_1118 (.A(n_0_2_1130), .B(n_0_2_1078), .ZN(n_0_2_1077));
   NAND3_X1 i_0_2_1119 (.A1(n_0_2_1132), .A2(n_0_2_1127), .A3(n_0_2_1123), 
      .ZN(n_0_2_1078));
   OR2_X1 i_0_2_1120 (.A1(n_0_2_458), .A2(n_0_2_1081), .ZN(n_0_2_1079));
   NAND2_X1 i_0_2_1121 (.A1(n_0_2_458), .A2(n_0_2_1081), .ZN(n_0_2_1080));
   AOI22_X1 i_0_2_1122 (.A1(n_0_2_1415), .A2(n_0_2_1121), .B1(n_0_2_1120), 
      .B2(n_0_2_1082), .ZN(n_0_2_1081));
   AOI22_X1 i_0_2_1123 (.A1(n_0_2_363), .A2(n_0_2_1117), .B1(n_0_2_1116), 
      .B2(n_0_2_1083), .ZN(n_0_2_1082));
   AOI22_X1 i_0_2_1124 (.A1(n_0_2_1410), .A2(n_0_2_1113), .B1(n_0_2_1112), 
      .B2(n_0_2_1084), .ZN(n_0_2_1083));
   INV_X1 i_0_2_1125 (.A(n_0_2_1085), .ZN(n_0_2_1084));
   AOI22_X1 i_0_2_1126 (.A1(n_0_2_1408), .A2(n_0_2_1110), .B1(n_0_2_1109), 
      .B2(n_0_2_1086), .ZN(n_0_2_1085));
   AOI22_X1 i_0_2_1127 (.A1(n_0_2_147), .A2(n_0_2_1107), .B1(n_0_2_1088), 
      .B2(n_0_2_1087), .ZN(n_0_2_1086));
   XNOR2_X1 i_0_2_1128 (.A(n_0_2_1406), .B(n_0_2_1107), .ZN(n_0_2_1087));
   AOI22_X1 i_0_2_1129 (.A1(n_0_2_1403), .A2(n_0_2_1104), .B1(n_0_2_1103), 
      .B2(n_0_2_1089), .ZN(n_0_2_1088));
   AOI21_X1 i_0_2_1130 (.A(n_0_2_1093), .B1(n_0_2_1094), .B2(n_0_2_1090), 
      .ZN(n_0_2_1089));
   XNOR2_X1 i_0_2_1131 (.A(n_0_2_1166), .B(n_0_2_1092), .ZN(n_0_2_1090));
   NAND3_X1 i_0_2_1132 (.A1(n_0_2_1168), .A2(n_0_2_1165), .A3(n_0_2_1123), 
      .ZN(n_0_2_1092));
   NOR2_X1 i_0_2_1133 (.A1(n_0_2_1400), .A2(n_0_2_1095), .ZN(n_0_2_1093));
   NAND2_X1 i_0_2_1134 (.A1(n_0_2_1400), .A2(n_0_2_1095), .ZN(n_0_2_1094));
   AOI21_X1 i_0_2_1135 (.A(n_0_2_1096), .B1(n_0_2_1100), .B2(n_0_2_1098), 
      .ZN(n_0_2_1095));
   INV_X1 i_0_2_1136 (.A(n_0_2_1097), .ZN(n_0_2_1096));
   AOI21_X1 i_0_2_1137 (.A(n_0_2_1397), .B1(n_0_2_49), .B2(n_0_2_1101), .ZN(
      n_0_2_1097));
   XNOR2_X1 i_0_2_1138 (.A(n_0_2_1169), .B(n_0_2_1099), .ZN(n_0_2_1098));
   NAND2_X1 i_0_2_1139 (.A1(in_b[0]), .A2(n_0_2_1123), .ZN(n_0_2_1099));
   OR2_X1 i_0_2_1140 (.A1(n_0_2_1367), .A2(n_0_2_1101), .ZN(n_0_2_1100));
   XNOR2_X1 i_0_2_1141 (.A(n_0_2_1447), .B(n_0_2_1102), .ZN(n_0_2_1101));
   NOR2_X1 i_0_2_1142 (.A1(n_0_2_1452), .A2(n_0_2_1390), .ZN(n_0_2_1102));
   AOI22_X1 i_0_2_1143 (.A1(n_0_2_1403), .A2(n_0_2_1104), .B1(n_0_2_96), 
      .B2(n_0_2_1105), .ZN(n_0_2_1103));
   INV_X1 i_0_2_1144 (.A(n_0_2_1105), .ZN(n_0_2_1104));
   XNOR2_X1 i_0_2_1145 (.A(n_0_2_1159), .B(n_0_2_1106), .ZN(n_0_2_1105));
   AOI211_X1 i_0_2_1146 (.A(n_0_2_1162), .B(n_0_2_1124), .C1(n_0_2_1400), 
      .C2(n_0_2_1163), .ZN(n_0_2_1106));
   XOR2_X1 i_0_2_1147 (.A(n_0_2_1154), .B(n_0_2_1108), .Z(n_0_2_1107));
   AOI211_X1 i_0_2_1148 (.A(n_0_2_1157), .B(n_0_2_1124), .C1(n_0_2_96), .C2(
      n_0_2_1158), .ZN(n_0_2_1108));
   XNOR2_X1 i_0_2_1149 (.A(n_0_2_209), .B(n_0_2_1110), .ZN(n_0_2_1109));
   XOR2_X1 i_0_2_1150 (.A(n_0_2_1149), .B(n_0_2_1111), .Z(n_0_2_1110));
   AOI211_X1 i_0_2_1151 (.A(n_0_2_1152), .B(n_0_2_1124), .C1(n_0_2_1406), 
      .C2(n_0_2_1153), .ZN(n_0_2_1111));
   AOI22_X1 i_0_2_1152 (.A1(n_0_2_1410), .A2(n_0_2_1113), .B1(n_0_2_281), 
      .B2(n_0_2_1114), .ZN(n_0_2_1112));
   INV_X1 i_0_2_1153 (.A(n_0_2_1114), .ZN(n_0_2_1113));
   XNOR2_X1 i_0_2_1154 (.A(n_0_2_1144), .B(n_0_2_1115), .ZN(n_0_2_1114));
   NAND3_X1 i_0_2_1155 (.A1(n_0_2_1147), .A2(n_0_2_1146), .A3(n_0_2_1123), 
      .ZN(n_0_2_1115));
   NAND2_X1 i_0_2_1156 (.A1(n_0_2_1413), .A2(n_0_2_1118), .ZN(n_0_2_1116));
   INV_X1 i_0_2_1157 (.A(n_0_2_1118), .ZN(n_0_2_1117));
   XNOR2_X1 i_0_2_1158 (.A(n_0_2_1139), .B(n_0_2_1119), .ZN(n_0_2_1118));
   AOI211_X1 i_0_2_1159 (.A(n_0_2_1142), .B(n_0_2_1124), .C1(n_0_2_1410), 
      .C2(n_0_2_1143), .ZN(n_0_2_1119));
   XNOR2_X1 i_0_2_1160 (.A(n_0_2_453), .B(n_0_2_1121), .ZN(n_0_2_1120));
   XNOR2_X1 i_0_2_1161 (.A(n_0_2_1134), .B(n_0_2_1122), .ZN(n_0_2_1121));
   NAND3_X1 i_0_2_1162 (.A1(n_0_2_1137), .A2(n_0_2_1136), .A3(n_0_2_1123), 
      .ZN(n_0_2_1122));
   NOR2_X1 i_0_2_1163 (.A1(n_0_2_1395), .A2(n_0_2_1124), .ZN(quotient[13]));
   INV_X1 i_0_2_1164 (.A(n_0_2_1124), .ZN(n_0_2_1123));
   OAI21_X1 i_0_2_1165 (.A(n_0_2_1125), .B1(n_0_2_458), .B2(n_0_2_1176), 
      .ZN(n_0_2_1124));
   NOR3_X1 i_0_2_1166 (.A1(n_0_2_1419), .A2(n_0_2_1418), .A3(n_0_2_1126), 
      .ZN(n_0_2_1125));
   AOI221_X1 i_0_2_1167 (.A(n_0_2_1128), .B1(n_0_2_453), .B2(n_0_2_1133), 
      .C1(n_0_2_1132), .C2(n_0_2_1130), .ZN(n_0_2_1126));
   NAND2_X1 i_0_2_1168 (.A1(n_0_2_453), .A2(n_0_2_1133), .ZN(n_0_2_1127));
   AOI21_X1 i_0_2_1169 (.A(n_0_2_1417), .B1(n_0_2_1370), .B2(n_0_2_1129), 
      .ZN(n_0_2_1128));
   NAND2_X1 i_0_2_1170 (.A1(n_0_2_1178), .A2(n_0_2_1173), .ZN(n_0_2_1129));
   XNOR2_X1 i_0_2_1171 (.A(n_0_2_1180), .B(n_0_2_1131), .ZN(n_0_2_1130));
   NAND3_X1 i_0_2_1172 (.A1(n_0_2_1182), .A2(n_0_2_1179), .A3(n_0_2_1172), 
      .ZN(n_0_2_1131));
   OR2_X1 i_0_2_1173 (.A1(n_0_2_453), .A2(n_0_2_1133), .ZN(n_0_2_1132));
   AOI22_X1 i_0_2_1174 (.A1(n_0_2_1413), .A2(n_0_2_1138), .B1(n_0_2_1137), 
      .B2(n_0_2_1134), .ZN(n_0_2_1133));
   XNOR2_X1 i_0_2_1175 (.A(n_0_2_1184), .B(n_0_2_1135), .ZN(n_0_2_1134));
   AND3_X1 i_0_2_1176 (.A1(n_0_2_1188), .A2(n_0_2_1186), .A3(n_0_2_1172), 
      .ZN(n_0_2_1135));
   NAND2_X1 i_0_2_1177 (.A1(n_0_2_1413), .A2(n_0_2_1138), .ZN(n_0_2_1136));
   OR2_X1 i_0_2_1178 (.A1(n_0_2_1413), .A2(n_0_2_1138), .ZN(n_0_2_1137));
   OAI21_X1 i_0_2_1179 (.A(n_0_2_1141), .B1(n_0_2_1142), .B2(n_0_2_1139), 
      .ZN(n_0_2_1138));
   XNOR2_X1 i_0_2_1180 (.A(n_0_2_1191), .B(n_0_2_1140), .ZN(n_0_2_1139));
   OAI211_X1 i_0_2_1181 (.A(n_0_2_1194), .B(n_0_2_1172), .C1(n_0_2_1408), 
      .C2(n_0_2_1195), .ZN(n_0_2_1140));
   NAND2_X1 i_0_2_1182 (.A1(n_0_2_1410), .A2(n_0_2_1143), .ZN(n_0_2_1141));
   NOR2_X1 i_0_2_1183 (.A1(n_0_2_1410), .A2(n_0_2_1143), .ZN(n_0_2_1142));
   AOI22_X1 i_0_2_1184 (.A1(n_0_2_209), .A2(n_0_2_1148), .B1(n_0_2_1146), 
      .B2(n_0_2_1144), .ZN(n_0_2_1143));
   XNOR2_X1 i_0_2_1185 (.A(n_0_2_1198), .B(n_0_2_1145), .ZN(n_0_2_1144));
   OAI211_X1 i_0_2_1186 (.A(n_0_2_1201), .B(n_0_2_1172), .C1(n_0_2_1406), 
      .C2(n_0_2_1202), .ZN(n_0_2_1145));
   OR2_X1 i_0_2_1187 (.A1(n_0_2_209), .A2(n_0_2_1148), .ZN(n_0_2_1146));
   NAND2_X1 i_0_2_1188 (.A1(n_0_2_209), .A2(n_0_2_1148), .ZN(n_0_2_1147));
   AOI22_X1 i_0_2_1189 (.A1(n_0_2_1406), .A2(n_0_2_1153), .B1(n_0_2_1151), 
      .B2(n_0_2_1149), .ZN(n_0_2_1148));
   XOR2_X1 i_0_2_1190 (.A(n_0_2_1203), .B(n_0_2_1150), .Z(n_0_2_1149));
   NAND3_X1 i_0_2_1191 (.A1(n_0_2_1206), .A2(n_0_2_1205), .A3(n_0_2_1172), 
      .ZN(n_0_2_1150));
   INV_X1 i_0_2_1192 (.A(n_0_2_1152), .ZN(n_0_2_1151));
   NOR2_X1 i_0_2_1193 (.A1(n_0_2_1406), .A2(n_0_2_1153), .ZN(n_0_2_1152));
   AOI22_X1 i_0_2_1194 (.A1(n_0_2_96), .A2(n_0_2_1158), .B1(n_0_2_1156), 
      .B2(n_0_2_1154), .ZN(n_0_2_1153));
   XNOR2_X1 i_0_2_1195 (.A(n_0_2_1208), .B(n_0_2_1155), .ZN(n_0_2_1154));
   AND3_X1 i_0_2_1196 (.A1(n_0_2_1212), .A2(n_0_2_1210), .A3(n_0_2_1172), 
      .ZN(n_0_2_1155));
   INV_X1 i_0_2_1197 (.A(n_0_2_1157), .ZN(n_0_2_1156));
   NOR2_X1 i_0_2_1198 (.A1(n_0_2_96), .A2(n_0_2_1158), .ZN(n_0_2_1157));
   AOI22_X1 i_0_2_1199 (.A1(n_0_2_1400), .A2(n_0_2_1163), .B1(n_0_2_1161), 
      .B2(n_0_2_1159), .ZN(n_0_2_1158));
   XNOR2_X1 i_0_2_1200 (.A(n_0_2_1215), .B(n_0_2_1160), .ZN(n_0_2_1159));
   OAI211_X1 i_0_2_1201 (.A(n_0_2_1217), .B(n_0_2_1172), .C1(n_0_2_1367), 
      .C2(n_0_2_1218), .ZN(n_0_2_1160));
   INV_X1 i_0_2_1202 (.A(n_0_2_1162), .ZN(n_0_2_1161));
   NOR2_X1 i_0_2_1203 (.A1(n_0_2_1400), .A2(n_0_2_1163), .ZN(n_0_2_1162));
   AOI21_X1 i_0_2_1204 (.A(n_0_2_1164), .B1(n_0_2_1168), .B2(n_0_2_1166), 
      .ZN(n_0_2_1163));
   INV_X1 i_0_2_1205 (.A(n_0_2_1165), .ZN(n_0_2_1164));
   AOI21_X1 i_0_2_1206 (.A(n_0_2_1397), .B1(n_0_2_49), .B2(n_0_2_1169), .ZN(
      n_0_2_1165));
   XNOR2_X1 i_0_2_1207 (.A(n_0_2_1218), .B(n_0_2_1167), .ZN(n_0_2_1166));
   NAND2_X1 i_0_2_1208 (.A1(in_b[0]), .A2(n_0_2_1172), .ZN(n_0_2_1167));
   NAND2_X1 i_0_2_1209 (.A1(n_0_2_1366), .A2(n_0_2_1170), .ZN(n_0_2_1168));
   INV_X1 i_0_2_1210 (.A(n_0_2_1170), .ZN(n_0_2_1169));
   XNOR2_X1 i_0_2_1211 (.A(in_a[6]), .B(n_0_2_1171), .ZN(n_0_2_1170));
   AOI21_X1 i_0_2_1212 (.A(n_0_2_1452), .B1(n_0_2_1447), .B2(n_0_2_1390), 
      .ZN(n_0_2_1171));
   AND2_X1 i_0_2_1213 (.A1(n_0_2_1394), .A2(n_0_2_1172), .ZN(quotient[14]));
   AOI21_X1 i_0_2_1214 (.A(n_0_2_1173), .B1(n_0_2_1415), .B2(n_0_2_1223), 
      .ZN(n_0_2_1172));
   INV_X1 i_0_2_1215 (.A(n_0_2_1174), .ZN(n_0_2_1173));
   AOI21_X1 i_0_2_1216 (.A(n_0_2_1416), .B1(n_0_2_1179), .B2(n_0_2_1175), 
      .ZN(n_0_2_1174));
   AOI22_X1 i_0_2_1217 (.A1(n_0_2_1182), .A2(n_0_2_1180), .B1(n_0_2_453), 
      .B2(n_0_2_1176), .ZN(n_0_2_1175));
   NAND2_X1 i_0_2_1218 (.A1(n_0_2_1370), .A2(n_0_2_1177), .ZN(n_0_2_1176));
   INV_X1 i_0_2_1219 (.A(n_0_2_1178), .ZN(n_0_2_1177));
   AOI211_X1 i_0_2_1220 (.A(n_0_2_1286), .B(n_0_2_1256), .C1(n_0_2_1414), 
      .C2(n_0_2_1221), .ZN(n_0_2_1178));
   OR2_X1 i_0_2_1221 (.A1(n_0_2_1413), .A2(n_0_2_1183), .ZN(n_0_2_1179));
   XOR2_X1 i_0_2_1222 (.A(n_0_2_1226), .B(n_0_2_1181), .Z(n_0_2_1180));
   AND3_X1 i_0_2_1223 (.A1(n_0_2_1228), .A2(n_0_2_1225), .A3(n_0_2_1219), 
      .ZN(n_0_2_1181));
   NAND2_X1 i_0_2_1224 (.A1(n_0_2_1413), .A2(n_0_2_1183), .ZN(n_0_2_1182));
   AOI21_X1 i_0_2_1225 (.A(n_0_2_1187), .B1(n_0_2_1188), .B2(n_0_2_1184), 
      .ZN(n_0_2_1183));
   XOR2_X1 i_0_2_1226 (.A(n_0_2_1230), .B(n_0_2_1185), .Z(n_0_2_1184));
   NAND3_X1 i_0_2_1227 (.A1(n_0_2_1233), .A2(n_0_2_1232), .A3(n_0_2_1219), 
      .ZN(n_0_2_1185));
   INV_X1 i_0_2_1228 (.A(n_0_2_1187), .ZN(n_0_2_1186));
   NOR2_X1 i_0_2_1229 (.A1(n_0_2_1410), .A2(n_0_2_1189), .ZN(n_0_2_1187));
   NAND2_X1 i_0_2_1230 (.A1(n_0_2_1410), .A2(n_0_2_1189), .ZN(n_0_2_1188));
   AOI21_X1 i_0_2_1231 (.A(n_0_2_1193), .B1(n_0_2_1194), .B2(n_0_2_1191), 
      .ZN(n_0_2_1189));
   XOR2_X1 i_0_2_1232 (.A(n_0_2_1235), .B(n_0_2_1192), .Z(n_0_2_1191));
   AND3_X1 i_0_2_1233 (.A1(n_0_2_1238), .A2(n_0_2_1237), .A3(n_0_2_1219), 
      .ZN(n_0_2_1192));
   NOR2_X1 i_0_2_1234 (.A1(n_0_2_1408), .A2(n_0_2_1195), .ZN(n_0_2_1193));
   NAND2_X1 i_0_2_1235 (.A1(n_0_2_1408), .A2(n_0_2_1195), .ZN(n_0_2_1194));
   AOI21_X1 i_0_2_1236 (.A(n_0_2_1200), .B1(n_0_2_1201), .B2(n_0_2_1198), 
      .ZN(n_0_2_1195));
   XNOR2_X1 i_0_2_1237 (.A(n_0_2_1240), .B(n_0_2_1199), .ZN(n_0_2_1198));
   AND3_X1 i_0_2_1238 (.A1(n_0_2_1243), .A2(n_0_2_1242), .A3(n_0_2_1219), 
      .ZN(n_0_2_1199));
   NOR2_X1 i_0_2_1239 (.A1(n_0_2_1406), .A2(n_0_2_1202), .ZN(n_0_2_1200));
   NAND2_X1 i_0_2_1240 (.A1(n_0_2_1406), .A2(n_0_2_1202), .ZN(n_0_2_1201));
   AOI22_X1 i_0_2_1241 (.A1(n_0_2_96), .A2(n_0_2_1207), .B1(n_0_2_1205), 
      .B2(n_0_2_1203), .ZN(n_0_2_1202));
   XNOR2_X1 i_0_2_1242 (.A(n_0_2_1245), .B(n_0_2_1204), .ZN(n_0_2_1203));
   NAND3_X1 i_0_2_1243 (.A1(n_0_2_1250), .A2(n_0_2_1249), .A3(n_0_2_1219), 
      .ZN(n_0_2_1204));
   OR2_X1 i_0_2_1244 (.A1(n_0_2_96), .A2(n_0_2_1207), .ZN(n_0_2_1205));
   NAND2_X1 i_0_2_1245 (.A1(n_0_2_96), .A2(n_0_2_1207), .ZN(n_0_2_1206));
   AOI21_X1 i_0_2_1246 (.A(n_0_2_1211), .B1(n_0_2_1212), .B2(n_0_2_1208), 
      .ZN(n_0_2_1207));
   XNOR2_X1 i_0_2_1247 (.A(n_0_2_1252), .B(n_0_2_1209), .ZN(n_0_2_1208));
   OAI211_X1 i_0_2_1248 (.A(n_0_2_1384), .B(n_0_2_1219), .C1(n_0_2_1385), 
      .C2(n_0_2_1367), .ZN(n_0_2_1209));
   INV_X1 i_0_2_1249 (.A(n_0_2_1211), .ZN(n_0_2_1210));
   NOR2_X1 i_0_2_1250 (.A1(n_0_2_54), .A2(n_0_2_1213), .ZN(n_0_2_1211));
   NAND2_X1 i_0_2_1251 (.A1(n_0_2_54), .A2(n_0_2_1213), .ZN(n_0_2_1212));
   AOI21_X1 i_0_2_1252 (.A(n_0_2_1214), .B1(n_0_2_1217), .B2(n_0_2_1215), 
      .ZN(n_0_2_1213));
   NOR2_X1 i_0_2_1253 (.A1(n_0_2_1367), .A2(n_0_2_1218), .ZN(n_0_2_1214));
   XNOR2_X1 i_0_2_1254 (.A(n_0_2_1386), .B(n_0_2_1216), .ZN(n_0_2_1215));
   NAND2_X1 i_0_2_1255 (.A1(in_b[0]), .A2(n_0_2_1219), .ZN(n_0_2_1216));
   AOI21_X1 i_0_2_1256 (.A(n_0_2_1397), .B1(n_0_2_49), .B2(n_0_2_1218), .ZN(
      n_0_2_1217));
   XNOR2_X1 i_0_2_1257 (.A(in_a[7]), .B(n_0_2_1388), .ZN(n_0_2_1218));
   AND2_X1 i_0_2_1258 (.A1(n_0_2_1394), .A2(n_0_2_1219), .ZN(quotient[15]));
   AOI21_X1 i_0_2_1259 (.A(n_0_2_1220), .B1(n_0_2_1413), .B2(n_0_2_1285), 
      .ZN(n_0_2_1219));
   NAND2_X1 i_0_2_1260 (.A1(n_0_2_1414), .A2(n_0_2_1221), .ZN(n_0_2_1220));
   NAND2_X1 i_0_2_1261 (.A1(n_0_2_1225), .A2(n_0_2_1222), .ZN(n_0_2_1221));
   AOI22_X1 i_0_2_1262 (.A1(n_0_2_1228), .A2(n_0_2_1226), .B1(n_0_2_363), 
      .B2(n_0_2_1224), .ZN(n_0_2_1222));
   INV_X1 i_0_2_1263 (.A(n_0_2_1224), .ZN(n_0_2_1223));
   OAI21_X1 i_0_2_1264 (.A(n_0_2_1370), .B1(n_0_2_1286), .B2(n_0_2_1256), 
      .ZN(n_0_2_1224));
   NAND2_X1 i_0_2_1265 (.A1(n_0_2_281), .A2(n_0_2_1229), .ZN(n_0_2_1225));
   XNOR2_X1 i_0_2_1266 (.A(n_0_2_1259), .B(n_0_2_1227), .ZN(n_0_2_1226));
   NAND3_X1 i_0_2_1267 (.A1(n_0_2_1262), .A2(n_0_2_1261), .A3(n_0_2_1254), 
      .ZN(n_0_2_1227));
   OR2_X1 i_0_2_1268 (.A1(n_0_2_281), .A2(n_0_2_1229), .ZN(n_0_2_1228));
   AOI22_X1 i_0_2_1269 (.A1(n_0_2_1408), .A2(n_0_2_1234), .B1(n_0_2_1232), 
      .B2(n_0_2_1230), .ZN(n_0_2_1229));
   XNOR2_X1 i_0_2_1270 (.A(n_0_2_1264), .B(n_0_2_1231), .ZN(n_0_2_1230));
   OAI211_X1 i_0_2_1271 (.A(n_0_2_1266), .B(n_0_2_1254), .C1(n_0_2_147), 
      .C2(n_0_2_1268), .ZN(n_0_2_1231));
   OR2_X1 i_0_2_1272 (.A1(n_0_2_1408), .A2(n_0_2_1234), .ZN(n_0_2_1232));
   NAND2_X1 i_0_2_1273 (.A1(n_0_2_1408), .A2(n_0_2_1234), .ZN(n_0_2_1233));
   AOI22_X1 i_0_2_1274 (.A1(n_0_2_147), .A2(n_0_2_1239), .B1(n_0_2_1238), 
      .B2(n_0_2_1235), .ZN(n_0_2_1234));
   XOR2_X1 i_0_2_1275 (.A(n_0_2_1269), .B(n_0_2_1236), .Z(n_0_2_1235));
   NAND3_X1 i_0_2_1276 (.A1(n_0_2_1272), .A2(n_0_2_1271), .A3(n_0_2_1254), 
      .ZN(n_0_2_1236));
   NAND2_X1 i_0_2_1277 (.A1(n_0_2_147), .A2(n_0_2_1239), .ZN(n_0_2_1237));
   OR2_X1 i_0_2_1278 (.A1(n_0_2_147), .A2(n_0_2_1239), .ZN(n_0_2_1238));
   AOI22_X1 i_0_2_1279 (.A1(n_0_2_1403), .A2(n_0_2_1244), .B1(n_0_2_1243), 
      .B2(n_0_2_1240), .ZN(n_0_2_1239));
   XOR2_X1 i_0_2_1280 (.A(n_0_2_1274), .B(n_0_2_1241), .Z(n_0_2_1240));
   NAND3_X1 i_0_2_1281 (.A1(n_0_2_1277), .A2(n_0_2_1276), .A3(n_0_2_1254), 
      .ZN(n_0_2_1241));
   NAND2_X1 i_0_2_1282 (.A1(n_0_2_1403), .A2(n_0_2_1244), .ZN(n_0_2_1242));
   OR2_X1 i_0_2_1283 (.A1(n_0_2_1403), .A2(n_0_2_1244), .ZN(n_0_2_1243));
   AOI22_X1 i_0_2_1284 (.A1(n_0_2_54), .A2(n_0_2_1251), .B1(n_0_2_1250), 
      .B2(n_0_2_1245), .ZN(n_0_2_1244));
   XOR2_X1 i_0_2_1285 (.A(n_0_2_1279), .B(n_0_2_1248), .Z(n_0_2_1245));
   OAI211_X1 i_0_2_1286 (.A(n_0_2_1284), .B(n_0_2_1254), .C1(n_0_2_1380), 
      .C2(n_0_2_1367), .ZN(n_0_2_1248));
   NAND2_X1 i_0_2_1287 (.A1(n_0_2_54), .A2(n_0_2_1251), .ZN(n_0_2_1249));
   OR2_X1 i_0_2_1288 (.A1(n_0_2_54), .A2(n_0_2_1251), .ZN(n_0_2_1250));
   AOI22_X1 i_0_2_1289 (.A1(n_0_2_1384), .A2(n_0_2_1252), .B1(n_0_2_1386), 
      .B2(n_0_2_1366), .ZN(n_0_2_1251));
   XNOR2_X1 i_0_2_1290 (.A(n_0_2_1381), .B(n_0_2_1253), .ZN(n_0_2_1252));
   NAND2_X1 i_0_2_1291 (.A1(in_b[0]), .A2(n_0_2_1254), .ZN(n_0_2_1253));
   AND2_X1 i_0_2_1292 (.A1(n_0_2_1257), .A2(n_0_2_1256), .ZN(n_0_2_1254));
   AOI21_X1 i_0_2_1293 (.A(n_0_2_1411), .B1(n_0_2_1410), .B2(n_0_2_1258), 
      .ZN(n_0_2_1256));
   OAI21_X1 i_0_2_1294 (.A(n_0_2_1285), .B1(n_0_2_1410), .B2(n_0_2_1258), 
      .ZN(n_0_2_1257));
   AOI22_X1 i_0_2_1295 (.A1(n_0_2_209), .A2(n_0_2_1263), .B1(n_0_2_1261), 
      .B2(n_0_2_1259), .ZN(n_0_2_1258));
   XNOR2_X1 i_0_2_1296 (.A(n_0_2_1290), .B(n_0_2_1260), .ZN(n_0_2_1259));
   NAND3_X1 i_0_2_1297 (.A1(n_0_2_1293), .A2(n_0_2_1292), .A3(n_0_2_1282), 
      .ZN(n_0_2_1260));
   OR2_X1 i_0_2_1298 (.A1(n_0_2_209), .A2(n_0_2_1263), .ZN(n_0_2_1261));
   NAND2_X1 i_0_2_1299 (.A1(n_0_2_209), .A2(n_0_2_1263), .ZN(n_0_2_1262));
   OAI21_X1 i_0_2_1300 (.A(n_0_2_1266), .B1(n_0_2_1267), .B2(n_0_2_1264), 
      .ZN(n_0_2_1263));
   XNOR2_X1 i_0_2_1301 (.A(n_0_2_1295), .B(n_0_2_1265), .ZN(n_0_2_1264));
   NAND3_X1 i_0_2_1302 (.A1(n_0_2_1298), .A2(n_0_2_1297), .A3(n_0_2_1282), 
      .ZN(n_0_2_1265));
   NAND2_X1 i_0_2_1303 (.A1(n_0_2_147), .A2(n_0_2_1268), .ZN(n_0_2_1266));
   NOR2_X1 i_0_2_1304 (.A1(n_0_2_147), .A2(n_0_2_1268), .ZN(n_0_2_1267));
   AOI22_X1 i_0_2_1305 (.A1(n_0_2_1403), .A2(n_0_2_1273), .B1(n_0_2_1272), 
      .B2(n_0_2_1269), .ZN(n_0_2_1268));
   XNOR2_X1 i_0_2_1306 (.A(n_0_2_1300), .B(n_0_2_1270), .ZN(n_0_2_1269));
   AOI211_X1 i_0_2_1307 (.A(n_0_2_1302), .B(n_0_2_1281), .C1(n_0_2_1400), 
      .C2(n_0_2_1304), .ZN(n_0_2_1270));
   NAND2_X1 i_0_2_1308 (.A1(n_0_2_1403), .A2(n_0_2_1273), .ZN(n_0_2_1271));
   OR2_X1 i_0_2_1309 (.A1(n_0_2_1403), .A2(n_0_2_1273), .ZN(n_0_2_1272));
   AOI22_X1 i_0_2_1310 (.A1(n_0_2_54), .A2(n_0_2_1278), .B1(n_0_2_1277), 
      .B2(n_0_2_1274), .ZN(n_0_2_1273));
   XNOR2_X1 i_0_2_1311 (.A(n_0_2_1307), .B(n_0_2_1275), .ZN(n_0_2_1274));
   NAND3_X1 i_0_2_1312 (.A1(n_0_2_1312), .A2(n_0_2_1306), .A3(n_0_2_1282), 
      .ZN(n_0_2_1275));
   NAND2_X1 i_0_2_1313 (.A1(n_0_2_54), .A2(n_0_2_1278), .ZN(n_0_2_1276));
   OR2_X1 i_0_2_1314 (.A1(n_0_2_54), .A2(n_0_2_1278), .ZN(n_0_2_1277));
   AOI22_X1 i_0_2_1315 (.A1(n_0_2_1284), .A2(n_0_2_1279), .B1(n_0_2_1381), 
      .B2(n_0_2_1366), .ZN(n_0_2_1278));
   XNOR2_X1 i_0_2_1316 (.A(n_0_2_1313), .B(n_0_2_1280), .ZN(n_0_2_1279));
   NOR2_X1 i_0_2_1317 (.A1(n_0_2_1405), .A2(n_0_2_1281), .ZN(n_0_2_1280));
   INV_X1 i_0_2_1318 (.A(n_0_2_1282), .ZN(n_0_2_1281));
   AOI21_X1 i_0_2_1319 (.A(n_0_2_1287), .B1(n_0_2_1314), .B2(n_0_2_1283), 
      .ZN(n_0_2_1282));
   NAND2_X1 i_0_2_1320 (.A1(n_0_2_209), .A2(n_0_2_1288), .ZN(n_0_2_1283));
   AOI21_X1 i_0_2_1321 (.A(n_0_2_1397), .B1(n_0_2_49), .B2(n_0_2_1380), .ZN(
      n_0_2_1284));
   AND2_X1 i_0_2_1322 (.A1(n_0_2_1370), .A2(n_0_2_1286), .ZN(n_0_2_1285));
   NAND2_X1 i_0_2_1323 (.A1(n_0_2_1315), .A2(n_0_2_1287), .ZN(n_0_2_1286));
   OAI21_X1 i_0_2_1324 (.A(n_0_2_1409), .B1(n_0_2_209), .B2(n_0_2_1288), 
      .ZN(n_0_2_1287));
   NAND2_X1 i_0_2_1325 (.A1(n_0_2_1292), .A2(n_0_2_1289), .ZN(n_0_2_1288));
   NAND2_X1 i_0_2_1326 (.A1(n_0_2_1293), .A2(n_0_2_1290), .ZN(n_0_2_1289));
   XNOR2_X1 i_0_2_1327 (.A(n_0_2_1318), .B(n_0_2_1291), .ZN(n_0_2_1290));
   NAND3_X1 i_0_2_1328 (.A1(n_0_2_1321), .A2(n_0_2_1320), .A3(n_0_2_1309), 
      .ZN(n_0_2_1291));
   NAND2_X1 i_0_2_1329 (.A1(n_0_2_147), .A2(n_0_2_1294), .ZN(n_0_2_1292));
   OR2_X1 i_0_2_1330 (.A1(n_0_2_147), .A2(n_0_2_1294), .ZN(n_0_2_1293));
   AOI22_X1 i_0_2_1331 (.A1(n_0_2_1403), .A2(n_0_2_1299), .B1(n_0_2_1297), 
      .B2(n_0_2_1295), .ZN(n_0_2_1294));
   XNOR2_X1 i_0_2_1332 (.A(n_0_2_1323), .B(n_0_2_1296), .ZN(n_0_2_1295));
   OAI211_X1 i_0_2_1333 (.A(n_0_2_1325), .B(n_0_2_1309), .C1(n_0_2_54), .C2(
      n_0_2_1327), .ZN(n_0_2_1296));
   OR2_X1 i_0_2_1334 (.A1(n_0_2_1403), .A2(n_0_2_1299), .ZN(n_0_2_1297));
   NAND2_X1 i_0_2_1335 (.A1(n_0_2_1403), .A2(n_0_2_1299), .ZN(n_0_2_1298));
   AOI21_X1 i_0_2_1336 (.A(n_0_2_1302), .B1(n_0_2_1303), .B2(n_0_2_1300), 
      .ZN(n_0_2_1299));
   XNOR2_X1 i_0_2_1337 (.A(n_0_2_1329), .B(n_0_2_1301), .ZN(n_0_2_1300));
   NOR3_X1 i_0_2_1338 (.A1(n_0_2_1349), .A2(n_0_2_1328), .A3(n_0_2_1310), 
      .ZN(n_0_2_1301));
   NOR2_X1 i_0_2_1339 (.A1(n_0_2_1400), .A2(n_0_2_1304), .ZN(n_0_2_1302));
   NAND2_X1 i_0_2_1340 (.A1(n_0_2_1400), .A2(n_0_2_1304), .ZN(n_0_2_1303));
   AOI21_X1 i_0_2_1341 (.A(n_0_2_1305), .B1(n_0_2_1312), .B2(n_0_2_1307), 
      .ZN(n_0_2_1304));
   INV_X1 i_0_2_1342 (.A(n_0_2_1306), .ZN(n_0_2_1305));
   AOI21_X1 i_0_2_1343 (.A(n_0_2_1397), .B1(n_0_2_49), .B2(n_0_2_1313), .ZN(
      n_0_2_1306));
   XNOR2_X1 i_0_2_1344 (.A(n_0_2_1351), .B(n_0_2_1308), .ZN(n_0_2_1307));
   NAND2_X1 i_0_2_1345 (.A1(in_b[0]), .A2(n_0_2_1309), .ZN(n_0_2_1308));
   INV_X1 i_0_2_1346 (.A(n_0_2_1310), .ZN(n_0_2_1309));
   NAND2_X1 i_0_2_1347 (.A1(n_0_2_1316), .A2(n_0_2_1311), .ZN(n_0_2_1310));
   OAI22_X1 i_0_2_1348 (.A1(n_0_2_1353), .A2(n_0_2_1333), .B1(n_0_2_1406), 
      .B2(n_0_2_1317), .ZN(n_0_2_1311));
   OR2_X1 i_0_2_1349 (.A1(n_0_2_1367), .A2(n_0_2_1313), .ZN(n_0_2_1312));
   XNOR2_X1 i_0_2_1350 (.A(in_a[10]), .B(n_0_2_1379), .ZN(n_0_2_1313));
   INV_X1 i_0_2_1351 (.A(n_0_2_1315), .ZN(n_0_2_1314));
   NOR2_X1 i_0_2_1352 (.A1(n_0_2_1353), .A2(n_0_2_1316), .ZN(n_0_2_1315));
   OAI21_X1 i_0_2_1353 (.A(n_0_2_1404), .B1(n_0_2_1407), .B2(n_0_2_1317), 
      .ZN(n_0_2_1316));
   AOI22_X1 i_0_2_1354 (.A1(n_0_2_96), .A2(n_0_2_1322), .B1(n_0_2_1321), 
      .B2(n_0_2_1318), .ZN(n_0_2_1317));
   XOR2_X1 i_0_2_1355 (.A(n_0_2_1337), .B(n_0_2_1319), .Z(n_0_2_1318));
   AND3_X1 i_0_2_1356 (.A1(n_0_2_1339), .A2(n_0_2_1336), .A3(n_0_2_1331), 
      .ZN(n_0_2_1319));
   NAND2_X1 i_0_2_1357 (.A1(n_0_2_96), .A2(n_0_2_1322), .ZN(n_0_2_1320));
   OR2_X1 i_0_2_1358 (.A1(n_0_2_96), .A2(n_0_2_1322), .ZN(n_0_2_1321));
   OAI21_X1 i_0_2_1359 (.A(n_0_2_1325), .B1(n_0_2_1326), .B2(n_0_2_1323), 
      .ZN(n_0_2_1322));
   XNOR2_X1 i_0_2_1360 (.A(n_0_2_1341), .B(n_0_2_1324), .ZN(n_0_2_1323));
   NAND3_X1 i_0_2_1361 (.A1(n_0_2_1346), .A2(n_0_2_1345), .A3(n_0_2_1331), 
      .ZN(n_0_2_1324));
   NAND2_X1 i_0_2_1362 (.A1(n_0_2_54), .A2(n_0_2_1327), .ZN(n_0_2_1325));
   NOR2_X1 i_0_2_1363 (.A1(n_0_2_54), .A2(n_0_2_1327), .ZN(n_0_2_1326));
   AOI21_X1 i_0_2_1364 (.A(n_0_2_1328), .B1(n_0_2_1350), .B2(n_0_2_1329), 
      .ZN(n_0_2_1327));
   NOR2_X1 i_0_2_1365 (.A1(n_0_2_1367), .A2(n_0_2_1351), .ZN(n_0_2_1328));
   XNOR2_X1 i_0_2_1366 (.A(n_0_2_1348), .B(n_0_2_1330), .ZN(n_0_2_1329));
   NAND2_X1 i_0_2_1367 (.A1(in_b[0]), .A2(n_0_2_1331), .ZN(n_0_2_1330));
   INV_X1 i_0_2_1368 (.A(n_0_2_1332), .ZN(n_0_2_1331));
   OAI21_X1 i_0_2_1369 (.A(n_0_2_1333), .B1(n_0_2_96), .B2(n_0_2_1335), .ZN(
      n_0_2_1332));
   AOI21_X1 i_0_2_1370 (.A(n_0_2_1404), .B1(n_0_2_1336), .B2(n_0_2_1334), 
      .ZN(n_0_2_1333));
   AOI22_X1 i_0_2_1371 (.A1(n_0_2_1339), .A2(n_0_2_1337), .B1(n_0_2_96), 
      .B2(n_0_2_1335), .ZN(n_0_2_1334));
   NAND2_X1 i_0_2_1372 (.A1(n_0_2_1370), .A2(n_0_2_1353), .ZN(n_0_2_1335));
   NAND2_X1 i_0_2_1373 (.A1(n_0_2_54), .A2(n_0_2_1340), .ZN(n_0_2_1336));
   XNOR2_X1 i_0_2_1374 (.A(n_0_2_1359), .B(n_0_2_1338), .ZN(n_0_2_1337));
   NAND3_X1 i_0_2_1375 (.A1(n_0_2_1357), .A2(n_0_2_1355), .A3(n_0_2_1343), 
      .ZN(n_0_2_1338));
   OR2_X1 i_0_2_1376 (.A1(n_0_2_54), .A2(n_0_2_1340), .ZN(n_0_2_1339));
   AOI22_X1 i_0_2_1377 (.A1(n_0_2_1366), .A2(n_0_2_1348), .B1(n_0_2_1346), 
      .B2(n_0_2_1341), .ZN(n_0_2_1340));
   XNOR2_X1 i_0_2_1378 (.A(n_0_2_1358), .B(n_0_2_1342), .ZN(n_0_2_1341));
   NAND2_X1 i_0_2_1379 (.A1(in_b[0]), .A2(n_0_2_1343), .ZN(n_0_2_1342));
   NOR3_X1 i_0_2_1380 (.A1(n_0_2_1401), .A2(n_0_2_1354), .A3(n_0_2_1344), 
      .ZN(n_0_2_1343));
   NOR2_X1 i_0_2_1381 (.A1(n_0_2_54), .A2(n_0_2_1363), .ZN(n_0_2_1344));
   NAND2_X1 i_0_2_1382 (.A1(n_0_2_1366), .A2(n_0_2_1348), .ZN(n_0_2_1345));
   INV_X1 i_0_2_1383 (.A(n_0_2_1347), .ZN(n_0_2_1346));
   AOI21_X1 i_0_2_1384 (.A(n_0_2_1398), .B1(in_b[0]), .B2(n_0_2_1348), .ZN(
      n_0_2_1347));
   XOR2_X1 i_0_2_1385 (.A(in_a[12]), .B(n_0_2_1377), .Z(n_0_2_1348));
   INV_X1 i_0_2_1386 (.A(n_0_2_1350), .ZN(n_0_2_1349));
   AOI21_X1 i_0_2_1387 (.A(n_0_2_1397), .B1(n_0_2_49), .B2(n_0_2_1351), .ZN(
      n_0_2_1350));
   XOR2_X1 i_0_2_1388 (.A(in_a[11]), .B(n_0_2_1378), .Z(n_0_2_1351));
   OAI21_X1 i_0_2_1389 (.A(n_0_2_1363), .B1(n_0_2_1401), .B2(n_0_2_1354), 
      .ZN(n_0_2_1353));
   AOI221_X1 i_0_2_1390 (.A(n_0_2_1356), .B1(n_0_2_54), .B2(n_0_2_1363), 
      .C1(n_0_2_1359), .C2(n_0_2_1357), .ZN(n_0_2_1354));
   INV_X1 i_0_2_1391 (.A(n_0_2_1356), .ZN(n_0_2_1355));
   OAI21_X1 i_0_2_1392 (.A(n_0_2_1412), .B1(n_0_2_1398), .B2(n_0_2_1358), 
      .ZN(n_0_2_1356));
   NAND2_X1 i_0_2_1393 (.A1(n_0_2_1366), .A2(n_0_2_1358), .ZN(n_0_2_1357));
   XOR2_X1 i_0_2_1394 (.A(in_a[13]), .B(n_0_2_1375), .Z(n_0_2_1358));
   AOI21_X1 i_0_2_1395 (.A(n_0_2_1365), .B1(in_b[0]), .B2(n_0_2_1360), .ZN(
      n_0_2_1359));
   INV_X1 i_0_2_1396 (.A(n_0_2_1361), .ZN(n_0_2_1360));
   OAI21_X1 i_0_2_1397 (.A(n_0_2_1364), .B1(n_0_2_1369), .B2(n_0_2_1362), 
      .ZN(n_0_2_1361));
   AOI21_X1 i_0_2_1398 (.A(n_0_2_1398), .B1(in_b[0]), .B2(n_0_2_1365), .ZN(
      n_0_2_1362));
   AOI21_X1 i_0_2_1399 (.A(n_0_2_1368), .B1(n_0_2_1398), .B2(n_0_2_1364), 
      .ZN(n_0_2_1363));
   AOI21_X1 i_0_2_1400 (.A(n_0_2_1399), .B1(n_0_2_1366), .B2(n_0_2_1365), 
      .ZN(n_0_2_1364));
   XNOR2_X1 i_0_2_1401 (.A(in_a[14]), .B(n_0_2_1374), .ZN(n_0_2_1365));
   INV_X1 i_0_2_1402 (.A(n_0_2_1367), .ZN(n_0_2_1366));
   NAND2_X1 i_0_2_1403 (.A1(in_b[0]), .A2(n_0_2_1398), .ZN(n_0_2_1367));
   INV_X1 i_0_2_1404 (.A(n_0_2_1369), .ZN(n_0_2_1368));
   AOI21_X1 i_0_2_1405 (.A(n_0_2_1372), .B1(in_b[0]), .B2(n_0_2_1396), .ZN(
      n_0_2_1369));
   NAND2_X1 i_0_2_1406 (.A1(n_0_2_1395), .A2(n_0_2_1371), .ZN(n_0_2_1370));
   INV_X1 i_0_2_1407 (.A(n_0_2_1372), .ZN(n_0_2_1371));
   XNOR2_X1 i_0_2_1408 (.A(n_0_2_1451), .B(n_0_2_1373), .ZN(n_0_2_1372));
   AOI21_X1 i_0_2_1409 (.A(n_0_2_1374), .B1(in_a[63]), .B2(in_a[14]), .ZN(
      n_0_2_1373));
   AOI21_X1 i_0_2_1410 (.A(n_0_2_1452), .B1(n_0_2_1450), .B2(n_0_2_1375), 
      .ZN(n_0_2_1374));
   OAI21_X1 i_0_2_1411 (.A(in_a[63]), .B1(in_a[12]), .B2(n_0_2_1376), .ZN(
      n_0_2_1375));
   INV_X1 i_0_2_1412 (.A(n_0_2_1377), .ZN(n_0_2_1376));
   OAI21_X1 i_0_2_1413 (.A(in_a[63]), .B1(in_a[11]), .B2(n_0_2_1378), .ZN(
      n_0_2_1377));
   AOI21_X1 i_0_2_1414 (.A(n_0_2_1452), .B1(n_0_2_1449), .B2(n_0_2_1379), 
      .ZN(n_0_2_1378));
   AOI21_X1 i_0_2_1415 (.A(n_0_2_1382), .B1(in_a[63]), .B2(in_a[9]), .ZN(
      n_0_2_1379));
   INV_X1 i_0_2_1416 (.A(n_0_2_1381), .ZN(n_0_2_1380));
   XNOR2_X1 i_0_2_1417 (.A(in_a[9]), .B(n_0_2_1382), .ZN(n_0_2_1381));
   NAND2_X1 i_0_2_1418 (.A1(n_0_2_1388), .A2(n_0_2_1383), .ZN(n_0_2_1382));
   OAI21_X1 i_0_2_1419 (.A(in_a[63]), .B1(in_a[8]), .B2(in_a[7]), .ZN(n_0_2_1383));
   AOI21_X1 i_0_2_1420 (.A(n_0_2_1397), .B1(n_0_2_49), .B2(n_0_2_1385), .ZN(
      n_0_2_1384));
   INV_X1 i_0_2_1421 (.A(n_0_2_1386), .ZN(n_0_2_1385));
   XNOR2_X1 i_0_2_1422 (.A(in_a[8]), .B(n_0_2_1387), .ZN(n_0_2_1386));
   AOI21_X1 i_0_2_1423 (.A(n_0_2_1452), .B1(n_0_2_1448), .B2(n_0_2_1388), 
      .ZN(n_0_2_1387));
   OAI21_X1 i_0_2_1424 (.A(in_a[63]), .B1(in_a[6]), .B2(n_0_2_1389), .ZN(
      n_0_2_1388));
   NAND2_X1 i_0_2_1425 (.A1(n_0_2_1447), .A2(n_0_2_1390), .ZN(n_0_2_1389));
   NOR2_X1 i_0_2_1426 (.A1(in_a[4]), .A2(n_0_2_1391), .ZN(n_0_2_1390));
   NAND3_X1 i_0_2_1427 (.A1(n_0_2_1445), .A2(n_0_2_1392), .A3(n_0_2_1446), 
      .ZN(n_0_2_1391));
   NOR2_X1 i_0_2_1428 (.A1(in_a[1]), .A2(n_0_2_1393), .ZN(n_0_2_1392));
   NOR2_X1 i_0_2_1429 (.A1(n_0_2_1452), .A2(n_0_2_1444), .ZN(n_0_2_1393));
   INV_X1 i_0_2_1430 (.A(n_0_2_1395), .ZN(n_0_2_1394));
   NOR2_X1 i_0_2_1431 (.A1(n_0_2_1399), .A2(n_0_2_1412), .ZN(n_0_2_1395));
   NOR2_X1 i_0_2_1432 (.A1(n_0_2_1399), .A2(n_0_2_1398), .ZN(n_0_2_1396));
   INV_X1 i_0_2_1433 (.A(n_0_2_1412), .ZN(n_0_2_1397));
   NAND2_X1 i_0_2_1434 (.A1(n_0_2_1405), .A2(n_0_2_49), .ZN(n_0_2_1412));
   INV_X1 i_0_2_1435 (.A(n_0_2_49), .ZN(n_0_2_1398));
   AOI22_X1 i_0_2_1436 (.A1(in_b[63]), .A2(n_0_1), .B1(n_0_2_1454), .B2(in_b[1]), 
      .ZN(n_0_2_49));
   NAND2_X1 i_0_2_1437 (.A1(n_0_2_1402), .A2(n_0_2_54), .ZN(n_0_2_1399));
   INV_X1 i_0_2_1438 (.A(n_0_2_54), .ZN(n_0_2_1400));
   OAI22_X1 i_0_2_1439 (.A1(in_b[63]), .A2(in_b[2]), .B1(n_0_2_1454), .B2(n_0_2), 
      .ZN(n_0_2_54));
   INV_X1 i_0_2_1440 (.A(n_0_2_1402), .ZN(n_0_2_1401));
   NOR2_X1 i_0_2_1441 (.A1(n_0_2_1404), .A2(n_0_2_1403), .ZN(n_0_2_1402));
   INV_X1 i_0_2_1442 (.A(n_0_2_96), .ZN(n_0_2_1403));
   AOI22_X1 i_0_2_1443 (.A1(in_b[63]), .A2(n_0_3), .B1(n_0_2_1454), .B2(in_b[3]), 
      .ZN(n_0_2_96));
   OR2_X1 i_0_2_1444 (.A1(n_0_2_1407), .A2(n_0_2_1406), .ZN(n_0_2_1404));
   INV_X1 i_0_2_1445 (.A(n_0_2_147), .ZN(n_0_2_1406));
   AOI22_X1 i_0_2_1446 (.A1(in_b[63]), .A2(n_0_4), .B1(n_0_2_1454), .B2(in_b[4]), 
      .ZN(n_0_2_147));
   NAND2_X1 i_0_2_1447 (.A1(n_0_2_1409), .A2(n_0_2_209), .ZN(n_0_2_1407));
   INV_X1 i_0_2_1448 (.A(n_0_2_209), .ZN(n_0_2_1408));
   AOI22_X1 i_0_2_1449 (.A1(in_b[63]), .A2(n_0_5), .B1(n_0_2_1454), .B2(in_b[5]), 
      .ZN(n_0_2_209));
   NOR2_X1 i_0_2_1450 (.A1(n_0_2_1411), .A2(n_0_2_1410), .ZN(n_0_2_1409));
   INV_X1 i_0_2_1451 (.A(n_0_2_281), .ZN(n_0_2_1410));
   AOI22_X1 i_0_2_1452 (.A1(in_b[63]), .A2(n_0_6), .B1(n_0_2_1454), .B2(in_b[6]), 
      .ZN(n_0_2_281));
   NAND2_X1 i_0_2_1453 (.A1(n_0_2_1414), .A2(n_0_2_363), .ZN(n_0_2_1411));
   INV_X1 i_0_2_1454 (.A(n_0_2_363), .ZN(n_0_2_1413));
   AOI22_X1 i_0_2_1455 (.A1(in_b[63]), .A2(n_0_7), .B1(n_0_2_1454), .B2(in_b[7]), 
      .ZN(n_0_2_363));
   NOR2_X1 i_0_2_1456 (.A1(n_0_2_1416), .A2(n_0_2_1415), .ZN(n_0_2_1414));
   INV_X1 i_0_2_1457 (.A(n_0_2_453), .ZN(n_0_2_1415));
   AOI22_X1 i_0_2_1458 (.A1(in_b[63]), .A2(n_0_8), .B1(n_0_2_1454), .B2(in_b[8]), 
      .ZN(n_0_2_453));
   OR3_X1 i_0_2_1459 (.A1(n_0_2_1419), .A2(n_0_2_1418), .A3(n_0_2_1417), 
      .ZN(n_0_2_1416));
   INV_X1 i_0_2_1460 (.A(n_0_2_458), .ZN(n_0_2_1417));
   OAI22_X1 i_0_2_1461 (.A1(in_b[63]), .A2(in_b[9]), .B1(n_0_2_1454), .B2(n_0_9), 
      .ZN(n_0_2_458));
   INV_X1 i_0_2_1462 (.A(n_0_2_660), .ZN(n_0_2_1418));
   OAI22_X1 i_0_2_1463 (.A1(in_b[63]), .A2(in_b[10]), .B1(n_0_2_1454), .B2(
      n_0_10), .ZN(n_0_2_660));
   OR2_X1 i_0_2_1464 (.A1(n_0_2_1440), .A2(n_0_2_1420), .ZN(n_0_2_1419));
   NAND2_X1 i_0_2_1465 (.A1(n_0_2_1423), .A2(n_0_2_907), .ZN(n_0_2_1420));
   INV_X1 i_0_2_1466 (.A(n_0_2_907), .ZN(n_0_2_1421));
   OAI22_X1 i_0_2_1467 (.A1(in_b[63]), .A2(in_b[12]), .B1(n_0_2_1454), .B2(
      n_0_12), .ZN(n_0_2_907));
   INV_X1 i_0_2_1468 (.A(n_0_2_1423), .ZN(n_0_2_1422));
   NOR2_X1 i_0_2_1469 (.A1(n_0_2_1425), .A2(n_0_2_1424), .ZN(n_0_2_1423));
   INV_X1 i_0_2_1470 (.A(n_0_2_1044), .ZN(n_0_2_1424));
   OAI22_X1 i_0_2_1471 (.A1(in_b[63]), .A2(in_b[13]), .B1(n_0_2_1454), .B2(
      n_0_13), .ZN(n_0_2_1044));
   NAND3_X1 i_0_2_1472 (.A1(n_0_2_1190), .A2(n_0_2_1426), .A3(n_0_2_1430), 
      .ZN(n_0_2_1425));
   NOR2_X1 i_0_2_1473 (.A1(n_0_2_1428), .A2(n_0_2_1427), .ZN(n_0_2_1426));
   INV_X1 i_0_2_1474 (.A(n_0_2_1352), .ZN(n_0_2_1427));
   OAI22_X1 i_0_2_1475 (.A1(in_b[63]), .A2(in_b[15]), .B1(n_0_2_1454), .B2(
      n_0_15), .ZN(n_0_2_1352));
   INV_X1 i_0_2_1476 (.A(n_0_2_1516), .ZN(n_0_2_1428));
   OAI22_X1 i_0_2_1477 (.A1(in_b[63]), .A2(in_b[16]), .B1(n_0_2_1454), .B2(
      n_0_16), .ZN(n_0_2_1516));
   INV_X1 i_0_2_1478 (.A(n_0_2_1190), .ZN(n_0_2_1429));
   OAI22_X1 i_0_2_1479 (.A1(in_b[63]), .A2(in_b[14]), .B1(n_0_2_1454), .B2(
      n_0_14), .ZN(n_0_2_1190));
   AND2_X1 i_0_2_1480 (.A1(n_0_2_154), .A2(n_0_2_1431), .ZN(n_0_2_1430));
   NOR2_X1 i_0_2_1481 (.A1(n_0_2_1433), .A2(n_0_2_1432), .ZN(n_0_2_1431));
   INV_X1 i_0_2_1482 (.A(n_0_2_667), .ZN(n_0_2_1432));
   OAI22_X1 i_0_2_1483 (.A1(in_b[63]), .A2(in_b[22]), .B1(n_0_2_1454), .B2(
      n_0_22), .ZN(n_0_2_667));
   INV_X1 i_0_2_1484 (.A(n_0_2_50), .ZN(n_0_2_1433));
   OAI22_X1 i_0_2_1485 (.A1(in_b[63]), .A2(in_b[21]), .B1(n_0_2_1454), .B2(
      n_0_21), .ZN(n_0_2_50));
   INV_X1 i_0_2_1486 (.A(n_0_2_51), .ZN(n_0_2_154));
   NAND2_X1 i_0_2_1487 (.A1(n_0_2_1197), .A2(n_0_2_52), .ZN(n_0_2_51));
   INV_X1 i_0_2_1488 (.A(n_0_2_52), .ZN(n_0_2_1434));
   OAI22_X1 i_0_2_1489 (.A1(in_b[63]), .A2(in_b[17]), .B1(n_0_2_1454), .B2(
      n_0_17), .ZN(n_0_2_52));
   INV_X1 i_0_2_1490 (.A(n_0_2_1435), .ZN(n_0_2_1197));
   NAND2_X1 i_0_2_1491 (.A1(n_0_2_1437), .A2(n_0_2_53), .ZN(n_0_2_1435));
   INV_X1 i_0_2_1492 (.A(n_0_2_53), .ZN(n_0_2_1436));
   OAI22_X1 i_0_2_1493 (.A1(in_b[63]), .A2(in_b[18]), .B1(n_0_2_1454), .B2(
      n_0_18), .ZN(n_0_2_53));
   NOR2_X1 i_0_2_1494 (.A1(n_0_2_1439), .A2(n_0_2_1438), .ZN(n_0_2_1437));
   INV_X1 i_0_2_1495 (.A(n_0_2_55), .ZN(n_0_2_1438));
   OAI22_X1 i_0_2_1496 (.A1(in_b[63]), .A2(in_b[19]), .B1(n_0_2_1454), .B2(
      n_0_19), .ZN(n_0_2_55));
   INV_X1 i_0_2_1497 (.A(n_0_2_56), .ZN(n_0_2_1439));
   OAI22_X1 i_0_2_1498 (.A1(in_b[63]), .A2(in_b[20]), .B1(n_0_2_1454), .B2(
      n_0_20), .ZN(n_0_2_56));
   INV_X1 i_0_2_1499 (.A(n_0_2_780), .ZN(n_0_2_1440));
   OAI22_X1 i_0_2_1500 (.A1(in_b[63]), .A2(in_b[11]), .B1(n_0_2_1454), .B2(
      n_0_11), .ZN(n_0_2_780));
   OR2_X1 i_0_2_1501 (.A1(ovfl_flag), .A2(divide_by_zero_error), .ZN(err));
   INV_X1 i_0_2_1502 (.A(n_0_28), .ZN(n_0_2_1441));
   INV_X1 i_0_2_1503 (.A(n_0_29), .ZN(n_0_2_1442));
   INV_X1 i_0_2_1504 (.A(n_0_30), .ZN(n_0_2_1443));
   INV_X1 i_0_2_1505 (.A(in_a[0]), .ZN(n_0_2_1444));
   INV_X1 i_0_2_1506 (.A(in_a[2]), .ZN(n_0_2_1445));
   INV_X1 i_0_2_1507 (.A(in_a[3]), .ZN(n_0_2_1446));
   INV_X1 i_0_2_1508 (.A(in_a[5]), .ZN(n_0_2_1447));
   INV_X1 i_0_2_1509 (.A(in_a[7]), .ZN(n_0_2_1448));
   INV_X1 i_0_2_1510 (.A(in_a[10]), .ZN(n_0_2_1449));
   INV_X1 i_0_2_1511 (.A(in_a[13]), .ZN(n_0_2_1450));
   INV_X1 i_0_2_1512 (.A(in_a[15]), .ZN(n_0_2_1451));
   INV_X1 i_0_2_1513 (.A(in_a[63]), .ZN(n_0_2_1452));
   INV_X1 i_0_2_1514 (.A(in_b[0]), .ZN(n_0_2_1405));
   INV_X1 i_0_2_1515 (.A(in_b[8]), .ZN(n_0_2_1453));
   INV_X1 i_0_2_1516 (.A(in_b[63]), .ZN(n_0_2_1454));
   AND2_X1 i_0_2_1517 (.A1(n_0_2_30), .A2(n_0_2_316), .ZN(n_0_2_1455));
   OAI22_X1 i_0_2_1518 (.A1(n_0_2_1455), .A2(n_0_2_281), .B1(n_0_2_30), .B2(
      n_0_2_316), .ZN(n_0_2_1456));
   AOI21_X1 i_0_2_1519 (.A(n_0_2_315), .B1(n_0_2_1456), .B2(n_0_2_340), .ZN(
      n_0_2_1457));
   OR2_X1 i_0_2_1520 (.A1(n_0_2_32), .A2(n_0_2_453), .ZN(n_0_2_1458));
   AOI22_X1 i_0_2_1521 (.A1(n_0_2_1457), .A2(n_0_2_1458), .B1(n_0_2_32), 
      .B2(n_0_2_453), .ZN(n_0_2_1459));
   AOI21_X1 i_0_2_1522 (.A(n_0_2_314), .B1(n_0_2_1459), .B2(n_0_2_345), .ZN(
      n_0_2_1460));
   AND2_X1 i_0_2_1523 (.A1(n_0_2_34), .A2(n_0_2_660), .ZN(n_0_2_1461));
   OAI22_X1 i_0_2_1524 (.A1(n_0_2_1460), .A2(n_0_2_1461), .B1(n_0_2_34), 
      .B2(n_0_2_660), .ZN(n_0_2_1462));
   AOI21_X1 i_0_2_1525 (.A(n_0_2_313), .B1(n_0_2_1462), .B2(n_0_2_350), .ZN(
      n_0_2_1463));
   OR2_X1 i_0_2_1526 (.A1(n_0_2_36), .A2(n_0_2_907), .ZN(n_0_2_1464));
   AOI22_X1 i_0_2_1527 (.A1(n_0_2_1463), .A2(n_0_2_1464), .B1(n_0_2_36), 
      .B2(n_0_2_907), .ZN(n_0_2_1465));
   AOI21_X1 i_0_2_1528 (.A(n_0_2_312), .B1(n_0_2_1465), .B2(n_0_2_355), .ZN(
      n_0_2_1466));
   OR2_X1 i_0_2_1529 (.A1(n_0_2_1190), .A2(n_0_2_38), .ZN(n_0_2_1467));
   AOI22_X1 i_0_2_1530 (.A1(n_0_2_1466), .A2(n_0_2_1467), .B1(n_0_2_1190), 
      .B2(n_0_2_38), .ZN(n_0_2_1468));
   AOI21_X1 i_0_2_1531 (.A(n_0_2_311), .B1(n_0_2_1468), .B2(n_0_2_360), .ZN(
      n_0_2_1469));
   OR2_X1 i_0_2_1532 (.A1(n_0_2_1516), .A2(n_0_2_40), .ZN(n_0_2_1470));
   AOI22_X1 i_0_2_1533 (.A1(n_0_2_1469), .A2(n_0_2_1470), .B1(n_0_2_1516), 
      .B2(n_0_2_40), .ZN(n_0_2_1471));
   AOI21_X1 i_0_2_1534 (.A(n_0_2_310), .B1(n_0_2_1471), .B2(n_0_2_366), .ZN(
      n_0_2_1472));
   AND2_X1 i_0_2_1535 (.A1(n_0_2_53), .A2(n_0_2_42), .ZN(n_0_2_1473));
   OAI22_X1 i_0_2_1536 (.A1(n_0_2_1472), .A2(n_0_2_1473), .B1(n_0_2_53), 
      .B2(n_0_2_42), .ZN(n_0_2_1474));
   AOI21_X1 i_0_2_1537 (.A(n_0_2_309), .B1(n_0_2_1474), .B2(n_0_2_371), .ZN(
      n_0_2_1475));
   INV_X1 i_0_2_1538 (.A(n_0_2_56), .ZN(n_0_2_1476));
   INV_X1 i_0_2_1539 (.A(n_0_2_44), .ZN(n_0_2_1477));
   NAND2_X1 i_0_2_1540 (.A1(n_0_2_1476), .A2(n_0_2_1477), .ZN(n_0_2_1478));
   AOI22_X1 i_0_2_1541 (.A1(n_0_2_1475), .A2(n_0_2_1478), .B1(n_0_2_56), 
      .B2(n_0_2_44), .ZN(n_0_2_1479));
   AOI211_X1 i_0_2_1542 (.A(n_0_2_305), .B(n_0_2_1432), .C1(n_0_2_1479), 
      .C2(n_0_2_306), .ZN(n_0_2_1480));
   INV_X1 i_0_2_1543 (.A(n_0_2_1480), .ZN(n_0_2_1481));
   NOR2_X1 i_0_2_1544 (.A1(n_0_2_1481), .A2(n_0_2_1395), .ZN(quotient[1]));
   INV_X1 i_0_2_1545 (.A(n_0_2_847), .ZN(n_0_2_1482));
   OAI22_X1 i_0_2_1546 (.A1(quotient[1]), .A2(n_0_2_847), .B1(n_0_23), .B2(
      n_0_2_1482), .ZN(n_0_2_1483));
   INV_X1 i_0_2_1547 (.A(n_0_2_1483), .ZN(n_0_42));
   XOR2_X1 i_0_2_1548 (.A(n_0_2_1479), .B(n_0_2_278), .Z(n_0_2_1484));
   INV_X1 i_0_2_1549 (.A(n_0_2_24), .ZN(n_0_2_1485));
   OAI22_X1 i_0_2_1550 (.A1(n_0_2_1481), .A2(n_0_2_1484), .B1(n_0_2_1480), 
      .B2(n_0_2_1485), .ZN(n_0_2_1486));
   OAI21_X1 i_0_2_1551 (.A(n_0_2_1394), .B1(n_0_2_1486), .B2(n_0_2_667), 
      .ZN(n_0_2_1487));
   XNOR2_X1 i_0_2_1552 (.A(n_0_2_1466), .B(n_0_2_286), .ZN(n_0_2_1488));
   AOI22_X1 i_0_2_1553 (.A1(n_0_2_1481), .A2(n_0_2_38), .B1(n_0_2_1480), 
      .B2(n_0_2_1488), .ZN(n_0_2_1489));
   INV_X1 i_0_2_1554 (.A(n_0_2_1352), .ZN(n_0_2_1490));
   XNOR2_X1 i_0_2_1555 (.A(n_0_2_1465), .B(n_0_2_288), .ZN(n_0_2_1491));
   AOI22_X1 i_0_2_1556 (.A1(n_0_2_1481), .A2(n_0_2_37), .B1(n_0_2_1480), 
      .B2(n_0_2_1491), .ZN(n_0_2_1492));
   INV_X1 i_0_2_1557 (.A(n_0_2_1190), .ZN(n_0_2_1493));
   AOI22_X1 i_0_2_1558 (.A1(n_0_2_1489), .A2(n_0_2_1490), .B1(n_0_2_1492), 
      .B2(n_0_2_1493), .ZN(n_0_2_1494));
   AOI22_X1 i_0_2_1559 (.A1(n_0_2_1481), .A2(n_0_2_28), .B1(n_0_2_1480), 
      .B2(n_0_2_298), .ZN(n_0_2_1495));
   INV_X1 i_0_2_1560 (.A(n_0_2_209), .ZN(n_0_2_1496));
   AOI22_X1 i_0_2_1561 (.A1(n_0_2_1481), .A2(n_0_2_29), .B1(n_0_2_1480), 
      .B2(n_0_2_296), .ZN(n_0_2_1497));
   INV_X1 i_0_2_1562 (.A(n_0_2_281), .ZN(n_0_2_1498));
   AOI22_X1 i_0_2_1563 (.A1(n_0_2_1495), .A2(n_0_2_1496), .B1(n_0_2_1497), 
      .B2(n_0_2_1498), .ZN(n_0_2_1499));
   OAI21_X1 i_0_2_1564 (.A(in_b[0]), .B1(n_0_2_49), .B2(n_0_2_1405), .ZN(
      n_0_2_1500));
   OAI21_X1 i_0_2_1565 (.A(n_0_2_1412), .B1(n_0_2_1481), .B2(n_0_2_1500), 
      .ZN(n_0_2_1501));
   NOR2_X1 i_0_2_1566 (.A1(n_0_2_1501), .A2(n_0_2_54), .ZN(n_0_2_1502));
   AOI222_X1 i_0_2_1567 (.A1(n_0_2_1501), .A2(n_0_2_54), .B1(n_0_2_1481), 
      .B2(n_0_2_25), .C1(n_0_2_1480), .C2(n_0_2_304), .ZN(n_0_2_1503));
   AOI22_X1 i_0_2_1568 (.A1(n_0_2_1481), .A2(n_0_2_26), .B1(n_0_2_1480), 
      .B2(n_0_2_302), .ZN(n_0_2_1504));
   INV_X1 i_0_2_1569 (.A(n_0_2_96), .ZN(n_0_2_1505));
   AOI211_X1 i_0_2_1570 (.A(n_0_2_1502), .B(n_0_2_1503), .C1(n_0_2_1504), 
      .C2(n_0_2_1505), .ZN(n_0_2_1506));
   INV_X1 i_0_2_1571 (.A(n_0_2_1504), .ZN(n_0_2_1507));
   AOI21_X1 i_0_2_1572 (.A(n_0_2_1506), .B1(n_0_2_1507), .B2(n_0_2_96), .ZN(
      n_0_2_1508));
   INV_X1 i_0_2_1573 (.A(n_0_2_147), .ZN(n_0_2_1509));
   AOI22_X1 i_0_2_1574 (.A1(n_0_2_1481), .A2(n_0_2_27), .B1(n_0_2_1480), 
      .B2(n_0_2_300), .ZN(n_0_2_1510));
   AOI21_X1 i_0_2_1575 (.A(n_0_2_1508), .B1(n_0_2_1509), .B2(n_0_2_1510), 
      .ZN(n_0_2_1511));
   OAI22_X1 i_0_2_1576 (.A1(n_0_2_1495), .A2(n_0_2_1496), .B1(n_0_2_1510), 
      .B2(n_0_2_1509), .ZN(n_0_2_1512));
   OAI21_X1 i_0_2_1577 (.A(n_0_2_1499), .B1(n_0_2_1511), .B2(n_0_2_1512), 
      .ZN(n_0_2_1513));
   INV_X1 i_0_2_1578 (.A(n_0_2_295), .ZN(n_0_2_1514));
   INV_X1 i_0_2_1579 (.A(n_0_2_316), .ZN(n_0_2_1515));
   OAI221_X1 i_0_2_1580 (.A(n_0_2_1480), .B1(n_0_2_295), .B2(n_0_2_316), 
      .C1(n_0_2_1514), .C2(n_0_2_1515), .ZN(n_0_2_1517));
   OAI21_X1 i_0_2_1581 (.A(n_0_2_1517), .B1(n_0_2_30), .B2(n_0_2_1480), .ZN(
      n_0_2_1518));
   INV_X1 i_0_2_1582 (.A(n_0_2_363), .ZN(n_0_2_1519));
   OAI221_X1 i_0_2_1583 (.A(n_0_2_1513), .B1(n_0_2_1518), .B2(n_0_2_1519), 
      .C1(n_0_2_1498), .C2(n_0_2_1497), .ZN(n_0_2_1520));
   INV_X1 i_0_2_1584 (.A(n_0_2_1518), .ZN(n_0_2_1521));
   XOR2_X1 i_0_2_1585 (.A(n_0_2_1456), .B(n_0_2_294), .Z(n_0_2_1523));
   INV_X1 i_0_2_1586 (.A(n_0_2_31), .ZN(n_0_2_1524));
   OAI22_X1 i_0_2_1587 (.A1(n_0_2_1481), .A2(n_0_2_1523), .B1(n_0_2_1480), 
      .B2(n_0_2_1524), .ZN(n_0_2_1526));
   OAI221_X1 i_0_2_1588 (.A(n_0_2_1520), .B1(n_0_2_363), .B2(n_0_2_1521), 
      .C1(n_0_2_453), .C2(n_0_2_1526), .ZN(n_0_2_1527));
   XNOR2_X1 i_0_2_1589 (.A(n_0_2_1457), .B(n_0_2_293), .ZN(n_0_2_1529));
   AOI22_X1 i_0_2_1590 (.A1(n_0_2_1481), .A2(n_0_2_32), .B1(n_0_2_1480), 
      .B2(n_0_2_1529), .ZN(n_0_2_1530));
   INV_X1 i_0_2_1591 (.A(n_0_2_1530), .ZN(n_0_2_1532));
   AOI22_X1 i_0_2_1592 (.A1(n_0_2_1532), .A2(n_0_2_458), .B1(n_0_2_1526), 
      .B2(n_0_2_453), .ZN(n_0_2_1533));
   INV_X1 i_0_2_1593 (.A(n_0_2_660), .ZN(n_0_2_1535));
   XNOR2_X1 i_0_2_1594 (.A(n_0_2_1459), .B(n_0_2_292), .ZN(n_0_2_1536));
   AOI22_X1 i_0_2_1595 (.A1(n_0_2_1481), .A2(n_0_2_33), .B1(n_0_2_1480), 
      .B2(n_0_2_1536), .ZN(n_0_2_1538));
   INV_X1 i_0_2_1596 (.A(n_0_2_458), .ZN(n_0_2_1539));
   AOI222_X1 i_0_2_1597 (.A1(n_0_2_1527), .A2(n_0_2_1533), .B1(n_0_2_1535), 
      .B2(n_0_2_1538), .C1(n_0_2_1539), .C2(n_0_2_1530), .ZN(n_0_2_1541));
   XNOR2_X1 i_0_2_1598 (.A(n_0_2_1460), .B(n_0_2_291), .ZN(n_0_2_1542));
   AOI22_X1 i_0_2_1599 (.A1(n_0_2_1481), .A2(n_0_2_34), .B1(n_0_2_1480), 
      .B2(n_0_2_1542), .ZN(n_0_2_1544));
   INV_X1 i_0_2_1600 (.A(n_0_2_780), .ZN(n_0_2_1545));
   OAI22_X1 i_0_2_1601 (.A1(n_0_2_1544), .A2(n_0_2_1545), .B1(n_0_2_1538), 
      .B2(n_0_2_1535), .ZN(n_0_2_1547));
   XOR2_X1 i_0_2_1602 (.A(n_0_2_1462), .B(n_0_2_290), .Z(n_0_2_1548));
   INV_X1 i_0_2_1603 (.A(n_0_2_35), .ZN(n_0_2_1550));
   OAI22_X1 i_0_2_1604 (.A1(n_0_2_1481), .A2(n_0_2_1548), .B1(n_0_2_1480), 
      .B2(n_0_2_1550), .ZN(n_0_2_1551));
   INV_X1 i_0_2_1605 (.A(n_0_2_1544), .ZN(n_0_2_1553));
   OAI222_X1 i_0_2_1606 (.A1(n_0_2_1541), .A2(n_0_2_1547), .B1(n_0_2_907), 
      .B2(n_0_2_1551), .C1(n_0_2_780), .C2(n_0_2_1553), .ZN(n_0_2_1554));
   NAND2_X1 i_0_2_1607 (.A1(n_0_2_1551), .A2(n_0_2_907), .ZN(n_0_2_1556));
   XNOR2_X1 i_0_2_1608 (.A(n_0_2_1463), .B(n_0_2_289), .ZN(n_0_2_1557));
   AOI22_X1 i_0_2_1609 (.A1(n_0_2_1481), .A2(n_0_2_36), .B1(n_0_2_1480), 
      .B2(n_0_2_1557), .ZN(n_0_2_1559));
   INV_X1 i_0_2_1610 (.A(n_0_2_1044), .ZN(n_0_2_1560));
   AOI22_X1 i_0_2_1611 (.A1(n_0_2_1554), .A2(n_0_2_1556), .B1(n_0_2_1559), 
      .B2(n_0_2_1560), .ZN(n_0_2_1562));
   OAI22_X1 i_0_2_1612 (.A1(n_0_2_1492), .A2(n_0_2_1493), .B1(n_0_2_1559), 
      .B2(n_0_2_1560), .ZN(n_0_2_1563));
   OAI21_X1 i_0_2_1613 (.A(n_0_2_1494), .B1(n_0_2_1562), .B2(n_0_2_1563), 
      .ZN(n_0_2_1565));
   INV_X1 i_0_2_1614 (.A(n_0_2_1516), .ZN(n_0_2_1566));
   XNOR2_X1 i_0_2_1615 (.A(n_0_2_1468), .B(n_0_2_285), .ZN(n_0_2_1568));
   AOI22_X1 i_0_2_1616 (.A1(n_0_2_1481), .A2(n_0_2_39), .B1(n_0_2_1480), 
      .B2(n_0_2_1568), .ZN(n_0_2_1569));
   OAI221_X1 i_0_2_1617 (.A(n_0_2_1565), .B1(n_0_2_1566), .B2(n_0_2_1569), 
      .C1(n_0_2_1490), .C2(n_0_2_1489), .ZN(n_0_2_1571));
   XNOR2_X1 i_0_2_1618 (.A(n_0_2_1469), .B(n_0_2_284), .ZN(n_0_2_1572));
   AOI22_X1 i_0_2_1619 (.A1(n_0_2_1481), .A2(n_0_2_40), .B1(n_0_2_1480), 
      .B2(n_0_2_1572), .ZN(n_0_2_1574));
   INV_X1 i_0_2_1620 (.A(n_0_2_52), .ZN(n_0_2_1575));
   AOI22_X1 i_0_2_1621 (.A1(n_0_2_1574), .A2(n_0_2_1575), .B1(n_0_2_1569), 
      .B2(n_0_2_1566), .ZN(n_0_2_1576));
   INV_X1 i_0_2_1622 (.A(n_0_2_1574), .ZN(n_0_2_1577));
   XOR2_X1 i_0_2_1623 (.A(n_0_2_1471), .B(n_0_2_283), .Z(n_0_2_1578));
   INV_X1 i_0_2_1624 (.A(n_0_2_41), .ZN(n_0_2_1580));
   OAI22_X1 i_0_2_1625 (.A1(n_0_2_1481), .A2(n_0_2_1578), .B1(n_0_2_1480), 
      .B2(n_0_2_1580), .ZN(n_0_2_1581));
   AOI222_X1 i_0_2_1626 (.A1(n_0_2_1571), .A2(n_0_2_1576), .B1(n_0_2_52), 
      .B2(n_0_2_1577), .C1(n_0_2_53), .C2(n_0_2_1581), .ZN(n_0_2_1582));
   XNOR2_X1 i_0_2_1627 (.A(n_0_2_1472), .B(n_0_2_282), .ZN(n_0_2_1583));
   AOI22_X1 i_0_2_1628 (.A1(n_0_2_1481), .A2(n_0_2_42), .B1(n_0_2_1480), 
      .B2(n_0_2_1583), .ZN(n_0_2_1584));
   INV_X1 i_0_2_1629 (.A(n_0_2_1584), .ZN(n_0_2_1586));
   OAI22_X1 i_0_2_1630 (.A1(n_0_2_1581), .A2(n_0_2_53), .B1(n_0_2_1586), 
      .B2(n_0_2_55), .ZN(n_0_2_1587));
   XNOR2_X1 i_0_2_1631 (.A(n_0_2_1474), .B(n_0_2_280), .ZN(n_0_2_1592));
   AOI22_X1 i_0_2_1632 (.A1(n_0_2_1481), .A2(n_0_2_43), .B1(n_0_2_1480), 
      .B2(n_0_2_1592), .ZN(n_0_2_1593));
   INV_X1 i_0_2_1633 (.A(n_0_2_55), .ZN(n_0_2_1594));
   OAI222_X1 i_0_2_1634 (.A1(n_0_2_1582), .A2(n_0_2_1587), .B1(n_0_2_1476), 
      .B2(n_0_2_1593), .C1(n_0_2_1594), .C2(n_0_2_1584), .ZN(n_0_2_1596));
   INV_X1 i_0_2_1635 (.A(n_0_2_1593), .ZN(n_0_2_1597));
   XOR2_X1 i_0_2_1636 (.A(n_0_2_1475), .B(n_0_2_279), .Z(n_0_2_1599));
   OAI22_X1 i_0_2_1637 (.A1(n_0_2_1481), .A2(n_0_2_1599), .B1(n_0_2_1480), 
      .B2(n_0_2_1477), .ZN(n_0_2_1600));
   OAI221_X1 i_0_2_1638 (.A(n_0_2_1596), .B1(n_0_2_1597), .B2(n_0_2_56), 
      .C1(n_0_2_50), .C2(n_0_2_1600), .ZN(n_0_2_1601));
   AOI22_X1 i_0_2_1639 (.A1(n_0_2_1486), .A2(n_0_2_667), .B1(n_0_2_1600), 
      .B2(n_0_2_50), .ZN(n_0_2_1603));
   AOI21_X1 i_0_2_1640 (.A(n_0_2_1487), .B1(n_0_2_1601), .B2(n_0_2_1603), 
      .ZN(quotient[0]));
endmodule
