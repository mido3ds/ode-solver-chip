/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sat Apr 25 19:54:56 2020
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 492112353 */

module datapath__1_13515(to_int6128, p_0);
   input [7:0]to_int6128;
   output p_0;

   NOR3_X1 i_0 (.A1(to_int6128[5]), .A2(n_0), .A3(to_int6128[6]), .ZN(p_0));
   OR4_X1 i_1 (.A1(to_int6128[2]), .A2(to_int6128[1]), .A3(to_int6128[3]), 
      .A4(to_int6128[4]), .ZN(n_0));
endmodule

module datapath__1_13522(to_int6128, p_0);
   input [7:0]to_int6128;
   output p_0;

   NOR3_X1 i_0 (.A1(to_int6128[5]), .A2(n_0), .A3(to_int6128[6]), .ZN(p_0));
   OR3_X1 i_1 (.A1(to_int6128[3]), .A2(to_int6128[2]), .A3(to_int6128[4]), 
      .ZN(n_0));
endmodule

module half_adder__3_459(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   INV_X1 i_2 (.A(a), .ZN(f));
endmodule

module half_adder__3_456(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;

   INV_X1 i_0_0 (.A(n_0_0), .ZN(f));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(n_0_4), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(n_0_3), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(a), .ZN(n_0_2));
   INV_X1 i_0_4 (.A(b), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(n_0_4), .ZN(cout));
   NAND2_X1 i_0_6 (.A1(a), .A2(b), .ZN(n_0_4));
endmodule

module half_adder__3_453(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(a), .A2(b), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_3), .A2(n_1_4), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module half_adder__3_450(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_0_0;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   INV_X1 i_0_0 (.A(n_0_0), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(n_0_0));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(a), .A2(b), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_3), .A2(n_1_4), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module half_adder__3_447(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_0_0;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   INV_X1 i_0_0 (.A(n_0_0), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(n_0_0));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(a), .A2(b), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_3), .A2(n_1_4), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module half_adder__3_444(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   AND2_X1 i_0_0 (.A1(b), .A2(a), .ZN(cout));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(b), .A2(a), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_4), .A2(n_1_3), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module half_adder__3_441(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(a), .A2(b), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_3), .A2(n_1_4), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module incrementor__3_460(a, enbl, c);
   input [6:0]a;
   input enbl;
   output [6:0]c;

   half_adder__3_459 half_adder_0_0_half_adder_0_i (.a(a[0]), .b(), .cout(), 
      .f(c[0]));
   half_adder__3_456 half_adder_0_1_half_adder_0_i (.a(a[1]), .b(a[0]), .cout(
      n_0), .f(c[1]));
   half_adder__3_453 half_adder_0_2_half_adder_0_i (.a(a[2]), .b(n_0), .cout(n_1), 
      .f(c[2]));
   half_adder__3_450 half_adder_0_3_half_adder_0_i (.a(a[3]), .b(n_1), .cout(n_2), 
      .f(c[3]));
   half_adder__3_447 half_adder_0_4_half_adder_0_i (.a(a[4]), .b(n_2), .cout(n_3), 
      .f(c[4]));
   half_adder__3_444 half_adder_0_5_half_adder_0_i (.a(a[5]), .b(n_3), .cout(n_4), 
      .f(c[5]));
   half_adder__3_441 half_adder_0_6_half_adder_0_i (.a(a[6]), .b(n_4), .cout(), 
      .f(c[6]));
endmodule

module full_adder__3_437(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(f));
   AND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(cout));
endmodule

module full_adder__3_433(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_6), .ZN(cout));
   NOR2_X1 i_0_1 (.A1(n_0_1), .A2(n_0_0), .ZN(f));
   AOI21_X1 i_0_2 (.A(cin), .B1(n_0_3), .B2(n_0_6), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_2), .ZN(n_0_1));
   NAND3_X1 i_0_4 (.A1(n_0_3), .A2(cin), .A3(n_0_6), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(n_0_4), .A2(n_0_5), .ZN(n_0_3));
   INV_X1 i_0_6 (.A(a), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(b), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(a), .A2(b), .ZN(n_0_6));
endmodule

module full_adder__3_429(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;

   NAND2_X1 i_0_11 (.A1(cin), .A2(b), .ZN(n_0_9));
   NAND2_X1 i_0_12 (.A1(n_0_11), .A2(n_0_0), .ZN(n_0_10));
   INV_X1 i_0_13 (.A(cin), .ZN(n_0_11));
   INV_X1 i_0_14 (.A(b), .ZN(n_0_0));
   OAI21_X1 i_0_0 (.A(n_0_1), .B1(n_0_2), .B2(n_0_3), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(n_0_1));
   NOR2_X1 i_0_2 (.A1(a), .A2(b), .ZN(n_0_2));
   INV_X1 i_0_3 (.A(cin), .ZN(n_0_3));
   INV_X1 i_0_4 (.A(n_0_4), .ZN(f));
   NAND2_X1 i_0_5 (.A1(n_0_6), .A2(n_0_5), .ZN(n_0_4));
   NAND3_X1 i_0_6 (.A1(a), .A2(n_0_9), .A3(n_0_10), .ZN(n_0_5));
   NAND2_X1 i_0_7 (.A1(n_0_8), .A2(n_0_7), .ZN(n_0_6));
   OAI21_X1 i_0_8 (.A(n_0_9), .B1(b), .B2(cin), .ZN(n_0_7));
   INV_X1 i_0_9 (.A(a), .ZN(n_0_8));
endmodule

module full_adder__3_425(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;

   INV_X1 i_0_0 (.A(n_0_1), .ZN(cout));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(f));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(n_0_1), .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(a), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_4), .A2(n_0_3), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(cin), .ZN(n_0_3));
   INV_X1 i_0_6 (.A(a), .ZN(n_0_4));
endmodule

module full_adder__3_421(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;

   INV_X1 i_0_0 (.A(n_0_1), .ZN(cout));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(f));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(n_0_1), .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(a), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_4), .A2(n_0_3), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(cin), .ZN(n_0_3));
   INV_X1 i_0_6 (.A(a), .ZN(n_0_4));
endmodule

module full_adder__3_417(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;

   INV_X1 i_0_0 (.A(n_0_1), .ZN(cout));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(f));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(n_0_1), .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(a), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_4), .A2(n_0_3), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(cin), .ZN(n_0_3));
   INV_X1 i_0_6 (.A(a), .ZN(n_0_4));
endmodule

module full_adder__3_413(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;

   INV_X1 i_0_0 (.A(n_0_0), .ZN(f));
   NAND2_X1 i_0_1 (.A1(n_0_2), .A2(n_0_1), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(a), .A2(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(n_0_3), .A2(n_0_4), .ZN(n_0_2));
   INV_X1 i_0_4 (.A(a), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(cin), .ZN(n_0_4));
endmodule

module int_adder__3_438(a, b, cin, enbl, c, cout);
   input [6:0]a;
   input [2:0]b;
   input cin;
   input enbl;
   output [6:0]c;
   output cout;

   full_adder__3_437 full_adder_0_0_full_adder_0_i (.a(a[0]), .b(b[0]), .cin(), 
      .f(c[0]), .cout(n_0));
   full_adder__3_433 full_adder_0_1_full_adder_0_i (.a(a[1]), .b(b[1]), .cin(n_0), 
      .f(c[1]), .cout(n_1));
   full_adder__3_429 full_adder_0_2_full_adder_0_i (.a(a[2]), .b(b[2]), .cin(n_1), 
      .f(c[2]), .cout(n_2));
   full_adder__3_425 full_adder_0_3_full_adder_0_i (.a(a[3]), .b(), .cin(n_2), 
      .f(c[3]), .cout(n_3));
   full_adder__3_421 full_adder_0_4_full_adder_0_i (.a(a[4]), .b(), .cin(n_3), 
      .f(c[4]), .cout(n_4));
   full_adder__3_417 full_adder_0_5_full_adder_0_i (.a(a[5]), .b(), .cin(n_4), 
      .f(c[5]), .cout(n_5));
   full_adder__3_413 full_adder_0_6_full_adder_0_i (.a(a[6]), .b(), .cin(n_5), 
      .f(c[6]), .cout());
endmodule

module range_extractor__3_461(in_a, in_size, out_a, out_b);
   input [6:0]in_a;
   input [2:0]in_size;
   output [6:0]out_a;
   output [6:0]out_b;

   incrementor__3_460 inc (.a(in_a), .enbl(), .c(out_a));
   int_adder__3_438 add (.a(out_a), .b(in_size), .cin(), .enbl(), .c(out_b), 
      .cout());
endmodule

module datapath__1_13511(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   NAND2_X1 i_0 (.A1(n_1), .A2(n_0), .ZN(p_0));
   NOR4_X1 i_1 (.A1(to_int5359[2]), .A2(to_int5359[0]), .A3(to_int5359[6]), 
      .A4(to_int5359[3]), .ZN(n_0));
   NOR3_X1 i_2 (.A1(to_int5359[5]), .A2(to_int5359[4]), .A3(to_int5359[1]), 
      .ZN(n_1));
endmodule

module datapath__1_7666(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NAND2_X1 i_0 (.A1(n_1), .A2(n_0), .ZN(p_0));
   NOR3_X1 i_1 (.A1(to_int6126[6]), .A2(to_int6126[5]), .A3(to_int6126[4]), 
      .ZN(n_0));
   NOR4_X1 i_2 (.A1(to_int6126[2]), .A2(to_int6126[0]), .A3(to_int6126[3]), 
      .A4(to_int6126[1]), .ZN(n_1));
endmodule

module datapath__1_7740(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NAND2_X1 i_0 (.A1(n_4), .A2(n_0), .ZN(p_0));
   NOR4_X1 i_1 (.A1(to_int6126[5]), .A2(to_int6126[4]), .A3(to_int6126[3]), 
      .A4(n_1), .ZN(n_0));
   NAND2_X1 i_2 (.A1(n_2), .A2(n_3), .ZN(n_1));
   NAND2_X1 i_3 (.A1(to_int6126[1]), .A2(to_int6126[0]), .ZN(n_2));
   INV_X1 i_4 (.A(to_int6126[2]), .ZN(n_3));
   INV_X1 i_5 (.A(to_int6126[6]), .ZN(n_4));
endmodule

module datapath__1_18134(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NOR2_X1 i_0 (.A1(n_1), .A2(n_0), .ZN(p_0));
   NAND3_X1 i_1 (.A1(to_int6126[6]), .A2(to_int6126[3]), .A3(to_int6126[1]), 
      .ZN(n_0));
   NAND4_X1 i_2 (.A1(to_int6126[2]), .A2(to_int6126[0]), .A3(to_int6126[5]), 
      .A4(to_int6126[4]), .ZN(n_1));
endmodule

module datapath__1_14001(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0));
   NAND2_X1 i_1 (.A1(to_int6126[6]), .A2(n_1), .ZN(n_0));
   INV_X1 i_2 (.A(n_2), .ZN(n_1));
   NAND4_X1 i_3 (.A1(to_int6126[5]), .A2(to_int6126[4]), .A3(to_int6126[3]), 
      .A4(n_3), .ZN(n_2));
   NAND2_X1 i_4 (.A1(n_5), .A2(n_4), .ZN(n_3));
   NAND2_X1 i_5 (.A1(to_int6126[1]), .A2(to_int6126[0]), .ZN(n_4));
   INV_X1 i_6 (.A(to_int6126[2]), .ZN(n_5));
endmodule

module datapath__1_13985(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   AND4_X1 i_0 (.A1(to_int6126[5]), .A2(n_0), .A3(to_int6126[6]), .A4(
      to_int6126[4]), .ZN(p_0));
   OR2_X1 i_1 (.A1(to_int6126[3]), .A2(n_1), .ZN(n_0));
   AND3_X1 i_2 (.A1(to_int6126[2]), .A2(to_int6126[1]), .A3(to_int6126[0]), 
      .ZN(n_1));
endmodule

module datapath__1_13961(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   AND4_X1 i_0 (.A1(to_int6126[5]), .A2(n_0), .A3(to_int6126[6]), .A4(
      to_int6126[4]), .ZN(p_0));
   OR4_X1 i_1 (.A1(to_int6126[2]), .A2(to_int6126[0]), .A3(to_int6126[3]), 
      .A4(to_int6126[1]), .ZN(n_0));
endmodule

module datapath__1_13953(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0));
   OAI211_X1 i_1 (.A(to_int6126[5]), .B(to_int6126[6]), .C1(to_int6126[4]), 
      .C2(n_1), .ZN(n_0));
   AND4_X1 i_2 (.A1(to_int6126[3]), .A2(to_int6126[2]), .A3(to_int6126[1]), 
      .A4(to_int6126[0]), .ZN(n_1));
endmodule

module datapath__1_13945(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   AOI21_X1 i_0 (.A(n_0), .B1(n_2), .B2(n_1), .ZN(p_0));
   NAND2_X1 i_1 (.A1(to_int6126[6]), .A2(to_int6126[5]), .ZN(n_0));
   OAI211_X1 i_2 (.A(to_int6126[3]), .B(to_int6126[2]), .C1(to_int6126[1]), 
      .C2(to_int6126[0]), .ZN(n_1));
   INV_X1 i_3 (.A(to_int6126[4]), .ZN(n_2));
endmodule

module datapath__1_13937(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0));
   OAI211_X1 i_1 (.A(to_int6126[5]), .B(to_int6126[6]), .C1(to_int6126[4]), 
      .C2(n_1), .ZN(n_0));
   NOR2_X1 i_2 (.A1(n_3), .A2(n_2), .ZN(n_1));
   AOI21_X1 i_3 (.A(to_int6126[2]), .B1(to_int6126[1]), .B2(to_int6126[0]), 
      .ZN(n_2));
   INV_X1 i_4 (.A(to_int6126[3]), .ZN(n_3));
endmodule

module datapath__1_13929(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   OR3_X1 i_0 (.A1(to_int6126[1]), .A2(to_int6126[0]), .A3(to_int6126[2]), 
      .ZN(n_0));
   AOI21_X1 i_1 (.A(to_int6126[4]), .B1(n_0), .B2(to_int6126[3]), .ZN(n_1));
   INV_X1 i_2 (.A(n_1), .ZN(n_2));
   AND3_X1 i_3 (.A1(n_2), .A2(to_int6126[5]), .A3(to_int6126[6]), .ZN(p_0));
endmodule

module datapath__1_13913(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NOR2_X1 i_0 (.A1(n_1), .A2(n_0), .ZN(p_0));
   NAND2_X1 i_1 (.A1(to_int6126[6]), .A2(to_int6126[5]), .ZN(n_0));
   AOI211_X1 i_2 (.A(to_int6126[4]), .B(to_int6126[3]), .C1(to_int6126[2]), 
      .C2(n_2), .ZN(n_1));
   OR2_X1 i_3 (.A1(to_int6126[1]), .A2(to_int6126[0]), .ZN(n_2));
endmodule

module datapath__1_13905(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   AND3_X1 i_0 (.A1(to_int6126[5]), .A2(n_0), .A3(to_int6126[6]), .ZN(p_0));
   OR4_X1 i_1 (.A1(to_int6126[2]), .A2(n_1), .A3(to_int6126[3]), .A4(
      to_int6126[4]), .ZN(n_0));
   AND2_X1 i_2 (.A1(to_int6126[1]), .A2(to_int6126[0]), .ZN(n_1));
endmodule

module datapath__1_13897(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   AOI21_X1 i_0 (.A(n_0), .B1(n_2), .B2(n_1), .ZN(p_0));
   NAND2_X1 i_1 (.A1(to_int6126[6]), .A2(to_int6126[5]), .ZN(n_0));
   NOR4_X1 i_2 (.A1(to_int6126[2]), .A2(to_int6126[0]), .A3(to_int6126[3]), 
      .A4(to_int6126[1]), .ZN(n_1));
   INV_X1 i_3 (.A(to_int6126[4]), .ZN(n_2));
endmodule

module datapath__1_13889(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   AND4_X1 i_0 (.A1(to_int6126[3]), .A2(to_int6126[2]), .A3(to_int6126[1]), 
      .A4(to_int6126[0]), .ZN(n_0));
   AOI21_X1 i_1 (.A(to_int6126[5]), .B1(n_0), .B2(to_int6126[4]), .ZN(n_1));
   INV_X1 i_2 (.A(to_int6126[6]), .ZN(n_2));
   NOR2_X1 i_3 (.A1(n_1), .A2(n_2), .ZN(p_0));
endmodule

module datapath__1_13881(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0));
   OAI21_X1 i_1 (.A(to_int6126[6]), .B1(to_int6126[5]), .B2(n_1), .ZN(n_0));
   AND4_X1 i_2 (.A1(to_int6126[3]), .A2(to_int6126[2]), .A3(n_2), .A4(
      to_int6126[4]), .ZN(n_1));
   OR2_X1 i_3 (.A1(to_int6126[1]), .A2(to_int6126[0]), .ZN(n_2));
endmodule

module datapath__1_13873(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NAND2_X1 i_3 (.A1(to_int6126[4]), .A2(to_int6126[3]), .ZN(n_2));
   AOI21_X1 i_4 (.A(to_int6126[2]), .B1(to_int6126[1]), .B2(to_int6126[0]), 
      .ZN(n_3));
   INV_X1 i_0 (.A(n_0), .ZN(p_0));
   NAND2_X1 i_1 (.A1(to_int6126[6]), .A2(n_1), .ZN(n_0));
   OAI21_X1 i_2 (.A(n_4), .B1(n_2), .B2(n_3), .ZN(n_1));
   INV_X1 i_5 (.A(to_int6126[5]), .ZN(n_4));
endmodule

module datapath__1_13865(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0));
   OAI21_X1 i_1 (.A(to_int6126[6]), .B1(to_int6126[5]), .B2(n_1), .ZN(n_0));
   AND3_X1 i_2 (.A1(to_int6126[3]), .A2(n_2), .A3(to_int6126[4]), .ZN(n_1));
   OR3_X1 i_3 (.A1(to_int6126[1]), .A2(to_int6126[0]), .A3(to_int6126[2]), 
      .ZN(n_2));
endmodule

module datapath__1_13857(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0));
   OAI21_X1 i_1 (.A(to_int6126[6]), .B1(to_int6126[5]), .B2(n_1), .ZN(n_0));
   INV_X1 i_2 (.A(n_2), .ZN(n_1));
   OAI21_X1 i_3 (.A(to_int6126[4]), .B1(to_int6126[3]), .B2(n_3), .ZN(n_2));
   AND3_X1 i_4 (.A1(to_int6126[2]), .A2(to_int6126[1]), .A3(to_int6126[0]), 
      .ZN(n_3));
endmodule

module datapath__1_13849(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0));
   OAI21_X1 i_1 (.A(to_int6126[6]), .B1(to_int6126[5]), .B2(n_1), .ZN(n_0));
   INV_X1 i_2 (.A(n_2), .ZN(n_1));
   OAI221_X1 i_3 (.A(to_int6126[4]), .B1(to_int6126[3]), .B2(n_3), .C1(
      to_int6126[3]), .C2(to_int6126[2]), .ZN(n_2));
   OR2_X1 i_4 (.A1(to_int6126[1]), .A2(to_int6126[0]), .ZN(n_3));
endmodule

module datapath__1_13841(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0));
   OAI21_X1 i_1 (.A(to_int6126[6]), .B1(to_int6126[5]), .B2(n_1), .ZN(n_0));
   INV_X1 i_2 (.A(n_2), .ZN(n_1));
   OAI21_X1 i_3 (.A(to_int6126[4]), .B1(to_int6126[3]), .B2(n_3), .ZN(n_2));
   INV_X1 i_4 (.A(n_4), .ZN(n_3));
   AOI21_X1 i_5 (.A(to_int6126[2]), .B1(to_int6126[1]), .B2(to_int6126[0]), 
      .ZN(n_4));
endmodule

module datapath__1_13833(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0));
   OAI21_X1 i_1 (.A(to_int6126[6]), .B1(to_int6126[5]), .B2(n_1), .ZN(n_0));
   INV_X1 i_2 (.A(n_2), .ZN(n_1));
   OAI21_X1 i_3 (.A(to_int6126[4]), .B1(to_int6126[1]), .B2(n_3), .ZN(n_2));
   OR3_X1 i_4 (.A1(to_int6126[2]), .A2(to_int6126[0]), .A3(to_int6126[3]), 
      .ZN(n_3));
endmodule

module datapath__1_13825(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   AND4_X1 i_0 (.A1(to_int6126[3]), .A2(to_int6126[2]), .A3(to_int6126[1]), 
      .A4(to_int6126[0]), .ZN(n_0));
   OR3_X1 i_1 (.A1(n_0), .A2(to_int6126[5]), .A3(to_int6126[4]), .ZN(n_1));
   AND2_X1 i_2 (.A1(n_1), .A2(to_int6126[6]), .ZN(p_0));
endmodule

module datapath__1_13817(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   AOI21_X1 i_0 (.A(n_2), .B1(n_1), .B2(n_0), .ZN(p_0));
   NOR2_X1 i_1 (.A1(to_int6126[5]), .A2(to_int6126[4]), .ZN(n_0));
   OAI211_X1 i_2 (.A(to_int6126[3]), .B(to_int6126[2]), .C1(to_int6126[1]), 
      .C2(to_int6126[0]), .ZN(n_1));
   INV_X1 i_3 (.A(to_int6126[6]), .ZN(n_2));
endmodule

module datapath__1_13809(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NOR2_X1 i_0 (.A1(n_3), .A2(n_0), .ZN(p_0));
   AOI211_X1 i_1 (.A(to_int6126[4]), .B(to_int6126[5]), .C1(to_int6126[3]), 
      .C2(n_1), .ZN(n_0));
   INV_X1 i_2 (.A(n_2), .ZN(n_1));
   AOI21_X1 i_3 (.A(to_int6126[2]), .B1(to_int6126[1]), .B2(to_int6126[0]), 
      .ZN(n_2));
   INV_X1 i_4 (.A(to_int6126[6]), .ZN(n_3));
endmodule

module datapath__1_13801(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NOR2_X1 i_0 (.A1(n_2), .A2(n_0), .ZN(p_0));
   AOI211_X1 i_1 (.A(to_int6126[4]), .B(to_int6126[5]), .C1(to_int6126[3]), 
      .C2(n_1), .ZN(n_0));
   OR3_X1 i_2 (.A1(to_int6126[1]), .A2(to_int6126[0]), .A3(to_int6126[2]), 
      .ZN(n_1));
   INV_X1 i_3 (.A(to_int6126[6]), .ZN(n_2));
endmodule

module datapath__1_13793(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   INV_X1 i_0 (.A(to_int6126[6]), .ZN(n_0));
   NAND3_X1 i_1 (.A1(to_int6126[2]), .A2(to_int6126[0]), .A3(to_int6126[1]), 
      .ZN(n_1));
   NOR3_X1 i_2 (.A1(to_int6126[4]), .A2(to_int6126[3]), .A3(to_int6126[5]), 
      .ZN(n_2));
   AOI21_X1 i_3 (.A(n_0), .B1(n_1), .B2(n_2), .ZN(p_0));
endmodule

module datapath__1_13785(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   AOI21_X1 i_0 (.A(n_2), .B1(n_1), .B2(n_0), .ZN(p_0));
   NOR3_X1 i_1 (.A1(to_int6126[4]), .A2(to_int6126[3]), .A3(to_int6126[5]), 
      .ZN(n_0));
   OAI21_X1 i_2 (.A(to_int6126[2]), .B1(to_int6126[1]), .B2(to_int6126[0]), 
      .ZN(n_1));
   INV_X1 i_3 (.A(to_int6126[6]), .ZN(n_2));
endmodule

module datapath__1_13777(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   INV_X1 i_0 (.A(to_int6126[6]), .ZN(n_0));
   NOR4_X1 i_1 (.A1(to_int6126[4]), .A2(to_int6126[3]), .A3(to_int6126[5]), 
      .A4(to_int6126[2]), .ZN(n_1));
   NAND2_X1 i_2 (.A1(to_int6126[1]), .A2(to_int6126[0]), .ZN(n_2));
   AOI21_X1 i_3 (.A(n_0), .B1(n_1), .B2(n_2), .ZN(p_0));
endmodule

module datapath__1_13769(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   INV_X1 i_0 (.A(to_int6126[6]), .ZN(n_0));
   NOR4_X1 i_1 (.A1(to_int6126[2]), .A2(to_int6126[0]), .A3(to_int6126[3]), 
      .A4(to_int6126[1]), .ZN(n_1));
   NOR2_X1 i_2 (.A1(to_int6126[5]), .A2(to_int6126[4]), .ZN(n_2));
   AOI21_X1 i_3 (.A(n_0), .B1(n_1), .B2(n_2), .ZN(p_0));
endmodule

module datapath__1_13762(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   OAI21_X1 i_0 (.A(n_2), .B1(n_1), .B2(n_0), .ZN(p_0));
   NAND2_X1 i_1 (.A1(to_int6126[5]), .A2(to_int6126[4]), .ZN(n_0));
   NAND4_X1 i_2 (.A1(to_int6126[3]), .A2(to_int6126[2]), .A3(to_int6126[1]), 
      .A4(to_int6126[0]), .ZN(n_1));
   INV_X1 i_3 (.A(to_int6126[6]), .ZN(n_2));
endmodule

module datapath__1_13754(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   OAI21_X1 i_0 (.A(n_2), .B1(n_1), .B2(n_0), .ZN(p_0));
   NAND4_X1 i_1 (.A1(to_int6126[4]), .A2(to_int6126[3]), .A3(to_int6126[5]), 
      .A4(to_int6126[2]), .ZN(n_0));
   NOR2_X1 i_2 (.A1(to_int6126[1]), .A2(to_int6126[0]), .ZN(n_1));
   INV_X1 i_3 (.A(to_int6126[6]), .ZN(n_2));
endmodule

module datapath__1_13746(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   OAI21_X1 i_0 (.A(n_2), .B1(n_1), .B2(n_0), .ZN(p_0));
   NAND3_X1 i_1 (.A1(to_int6126[4]), .A2(to_int6126[3]), .A3(to_int6126[5]), 
      .ZN(n_0));
   AOI21_X1 i_2 (.A(to_int6126[2]), .B1(to_int6126[1]), .B2(to_int6126[0]), 
      .ZN(n_1));
   INV_X1 i_3 (.A(to_int6126[6]), .ZN(n_2));
endmodule

module datapath__1_13738(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   OAI21_X1 i_0 (.A(n_2), .B1(n_1), .B2(n_0), .ZN(p_0));
   NAND3_X1 i_1 (.A1(to_int6126[4]), .A2(to_int6126[3]), .A3(to_int6126[5]), 
      .ZN(n_0));
   NOR3_X1 i_2 (.A1(to_int6126[1]), .A2(to_int6126[0]), .A3(to_int6126[2]), 
      .ZN(n_1));
   INV_X1 i_3 (.A(to_int6126[6]), .ZN(n_2));
endmodule

module datapath__1_13730(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NAND2_X1 i_0 (.A1(n_2), .A2(n_0), .ZN(p_0));
   OAI211_X1 i_1 (.A(to_int6126[4]), .B(to_int6126[5]), .C1(to_int6126[3]), 
      .C2(n_1), .ZN(n_0));
   AND3_X1 i_2 (.A1(to_int6126[1]), .A2(to_int6126[0]), .A3(to_int6126[2]), 
      .ZN(n_1));
   INV_X1 i_3 (.A(to_int6126[6]), .ZN(n_2));
endmodule

module datapath__1_13722(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NAND2_X1 i_0 (.A1(n_3), .A2(n_0), .ZN(p_0));
   OAI211_X1 i_1 (.A(to_int6126[4]), .B(to_int6126[5]), .C1(to_int6126[3]), 
      .C2(n_1), .ZN(n_0));
   INV_X1 i_2 (.A(n_2), .ZN(n_1));
   OAI21_X1 i_3 (.A(to_int6126[2]), .B1(to_int6126[1]), .B2(to_int6126[0]), 
      .ZN(n_2));
   INV_X1 i_4 (.A(to_int6126[6]), .ZN(n_3));
endmodule

module datapath__1_13714(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   OAI21_X1 i_0 (.A(n_2), .B1(n_1), .B2(n_0), .ZN(p_0));
   NAND2_X1 i_1 (.A1(to_int6126[5]), .A2(to_int6126[4]), .ZN(n_0));
   AOI211_X1 i_2 (.A(to_int6126[2]), .B(to_int6126[3]), .C1(to_int6126[1]), 
      .C2(to_int6126[0]), .ZN(n_1));
   INV_X1 i_3 (.A(to_int6126[6]), .ZN(n_2));
endmodule

module datapath__1_13706(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   OR2_X1 i_0 (.A1(to_int6126[6]), .A2(n_0), .ZN(p_0));
   AND3_X1 i_1 (.A1(to_int6126[4]), .A2(n_1), .A3(to_int6126[5]), .ZN(n_0));
   OR4_X1 i_2 (.A1(to_int6126[2]), .A2(to_int6126[0]), .A3(to_int6126[3]), 
      .A4(to_int6126[1]), .ZN(n_1));
endmodule

module datapath__1_13698(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   OAI21_X1 i_0 (.A(n_3), .B1(n_2), .B2(n_0), .ZN(p_0));
   AOI21_X1 i_1 (.A(to_int6126[4]), .B1(to_int6126[3]), .B2(n_1), .ZN(n_0));
   AND3_X1 i_2 (.A1(to_int6126[1]), .A2(to_int6126[0]), .A3(to_int6126[2]), 
      .ZN(n_1));
   INV_X1 i_3 (.A(to_int6126[5]), .ZN(n_2));
   INV_X1 i_4 (.A(to_int6126[6]), .ZN(n_3));
endmodule

module datapath__1_13690(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NAND2_X1 i_0 (.A1(n_3), .A2(n_0), .ZN(p_0));
   OAI21_X1 i_1 (.A(to_int6126[5]), .B1(to_int6126[4]), .B2(n_1), .ZN(n_0));
   INV_X1 i_2 (.A(n_2), .ZN(n_1));
   OAI211_X1 i_3 (.A(to_int6126[3]), .B(to_int6126[2]), .C1(to_int6126[1]), 
      .C2(to_int6126[0]), .ZN(n_2));
   INV_X1 i_4 (.A(to_int6126[6]), .ZN(n_3));
endmodule

module datapath__1_13682(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   OAI21_X1 i_0 (.A(n_4), .B1(n_3), .B2(n_0), .ZN(p_0));
   AOI21_X1 i_1 (.A(to_int6126[4]), .B1(to_int6126[3]), .B2(n_1), .ZN(n_0));
   INV_X1 i_2 (.A(n_2), .ZN(n_1));
   AOI21_X1 i_3 (.A(to_int6126[2]), .B1(to_int6126[1]), .B2(to_int6126[0]), 
      .ZN(n_2));
   INV_X1 i_4 (.A(to_int6126[5]), .ZN(n_3));
   INV_X1 i_5 (.A(to_int6126[6]), .ZN(n_4));
endmodule

module datapath__1_13674(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   OAI21_X1 i_0 (.A(n_3), .B1(n_2), .B2(n_0), .ZN(p_0));
   AOI21_X1 i_1 (.A(to_int6126[4]), .B1(to_int6126[3]), .B2(n_1), .ZN(n_0));
   OR3_X1 i_2 (.A1(to_int6126[1]), .A2(to_int6126[0]), .A3(to_int6126[2]), 
      .ZN(n_1));
   INV_X1 i_3 (.A(to_int6126[5]), .ZN(n_2));
   INV_X1 i_4 (.A(to_int6126[6]), .ZN(n_3));
endmodule

module datapath__1_13666(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NAND2_X1 i_0 (.A1(n_4), .A2(n_0), .ZN(p_0));
   OAI21_X1 i_1 (.A(to_int6126[5]), .B1(to_int6126[4]), .B2(n_1), .ZN(n_0));
   NAND2_X1 i_2 (.A1(n_3), .A2(n_2), .ZN(n_1));
   NAND3_X1 i_3 (.A1(to_int6126[2]), .A2(to_int6126[1]), .A3(to_int6126[0]), 
      .ZN(n_2));
   INV_X1 i_4 (.A(to_int6126[3]), .ZN(n_3));
   INV_X1 i_5 (.A(to_int6126[6]), .ZN(n_4));
endmodule

module datapath__1_13658(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   OAI21_X1 i_0 (.A(n_3), .B1(n_2), .B2(n_0), .ZN(p_0));
   AOI211_X1 i_1 (.A(to_int6126[4]), .B(to_int6126[3]), .C1(to_int6126[2]), 
      .C2(n_1), .ZN(n_0));
   OR2_X1 i_2 (.A1(to_int6126[1]), .A2(to_int6126[0]), .ZN(n_1));
   INV_X1 i_3 (.A(to_int6126[5]), .ZN(n_2));
   INV_X1 i_4 (.A(to_int6126[6]), .ZN(n_3));
endmodule

module datapath__1_13650(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   AND2_X1 i_0 (.A1(to_int6126[1]), .A2(to_int6126[0]), .ZN(n_0));
   NAND2_X1 i_1 (.A1(n_3), .A2(n_1), .ZN(p_0));
   OAI21_X1 i_2 (.A(to_int6126[5]), .B1(to_int6126[4]), .B2(n_2), .ZN(n_1));
   OR3_X1 i_3 (.A1(to_int6126[3]), .A2(to_int6126[2]), .A3(n_0), .ZN(n_2));
   INV_X1 i_4 (.A(to_int6126[6]), .ZN(n_3));
endmodule

module datapath__1_13642(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   OR2_X1 i_0 (.A1(to_int6126[2]), .A2(to_int6126[0]), .ZN(n_0));
   NAND2_X1 i_1 (.A1(n_3), .A2(n_1), .ZN(p_0));
   OAI21_X1 i_2 (.A(to_int6126[5]), .B1(to_int6126[4]), .B2(n_2), .ZN(n_1));
   OR3_X1 i_3 (.A1(to_int6126[3]), .A2(to_int6126[1]), .A3(n_0), .ZN(n_2));
   INV_X1 i_4 (.A(to_int6126[6]), .ZN(n_3));
endmodule

module datapath__1_13634(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   OAI21_X1 i_0 (.A(n_0), .B1(n_2), .B2(n_1), .ZN(p_0));
   NOR2_X1 i_1 (.A1(to_int6126[6]), .A2(to_int6126[5]), .ZN(n_0));
   NAND3_X1 i_2 (.A1(to_int6126[2]), .A2(to_int6126[1]), .A3(to_int6126[0]), 
      .ZN(n_1));
   NAND2_X1 i_3 (.A1(to_int6126[4]), .A2(to_int6126[3]), .ZN(n_2));
endmodule

module datapath__1_13626(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   OAI21_X1 i_0 (.A(n_0), .B1(n_2), .B2(n_1), .ZN(p_0));
   NOR2_X1 i_1 (.A1(to_int6126[6]), .A2(to_int6126[5]), .ZN(n_0));
   NAND3_X1 i_2 (.A1(to_int6126[4]), .A2(to_int6126[2]), .A3(to_int6126[3]), 
      .ZN(n_1));
   NOR2_X1 i_3 (.A1(to_int6126[1]), .A2(to_int6126[0]), .ZN(n_2));
endmodule

module datapath__1_13618(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   OAI21_X1 i_0 (.A(n_0), .B1(n_2), .B2(n_1), .ZN(p_0));
   NOR2_X1 i_1 (.A1(to_int6126[6]), .A2(to_int6126[5]), .ZN(n_0));
   NAND2_X1 i_2 (.A1(to_int6126[4]), .A2(to_int6126[3]), .ZN(n_1));
   AOI21_X1 i_3 (.A(to_int6126[2]), .B1(to_int6126[1]), .B2(to_int6126[0]), 
      .ZN(n_2));
endmodule

module datapath__1_13610(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   OR3_X1 i_0 (.A1(to_int6126[6]), .A2(to_int6126[5]), .A3(n_0), .ZN(p_0));
   AND3_X1 i_1 (.A1(to_int6126[3]), .A2(n_1), .A3(to_int6126[4]), .ZN(n_0));
   OR3_X1 i_2 (.A1(to_int6126[1]), .A2(to_int6126[0]), .A3(to_int6126[2]), 
      .ZN(n_1));
endmodule

module datapath__1_13602(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NAND2_X1 i_0 (.A1(n_1), .A2(n_0), .ZN(p_0));
   NOR2_X1 i_1 (.A1(to_int6126[6]), .A2(to_int6126[5]), .ZN(n_0));
   OAI21_X1 i_2 (.A(to_int6126[4]), .B1(to_int6126[3]), .B2(n_2), .ZN(n_1));
   AND3_X1 i_3 (.A1(to_int6126[2]), .A2(to_int6126[1]), .A3(to_int6126[0]), 
      .ZN(n_2));
endmodule

module datapath__1_13594(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   OAI21_X1 i_0 (.A(to_int6126[2]), .B1(to_int6126[1]), .B2(to_int6126[0]), 
      .ZN(n_0));
   INV_X1 i_1 (.A(n_0), .ZN(n_1));
   OAI21_X1 i_2 (.A(to_int6126[4]), .B1(n_1), .B2(to_int6126[3]), .ZN(n_2));
   NOR2_X1 i_3 (.A1(to_int6126[6]), .A2(to_int6126[5]), .ZN(n_3));
   NAND2_X1 i_4 (.A1(n_2), .A2(n_3), .ZN(p_0));
endmodule

module datapath__1_13586(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   OAI21_X1 i_0 (.A(n_0), .B1(n_2), .B2(n_1), .ZN(p_0));
   NOR2_X1 i_1 (.A1(to_int6126[6]), .A2(to_int6126[5]), .ZN(n_0));
   AOI211_X1 i_2 (.A(to_int6126[2]), .B(to_int6126[3]), .C1(to_int6126[1]), 
      .C2(to_int6126[0]), .ZN(n_1));
   INV_X1 i_3 (.A(to_int6126[4]), .ZN(n_2));
endmodule

module datapath__1_13578(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   OAI21_X1 i_0 (.A(n_0), .B1(n_2), .B2(n_1), .ZN(p_0));
   NOR2_X1 i_1 (.A1(to_int6126[6]), .A2(to_int6126[5]), .ZN(n_0));
   NOR4_X1 i_2 (.A1(to_int6126[2]), .A2(to_int6126[0]), .A3(to_int6126[3]), 
      .A4(to_int6126[1]), .ZN(n_1));
   INV_X1 i_3 (.A(to_int6126[4]), .ZN(n_2));
endmodule

module datapath__1_13562(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NAND2_X1 i_0 (.A1(n_3), .A2(n_0), .ZN(p_0));
   NOR3_X1 i_1 (.A1(to_int6126[5]), .A2(to_int6126[4]), .A3(n_1), .ZN(n_0));
   INV_X1 i_2 (.A(n_2), .ZN(n_1));
   OAI211_X1 i_3 (.A(to_int6126[3]), .B(to_int6126[2]), .C1(to_int6126[1]), 
      .C2(to_int6126[0]), .ZN(n_2));
   INV_X1 i_4 (.A(to_int6126[6]), .ZN(n_3));
endmodule

module datapath__1_13538(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NAND2_X1 i_0 (.A1(n_3), .A2(n_0), .ZN(p_0));
   NOR4_X1 i_1 (.A1(to_int6126[5]), .A2(to_int6126[4]), .A3(to_int6126[3]), 
      .A4(n_1), .ZN(n_0));
   INV_X1 i_2 (.A(n_2), .ZN(n_1));
   NAND3_X1 i_3 (.A1(to_int6126[2]), .A2(to_int6126[1]), .A3(to_int6126[0]), 
      .ZN(n_2));
   INV_X1 i_4 (.A(to_int6126[6]), .ZN(n_3));
endmodule

module datapath__1_13997(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NOR2_X1 i_0 (.A1(n_1), .A2(n_0), .ZN(p_0));
   OAI211_X1 i_1 (.A(to_int6126[4]), .B(to_int6126[3]), .C1(to_int6126[2]), 
      .C2(to_int6126[1]), .ZN(n_0));
   NAND2_X1 i_2 (.A1(to_int6126[6]), .A2(to_int6126[5]), .ZN(n_1));
endmodule

module datapath__1_13949(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0));
   OAI211_X1 i_1 (.A(to_int6126[6]), .B(to_int6126[5]), .C1(to_int6126[4]), 
      .C2(n_1), .ZN(n_0));
   AND3_X1 i_2 (.A1(to_int6126[3]), .A2(to_int6126[2]), .A3(to_int6126[1]), 
      .ZN(n_1));
endmodule

module datapath__1_13901(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   AND3_X1 i_0 (.A1(to_int6126[6]), .A2(to_int6126[5]), .A3(n_0), .ZN(p_0));
   OR4_X1 i_1 (.A1(to_int6126[3]), .A2(to_int6126[1]), .A3(to_int6126[4]), 
      .A4(to_int6126[2]), .ZN(n_0));
endmodule

module datapath__1_13885(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0));
   OAI21_X1 i_1 (.A(to_int6126[6]), .B1(to_int6126[5]), .B2(n_1), .ZN(n_0));
   AND4_X1 i_2 (.A1(to_int6126[4]), .A2(to_int6126[3]), .A3(to_int6126[2]), 
      .A4(to_int6126[1]), .ZN(n_1));
endmodule

module datapath__1_13869(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0));
   OAI21_X1 i_1 (.A(to_int6126[6]), .B1(to_int6126[5]), .B2(n_1), .ZN(n_0));
   INV_X1 i_2 (.A(n_2), .ZN(n_1));
   OAI211_X1 i_3 (.A(to_int6126[4]), .B(to_int6126[3]), .C1(to_int6126[2]), 
      .C2(to_int6126[1]), .ZN(n_2));
endmodule

module datapath__1_13853(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NOR2_X1 i_0 (.A1(n_3), .A2(n_0), .ZN(p_0));
   AOI21_X1 i_1 (.A(to_int6126[5]), .B1(to_int6126[4]), .B2(n_1), .ZN(n_0));
   INV_X1 i_2 (.A(n_2), .ZN(n_1));
   AOI21_X1 i_3 (.A(to_int6126[3]), .B1(to_int6126[2]), .B2(to_int6126[1]), 
      .ZN(n_2));
   INV_X1 i_4 (.A(to_int6126[6]), .ZN(n_3));
endmodule

module datapath__1_13837(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NOR2_X1 i_0 (.A1(n_2), .A2(n_0), .ZN(p_0));
   AOI21_X1 i_1 (.A(to_int6126[5]), .B1(to_int6126[4]), .B2(n_1), .ZN(n_0));
   OR3_X1 i_2 (.A1(to_int6126[2]), .A2(to_int6126[1]), .A3(to_int6126[3]), 
      .ZN(n_1));
   INV_X1 i_3 (.A(to_int6126[6]), .ZN(n_2));
endmodule

module datapath__1_13821(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   AND3_X1 i_0 (.A1(to_int6126[2]), .A2(to_int6126[1]), .A3(to_int6126[3]), 
      .ZN(n_0));
   OR3_X1 i_1 (.A1(n_0), .A2(to_int6126[4]), .A3(to_int6126[5]), .ZN(n_1));
   AND2_X1 i_2 (.A1(n_1), .A2(to_int6126[6]), .ZN(p_0));
endmodule

module datapath__1_13805(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NOR2_X1 i_0 (.A1(n_2), .A2(n_0), .ZN(p_0));
   AOI211_X1 i_1 (.A(to_int6126[5]), .B(to_int6126[4]), .C1(to_int6126[3]), 
      .C2(n_1), .ZN(n_0));
   OR2_X1 i_2 (.A1(to_int6126[2]), .A2(to_int6126[1]), .ZN(n_1));
   INV_X1 i_3 (.A(to_int6126[6]), .ZN(n_2));
endmodule

module datapath__1_13789(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   AOI21_X1 i_0 (.A(n_2), .B1(n_1), .B2(n_0), .ZN(p_0));
   NOR3_X1 i_1 (.A1(to_int6126[5]), .A2(to_int6126[3]), .A3(to_int6126[4]), 
      .ZN(n_0));
   NAND2_X1 i_2 (.A1(to_int6126[2]), .A2(to_int6126[1]), .ZN(n_1));
   INV_X1 i_3 (.A(to_int6126[6]), .ZN(n_2));
endmodule

module datapath__1_13773(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0));
   OAI21_X1 i_1 (.A(to_int6126[6]), .B1(to_int6126[2]), .B2(n_1), .ZN(n_0));
   OR4_X1 i_2 (.A1(to_int6126[5]), .A2(to_int6126[4]), .A3(to_int6126[3]), 
      .A4(to_int6126[1]), .ZN(n_1));
endmodule

module datapath__1_13758(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NAND4_X1 i_0 (.A1(to_int6126[3]), .A2(to_int6126[4]), .A3(to_int6126[2]), 
      .A4(to_int6126[1]), .ZN(n_0));
   NAND2_X1 i_1 (.A1(n_3), .A2(n_1), .ZN(p_0));
   NAND2_X1 i_2 (.A1(n_2), .A2(to_int6126[5]), .ZN(n_1));
   INV_X1 i_3 (.A(n_0), .ZN(n_2));
   INV_X1 i_4 (.A(to_int6126[6]), .ZN(n_3));
endmodule

module datapath__1_13742(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   OAI21_X1 i_0 (.A(n_2), .B1(n_1), .B2(n_0), .ZN(p_0));
   NAND3_X1 i_1 (.A1(to_int6126[5]), .A2(to_int6126[3]), .A3(to_int6126[4]), 
      .ZN(n_0));
   NOR2_X1 i_2 (.A1(to_int6126[2]), .A2(to_int6126[1]), .ZN(n_1));
   INV_X1 i_3 (.A(to_int6126[6]), .ZN(n_2));
endmodule

module datapath__1_13726(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   OAI21_X1 i_0 (.A(n_2), .B1(n_1), .B2(n_0), .ZN(p_0));
   NAND2_X1 i_1 (.A1(to_int6126[5]), .A2(to_int6126[4]), .ZN(n_0));
   AOI21_X1 i_2 (.A(to_int6126[3]), .B1(to_int6126[2]), .B2(to_int6126[1]), 
      .ZN(n_1));
   INV_X1 i_3 (.A(to_int6126[6]), .ZN(n_2));
endmodule

module datapath__1_13710(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   OR2_X1 i_0 (.A1(to_int6126[6]), .A2(n_0), .ZN(p_0));
   AND3_X1 i_1 (.A1(to_int6126[4]), .A2(n_1), .A3(to_int6126[5]), .ZN(n_0));
   OR3_X1 i_2 (.A1(to_int6126[2]), .A2(to_int6126[1]), .A3(to_int6126[3]), 
      .ZN(n_1));
endmodule

module datapath__1_13694(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NAND2_X1 i_0 (.A1(n_2), .A2(n_0), .ZN(p_0));
   OAI21_X1 i_1 (.A(to_int6126[5]), .B1(to_int6126[4]), .B2(n_1), .ZN(n_0));
   AND3_X1 i_2 (.A1(to_int6126[2]), .A2(to_int6126[1]), .A3(to_int6126[3]), 
      .ZN(n_1));
   INV_X1 i_3 (.A(to_int6126[6]), .ZN(n_2));
endmodule

module datapath__1_13678(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NAND2_X1 i_0 (.A1(n_3), .A2(n_0), .ZN(p_0));
   OAI21_X1 i_1 (.A(to_int6126[5]), .B1(to_int6126[4]), .B2(n_1), .ZN(n_0));
   INV_X1 i_2 (.A(n_2), .ZN(n_1));
   OAI21_X1 i_3 (.A(to_int6126[3]), .B1(to_int6126[2]), .B2(to_int6126[1]), 
      .ZN(n_2));
   INV_X1 i_4 (.A(to_int6126[6]), .ZN(n_3));
endmodule

module datapath__1_13662(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   OAI21_X1 i_0 (.A(n_2), .B1(n_1), .B2(n_0), .ZN(p_0));
   AOI211_X1 i_1 (.A(to_int6126[3]), .B(to_int6126[4]), .C1(to_int6126[2]), 
      .C2(to_int6126[1]), .ZN(n_0));
   INV_X1 i_2 (.A(to_int6126[5]), .ZN(n_1));
   INV_X1 i_3 (.A(to_int6126[6]), .ZN(n_2));
endmodule

module datapath__1_13646(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NAND2_X1 i_0 (.A1(n_2), .A2(n_0), .ZN(p_0));
   OAI21_X1 i_1 (.A(to_int6126[5]), .B1(to_int6126[4]), .B2(n_1), .ZN(n_0));
   OR3_X1 i_2 (.A1(to_int6126[3]), .A2(to_int6126[2]), .A3(to_int6126[1]), 
      .ZN(n_1));
   INV_X1 i_3 (.A(to_int6126[6]), .ZN(n_2));
endmodule

module datapath__1_13614(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NAND2_X1 i_0 (.A1(n_1), .A2(n_0), .ZN(p_0));
   NOR2_X1 i_1 (.A1(to_int6126[6]), .A2(to_int6126[5]), .ZN(n_0));
   OAI211_X1 i_2 (.A(to_int6126[4]), .B(to_int6126[3]), .C1(to_int6126[2]), 
      .C2(to_int6126[1]), .ZN(n_1));
endmodule

module datapath__1_13598(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   OAI21_X1 i_0 (.A(n_0), .B1(n_2), .B2(n_1), .ZN(p_0));
   NOR2_X1 i_1 (.A1(to_int6126[6]), .A2(to_int6126[5]), .ZN(n_0));
   AOI21_X1 i_2 (.A(to_int6126[3]), .B1(to_int6126[2]), .B2(to_int6126[1]), 
      .ZN(n_1));
   INV_X1 i_3 (.A(to_int6126[4]), .ZN(n_2));
endmodule

module datapath__1_13582(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   OAI21_X1 i_0 (.A(n_0), .B1(n_2), .B2(n_1), .ZN(p_0));
   NOR2_X1 i_1 (.A1(to_int6126[6]), .A2(to_int6126[5]), .ZN(n_0));
   NOR3_X1 i_2 (.A1(to_int6126[2]), .A2(to_int6126[1]), .A3(to_int6126[3]), 
      .ZN(n_1));
   INV_X1 i_3 (.A(to_int6126[4]), .ZN(n_2));
endmodule

module datapath__1_13566(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NAND2_X1 i_0 (.A1(n_3), .A2(n_0), .ZN(p_0));
   NOR3_X1 i_1 (.A1(to_int6126[5]), .A2(to_int6126[4]), .A3(n_1), .ZN(n_0));
   INV_X1 i_2 (.A(n_2), .ZN(n_1));
   NAND3_X1 i_3 (.A1(to_int6126[3]), .A2(to_int6126[2]), .A3(to_int6126[1]), 
      .ZN(n_2));
   INV_X1 i_4 (.A(to_int6126[6]), .ZN(n_3));
endmodule

module datapath__1_13550(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NAND2_X1 i_0 (.A1(n_2), .A2(n_0), .ZN(p_0));
   AOI211_X1 i_1 (.A(to_int6126[4]), .B(to_int6126[5]), .C1(to_int6126[3]), 
      .C2(n_1), .ZN(n_0));
   OR2_X1 i_2 (.A1(to_int6126[2]), .A2(to_int6126[1]), .ZN(n_1));
   INV_X1 i_3 (.A(to_int6126[6]), .ZN(n_2));
endmodule

module datapath__1_13534(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NAND2_X1 i_0 (.A1(n_1), .A2(n_0), .ZN(p_0));
   AOI211_X1 i_1 (.A(to_int6126[5]), .B(to_int6126[4]), .C1(to_int6126[2]), 
      .C2(to_int6126[1]), .ZN(n_0));
   NOR2_X1 i_2 (.A1(to_int6126[6]), .A2(to_int6126[3]), .ZN(n_1));
endmodule

module datapath__1_13519(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NAND2_X1 i_0 (.A1(n_1), .A2(n_0), .ZN(p_0));
   NOR4_X1 i_1 (.A1(to_int6126[6]), .A2(to_int6126[5]), .A3(to_int6126[4]), 
      .A4(to_int6126[1]), .ZN(n_0));
   NOR2_X1 i_2 (.A1(to_int6126[3]), .A2(to_int6126[2]), .ZN(n_1));
endmodule

module datapath__1_13909(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   AND3_X1 i_0 (.A1(to_int6126[5]), .A2(n_0), .A3(to_int6126[6]), .ZN(p_0));
   OR3_X1 i_1 (.A1(to_int6126[3]), .A2(to_int6126[2]), .A3(to_int6126[4]), 
      .ZN(n_0));
endmodule

module datapath__1_13877(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0));
   OAI21_X1 i_1 (.A(to_int6126[6]), .B1(to_int6126[5]), .B2(n_1), .ZN(n_0));
   AND3_X1 i_2 (.A1(to_int6126[4]), .A2(to_int6126[3]), .A3(to_int6126[2]), 
      .ZN(n_1));
endmodule

module datapath__1_13845(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0));
   NAND2_X1 i_1 (.A1(to_int6126[6]), .A2(n_1), .ZN(n_0));
   NAND2_X1 i_2 (.A1(n_2), .A2(n_3), .ZN(n_1));
   OAI21_X1 i_3 (.A(to_int6126[4]), .B1(to_int6126[3]), .B2(to_int6126[2]), 
      .ZN(n_2));
   INV_X1 i_4 (.A(to_int6126[5]), .ZN(n_3));
endmodule

module datapath__1_13813(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0));
   OAI21_X1 i_1 (.A(to_int6126[6]), .B1(to_int6126[5]), .B2(n_1), .ZN(n_0));
   INV_X1 i_2 (.A(n_2), .ZN(n_1));
   AOI21_X1 i_3 (.A(to_int6126[4]), .B1(to_int6126[3]), .B2(to_int6126[2]), 
      .ZN(n_2));
endmodule

module datapath__1_13781(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0));
   OAI21_X1 i_1 (.A(to_int6126[6]), .B1(to_int6126[3]), .B2(n_1), .ZN(n_0));
   OR3_X1 i_2 (.A1(to_int6126[4]), .A2(to_int6126[2]), .A3(to_int6126[5]), 
      .ZN(n_1));
endmodule

module datapath__1_13750(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NAND2_X1 i_0 (.A1(n_1), .A2(n_0), .ZN(p_0));
   NAND4_X1 i_1 (.A1(to_int6126[5]), .A2(to_int6126[4]), .A3(to_int6126[3]), 
      .A4(to_int6126[2]), .ZN(n_0));
   INV_X1 i_2 (.A(to_int6126[6]), .ZN(n_1));
endmodule

module datapath__1_13718(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NAND2_X1 i_0 (.A1(n_1), .A2(n_0), .ZN(p_0));
   OAI211_X1 i_1 (.A(to_int6126[5]), .B(to_int6126[4]), .C1(to_int6126[3]), 
      .C2(to_int6126[2]), .ZN(n_0));
   INV_X1 i_2 (.A(to_int6126[6]), .ZN(n_1));
endmodule

module datapath__1_13686(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   OAI21_X1 i_0 (.A(n_2), .B1(n_1), .B2(n_0), .ZN(p_0));
   AOI21_X1 i_1 (.A(to_int6126[4]), .B1(to_int6126[3]), .B2(to_int6126[2]), 
      .ZN(n_0));
   INV_X1 i_2 (.A(to_int6126[5]), .ZN(n_1));
   INV_X1 i_3 (.A(to_int6126[6]), .ZN(n_2));
endmodule

module datapath__1_13654(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NAND2_X1 i_0 (.A1(n_2), .A2(n_0), .ZN(p_0));
   OAI21_X1 i_1 (.A(to_int6126[5]), .B1(to_int6126[4]), .B2(n_1), .ZN(n_0));
   OR2_X1 i_2 (.A1(to_int6126[3]), .A2(to_int6126[2]), .ZN(n_1));
   INV_X1 i_3 (.A(to_int6126[6]), .ZN(n_2));
endmodule

module datapath__1_13622(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NAND2_X1 i_0 (.A1(n_3), .A2(n_0), .ZN(p_0));
   NOR2_X1 i_1 (.A1(to_int6126[5]), .A2(n_1), .ZN(n_0));
   INV_X1 i_2 (.A(n_2), .ZN(n_1));
   NAND3_X1 i_3 (.A1(to_int6126[4]), .A2(to_int6126[3]), .A3(to_int6126[2]), 
      .ZN(n_2));
   INV_X1 i_4 (.A(to_int6126[6]), .ZN(n_3));
endmodule

module datapath__1_13590(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   OAI21_X1 i_0 (.A(to_int6126[4]), .B1(to_int6126[3]), .B2(to_int6126[2]), 
      .ZN(n_0));
   NOR2_X1 i_1 (.A1(to_int6126[6]), .A2(to_int6126[5]), .ZN(n_1));
   NAND2_X1 i_2 (.A1(n_0), .A2(n_1), .ZN(p_0));
endmodule

module datapath__1_13558(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NAND2_X1 i_0 (.A1(n_3), .A2(n_0), .ZN(p_0));
   NOR3_X1 i_1 (.A1(to_int6126[5]), .A2(to_int6126[4]), .A3(n_1), .ZN(n_0));
   INV_X1 i_2 (.A(n_2), .ZN(n_1));
   NAND2_X1 i_3 (.A1(to_int6126[3]), .A2(to_int6126[2]), .ZN(n_2));
   INV_X1 i_4 (.A(to_int6126[6]), .ZN(n_3));
endmodule

module datapath__1_13526(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   OR4_X1 i_0 (.A1(to_int6126[4]), .A2(to_int6126[2]), .A3(to_int6126[5]), 
      .A4(to_int6126[3]), .ZN(n_0));
   OR2_X1 i_1 (.A1(n_0), .A2(to_int6126[6]), .ZN(p_0));
endmodule

module datapath__1_13925(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0));
   OAI211_X1 i_1 (.A(to_int6126[6]), .B(to_int6126[5]), .C1(to_int6126[4]), 
      .C2(to_int6126[3]), .ZN(n_0));
endmodule

module datapath__1_13861(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NOR2_X1 i_0 (.A1(n_1), .A2(n_0), .ZN(p_0));
   AOI21_X1 i_1 (.A(to_int6126[5]), .B1(to_int6126[4]), .B2(to_int6126[3]), 
      .ZN(n_0));
   INV_X1 i_2 (.A(to_int6126[6]), .ZN(n_1));
endmodule

module datapath__1_13797(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   OR3_X1 i_0 (.A1(to_int6126[4]), .A2(to_int6126[3]), .A3(to_int6126[5]), 
      .ZN(n_0));
   AND2_X1 i_1 (.A1(n_0), .A2(to_int6126[6]), .ZN(p_0));
endmodule

module datapath__1_13734(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   INV_X1 i_0 (.A(to_int6126[6]), .ZN(n_0));
   NAND3_X1 i_1 (.A1(to_int6126[4]), .A2(to_int6126[5]), .A3(to_int6126[3]), 
      .ZN(n_1));
   NAND2_X1 i_2 (.A1(n_1), .A2(n_0), .ZN(p_0));
endmodule

module datapath__1_13670(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NAND2_X1 i_0 (.A1(n_1), .A2(n_0), .ZN(p_0));
   OAI21_X1 i_1 (.A(to_int6126[5]), .B1(to_int6126[4]), .B2(to_int6126[3]), 
      .ZN(n_0));
   INV_X1 i_2 (.A(to_int6126[6]), .ZN(n_1));
endmodule

module datapath__1_13606(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NAND2_X1 i_0 (.A1(n_1), .A2(n_0), .ZN(p_0));
   AOI21_X1 i_1 (.A(to_int6126[5]), .B1(to_int6126[4]), .B2(to_int6126[3]), 
      .ZN(n_0));
   INV_X1 i_2 (.A(to_int6126[6]), .ZN(n_1));
endmodule

module datapath__1_13542(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NAND2_X1 i_0 (.A1(n_1), .A2(n_0), .ZN(p_0));
   NOR3_X1 i_1 (.A1(to_int6126[5]), .A2(to_int6126[4]), .A3(to_int6126[3]), 
      .ZN(n_0));
   INV_X1 i_2 (.A(to_int6126[6]), .ZN(n_1));
endmodule

module datapath__1_13702(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NAND2_X1 i_0 (.A1(n_1), .A2(n_0), .ZN(p_0));
   NAND2_X1 i_1 (.A1(to_int6126[5]), .A2(to_int6126[4]), .ZN(n_0));
   INV_X1 i_2 (.A(to_int6126[6]), .ZN(n_1));
endmodule

module datapath__1_13893(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   AND2_X1 i_0 (.A1(to_int6126[6]), .A2(to_int6126[5]), .ZN(p_0));
endmodule

module half_adder__3_82(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   INV_X1 i_2 (.A(a), .ZN(f));
endmodule

module half_adder__3_85(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_88(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(f));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(n_0_1), .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(a), .A2(b), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_3), .A2(n_0_4), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(a), .ZN(n_0_3));
   INV_X1 i_0_6 (.A(b), .ZN(n_0_4));
endmodule

module half_adder__3_91(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;

   INV_X1 i_0_0 (.A(n_0_0), .ZN(f));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(n_0_4), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(n_0_3), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(a), .ZN(n_0_2));
   INV_X1 i_0_4 (.A(b), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(n_0_4), .ZN(cout));
   NAND2_X1 i_0_6 (.A1(a), .A2(b), .ZN(n_0_4));
endmodule

module half_adder__3_94(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_0_0;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   INV_X1 i_0_0 (.A(n_0_0), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(n_0_0));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(a), .A2(b), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_3), .A2(n_1_4), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module half_adder__3_97(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(b), .A2(a), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_4), .A2(n_1_3), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module half_adder(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_4), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(b), .A2(a), .ZN(n_1_1));
   INV_X1 i_1_3 (.A(a), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(b), .ZN(n_1_3));
   NAND2_X1 i_1_5 (.A1(n_1_2), .A2(n_1_3), .ZN(n_1_4));
endmodule

module incrementor(a, enbl, c);
   input [6:0]a;
   input enbl;
   output [6:0]c;

   half_adder__3_82 half_adder_0_0_half_adder_0_i (.a(a[0]), .b(), .cout(), 
      .f(c[0]));
   half_adder__3_85 half_adder_0_1_half_adder_0_i (.a(a[1]), .b(a[0]), .cout(n_0), 
      .f(c[1]));
   half_adder__3_88 half_adder_0_2_half_adder_0_i (.a(a[2]), .b(n_0), .cout(n_1), 
      .f(c[2]));
   half_adder__3_91 half_adder_0_3_half_adder_0_i (.a(a[3]), .b(n_1), .cout(n_2), 
      .f(c[3]));
   half_adder__3_94 half_adder_0_4_half_adder_0_i (.a(a[4]), .b(n_2), .cout(n_3), 
      .f(c[4]));
   half_adder__3_97 half_adder_0_5_half_adder_0_i (.a(a[5]), .b(n_3), .cout(n_4), 
      .f(c[5]));
   half_adder half_adder_0_6_half_adder_0_i (.a(a[6]), .b(n_4), .cout(), 
      .f(c[6]));
endmodule

module full_adder__3_3(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(f));
   AND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(cout));
endmodule

module full_adder__3_7(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   NOR2_X1 i_0_0 (.A1(n_0_1), .A2(n_0_0), .ZN(f));
   AOI21_X1 i_0_1 (.A(cin), .B1(n_0_3), .B2(n_0_5), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_2), .ZN(n_0_1));
   NAND3_X1 i_0_3 (.A1(n_0_3), .A2(cin), .A3(n_0_5), .ZN(n_0_2));
   INV_X1 i_0_4 (.A(n_0_4), .ZN(n_0_3));
   OAI21_X1 i_0_5 (.A(n_0_5), .B1(n_0_4), .B2(n_0_6), .ZN(cout));
   NOR2_X1 i_0_6 (.A1(a), .A2(b), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(a), .A2(b), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(cin), .ZN(n_0_6));
endmodule

module full_adder__3_11(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   INV_X1 i_0_1 (.A(n_0_0), .ZN(f));
   NAND2_X1 i_0_2 (.A1(n_0_1), .A2(n_0_3), .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(n_0_2), .A2(n_0_5), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(cin), .ZN(n_0_2));
   NAND2_X1 i_0_0 (.A1(n_0_3), .A2(n_0_9), .ZN(cout));
   NAND2_X1 i_0_5 (.A1(cin), .A2(n_0_4), .ZN(n_0_3));
   INV_X1 i_0_6 (.A(n_0_5), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_9), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(n_0_7), .A2(n_0_8), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(a), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(b), .ZN(n_0_8));
   NAND2_X1 i_0_11 (.A1(a), .A2(b), .ZN(n_0_9));
endmodule

module full_adder__3_15(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;

   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(f));
   NAND2_X1 i_0_2 (.A1(cin), .A2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_3), .A2(a), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(cin), .ZN(n_0_3));
endmodule

module full_adder__3_19(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__3_23(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;

   INV_X1 i_0_0 (.A(n_0_1), .ZN(cout));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(f));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(n_0_1), .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(cin), .A2(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_3), .A2(n_0_4), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(cin), .ZN(n_0_3));
   INV_X1 i_0_6 (.A(a), .ZN(n_0_4));
endmodule

module full_adder__3_27(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(f));
   NAND2_X1 i_0_1 (.A1(a), .A2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(n_0_3), .A2(cin), .ZN(n_0_2));
   INV_X1 i_0_4 (.A(a), .ZN(n_0_3));
endmodule

module int_adder(a, b, cin, enbl, c, cout);
   input [6:0]a;
   input [2:0]b;
   input cin;
   input enbl;
   output [6:0]c;
   output cout;

   full_adder__3_3 full_adder_0_0_full_adder_0_i (.a(a[0]), .b(b[0]), .cin(), 
      .f(c[0]), .cout(n_0));
   full_adder__3_7 full_adder_0_1_full_adder_0_i (.a(a[1]), .b(b[1]), .cin(n_0), 
      .f(c[1]), .cout(n_1));
   full_adder__3_11 full_adder_0_2_full_adder_0_i (.a(a[2]), .b(b[2]), .cin(n_1), 
      .f(c[2]), .cout(n_2));
   full_adder__3_15 full_adder_0_3_full_adder_0_i (.a(a[3]), .b(), .cin(n_2), 
      .f(c[3]), .cout(n_3));
   full_adder__3_19 full_adder_0_4_full_adder_0_i (.a(a[4]), .b(), .cin(n_3), 
      .f(c[4]), .cout(n_4));
   full_adder__3_23 full_adder_0_5_full_adder_0_i (.a(a[5]), .b(), .cin(n_4), 
      .f(c[5]), .cout(n_5));
   full_adder__3_27 full_adder_0_6_full_adder_0_i (.a(a[6]), .b(), .cin(n_5), 
      .f(c[6]), .cout());
endmodule

module range_extractor(in_a, in_size, out_a, out_b);
   input [6:0]in_a;
   input [2:0]in_size;
   output [6:0]out_a;
   output [6:0]out_b;

   incrementor inc (.a(in_a), .enbl(), .c(out_a));
   int_adder add (.a(out_a), .b(in_size), .cin(), .enbl(), .c(out_b), .cout());
endmodule

module datapath__1_7663(\out_as[6] , \out_bs[6] , p_0);
   input [6:0]\out_as[6] ;
   input [6:0]\out_bs[6] ;
   output p_0;

   OAI21_X1 i_0 (.A(n_23), .B1(n_22), .B2(n_0), .ZN(p_0));
   NOR2_X1 i_1 (.A1(n_1), .A2(n_19), .ZN(n_0));
   AOI21_X1 i_2 (.A(n_2), .B1(n_18), .B2(\out_as[6] [5]), .ZN(n_1));
   NAND2_X1 i_3 (.A1(n_3), .A2(n_16), .ZN(n_2));
   OAI21_X1 i_4 (.A(n_4), .B1(n_17), .B2(\out_as[6] [4]), .ZN(n_3));
   AOI21_X1 i_5 (.A(n_5), .B1(n_15), .B2(\out_bs[6] [3]), .ZN(n_4));
   AOI21_X1 i_6 (.A(n_6), .B1(n_14), .B2(\out_as[6] [3]), .ZN(n_5));
   OAI21_X1 i_7 (.A(n_7), .B1(n_13), .B2(\out_bs[6] [2]), .ZN(n_6));
   NAND3_X1 i_8 (.A1(n_12), .A2(n_10), .A3(n_8), .ZN(n_7));
   OAI22_X1 i_9 (.A1(\out_bs[6] [1]), .A2(n_11), .B1(n_9), .B2(\out_bs[6] [0]), 
      .ZN(n_8));
   INV_X1 i_10 (.A(\out_as[6] [0]), .ZN(n_9));
   NAND2_X1 i_11 (.A1(\out_bs[6] [1]), .A2(n_11), .ZN(n_10));
   INV_X1 i_12 (.A(\out_as[6] [1]), .ZN(n_11));
   NAND2_X1 i_13 (.A1(\out_bs[6] [2]), .A2(n_13), .ZN(n_12));
   INV_X1 i_14 (.A(\out_as[6] [2]), .ZN(n_13));
   INV_X1 i_15 (.A(\out_bs[6] [3]), .ZN(n_14));
   INV_X1 i_16 (.A(\out_as[6] [3]), .ZN(n_15));
   NAND2_X1 i_17 (.A1(n_17), .A2(\out_as[6] [4]), .ZN(n_16));
   INV_X1 i_18 (.A(\out_bs[6] [4]), .ZN(n_17));
   INV_X1 i_19 (.A(\out_bs[6] [5]), .ZN(n_18));
   INV_X1 i_20 (.A(n_20), .ZN(n_19));
   NAND2_X1 i_21 (.A1(\out_bs[6] [5]), .A2(n_21), .ZN(n_20));
   INV_X1 i_22 (.A(\out_as[6] [5]), .ZN(n_21));
   NOR2_X1 i_23 (.A1(\out_bs[6] [6]), .A2(n_24), .ZN(n_22));
   NAND2_X1 i_24 (.A1(\out_bs[6] [6]), .A2(n_24), .ZN(n_23));
   INV_X1 i_25 (.A(\out_as[6] [6]), .ZN(n_24));
endmodule

module datapath__1_12443(\out_as[7] , \out_bs[7] , p_0);
   input [6:0]\out_as[7] ;
   input [6:0]\out_bs[7] ;
   output p_0;

   INV_X1 i_2 (.A(\out_as[7] [6]), .ZN(n_0));
   INV_X1 i_18 (.A(n_18), .ZN(n_17));
   OAI21_X1 i_19 (.A(n_19), .B1(n_23), .B2(\out_bs[7] [2]), .ZN(n_18));
   NAND2_X1 i_20 (.A1(n_22), .A2(\out_as[7] [1]), .ZN(n_19));
   OAI211_X1 i_21 (.A(\out_as[7] [0]), .B(n_21), .C1(n_22), .C2(\out_as[7] [1]), 
      .ZN(n_20));
   INV_X1 i_22 (.A(\out_bs[7] [0]), .ZN(n_21));
   INV_X1 i_23 (.A(\out_bs[7] [1]), .ZN(n_22));
   INV_X1 i_24 (.A(\out_as[7] [2]), .ZN(n_23));
   NAND2_X1 i_17 (.A1(\out_bs[7] [2]), .A2(n_23), .ZN(n_1));
   NAND2_X1 i_25 (.A1(n_17), .A2(n_20), .ZN(n_2));
   NAND2_X1 i_0 (.A1(n_4), .A2(n_3), .ZN(p_0));
   OR2_X1 i_1 (.A1(n_6), .A2(\out_as[7] [6]), .ZN(n_3));
   NAND2_X1 i_3 (.A1(\out_bs[7] [6]), .A2(n_5), .ZN(n_4));
   NAND2_X1 i_4 (.A1(n_6), .A2(n_16), .ZN(n_5));
   AOI22_X1 i_5 (.A1(n_7), .A2(n_9), .B1(n_15), .B2(\out_bs[7] [5]), .ZN(n_6));
   AOI22_X1 i_6 (.A1(n_8), .A2(\out_as[7] [5]), .B1(\out_as[7] [4]), .B2(n_14), 
      .ZN(n_7));
   INV_X1 i_7 (.A(\out_bs[7] [5]), .ZN(n_8));
   OAI211_X1 i_8 (.A(n_11), .B(n_10), .C1(n_14), .C2(\out_as[7] [4]), .ZN(n_9));
   NAND2_X1 i_9 (.A1(\out_bs[7] [3]), .A2(n_13), .ZN(n_10));
   OAI21_X1 i_10 (.A(n_12), .B1(n_13), .B2(\out_bs[7] [3]), .ZN(n_11));
   NAND2_X1 i_11 (.A1(n_2), .A2(n_1), .ZN(n_12));
   INV_X1 i_12 (.A(\out_as[7] [3]), .ZN(n_13));
   INV_X1 i_13 (.A(\out_bs[7] [4]), .ZN(n_14));
   INV_X1 i_14 (.A(\out_as[7] [5]), .ZN(n_15));
   INV_X1 i_15 (.A(n_0), .ZN(n_16));
endmodule

module datapath__1_14009(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NOR2_X1 i_0 (.A1(n_1), .A2(n_0), .ZN(p_0));
   OAI21_X1 i_1 (.A(to_int6126[3]), .B1(to_int6126[1]), .B2(to_int6126[0]), 
      .ZN(n_0));
   NAND4_X1 i_2 (.A1(to_int6126[6]), .A2(to_int6126[5]), .A3(to_int6126[4]), 
      .A4(to_int6126[2]), .ZN(n_1));
endmodule

module datapath__1_13993(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NAND4_X1 i_3 (.A1(to_int6126[5]), .A2(to_int6126[4]), .A3(to_int6126[3]), 
      .A4(n_0), .ZN(n_2));
   OR3_X1 i_4 (.A1(to_int6126[2]), .A2(to_int6126[1]), .A3(to_int6126[0]), 
      .ZN(n_0));
   INV_X1 i_0 (.A(to_int6126[6]), .ZN(n_1));
   NOR2_X1 i_1 (.A1(n_1), .A2(n_2), .ZN(p_0));
endmodule

module datapath__1_13977(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0));
   NAND2_X1 i_1 (.A1(to_int6126[6]), .A2(n_1), .ZN(n_0));
   INV_X1 i_2 (.A(n_2), .ZN(n_1));
   OAI211_X1 i_3 (.A(to_int6126[5]), .B(to_int6126[4]), .C1(to_int6126[3]), 
      .C2(n_3), .ZN(n_2));
   INV_X1 i_4 (.A(n_4), .ZN(n_3));
   OAI21_X1 i_5 (.A(to_int6126[2]), .B1(to_int6126[1]), .B2(to_int6126[0]), 
      .ZN(n_4));
endmodule

module datapath__1_13969(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NOR2_X1 i_0 (.A1(n_1), .A2(n_0), .ZN(p_0));
   NAND3_X1 i_1 (.A1(to_int6126[5]), .A2(to_int6126[4]), .A3(to_int6126[6]), 
      .ZN(n_0));
   AOI211_X1 i_2 (.A(to_int6126[2]), .B(to_int6126[3]), .C1(to_int6126[1]), 
      .C2(to_int6126[0]), .ZN(n_1));
endmodule

module datapath__1_13921(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   AND3_X1 i_0 (.A1(to_int6126[5]), .A2(n_0), .A3(to_int6126[6]), .ZN(p_0));
   OR3_X1 i_1 (.A1(to_int6126[3]), .A2(n_1), .A3(to_int6126[4]), .ZN(n_0));
   AND3_X1 i_2 (.A1(to_int6126[1]), .A2(to_int6126[0]), .A3(to_int6126[2]), 
      .ZN(n_1));
endmodule

module datapath__1_14013(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0));
   NAND2_X1 i_1 (.A1(to_int6126[6]), .A2(n_1), .ZN(n_0));
   INV_X1 i_2 (.A(n_2), .ZN(n_1));
   NAND3_X1 i_3 (.A1(to_int6126[5]), .A2(to_int6126[4]), .A3(n_3), .ZN(n_2));
   INV_X1 i_4 (.A(n_4), .ZN(n_3));
   NAND3_X1 i_5 (.A1(to_int6126[3]), .A2(to_int6126[2]), .A3(to_int6126[1]), 
      .ZN(n_4));
endmodule

module datapath__1_13981(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NOR2_X1 i_0 (.A1(n_1), .A2(n_0), .ZN(p_0));
   NAND3_X1 i_1 (.A1(to_int6126[5]), .A2(to_int6126[4]), .A3(to_int6126[6]), 
      .ZN(n_0));
   AOI21_X1 i_2 (.A(to_int6126[3]), .B1(to_int6126[2]), .B2(to_int6126[1]), 
      .ZN(n_1));
endmodule

module datapath__1_13965(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   AND4_X1 i_0 (.A1(to_int6126[5]), .A2(to_int6126[4]), .A3(to_int6126[6]), 
      .A4(n_0), .ZN(p_0));
   OR3_X1 i_1 (.A1(to_int6126[2]), .A2(to_int6126[1]), .A3(to_int6126[3]), 
      .ZN(n_0));
endmodule

module datapath__1_13933(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   AOI21_X1 i_0 (.A(n_0), .B1(n_2), .B2(n_1), .ZN(p_0));
   NAND2_X1 i_1 (.A1(to_int6126[6]), .A2(to_int6126[5]), .ZN(n_0));
   OAI21_X1 i_2 (.A(to_int6126[3]), .B1(to_int6126[2]), .B2(to_int6126[1]), 
      .ZN(n_1));
   INV_X1 i_3 (.A(to_int6126[4]), .ZN(n_2));
endmodule

module datapath__1_13917(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   AOI211_X1 i_0 (.A(to_int6126[3]), .B(to_int6126[4]), .C1(to_int6126[2]), 
      .C2(to_int6126[1]), .ZN(n_0));
   NAND2_X1 i_1 (.A1(to_int6126[6]), .A2(to_int6126[5]), .ZN(n_1));
   NOR2_X1 i_2 (.A1(n_1), .A2(n_0), .ZN(p_0));
endmodule

module datapath__1_14005(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   AND4_X1 i_0 (.A1(to_int6126[5]), .A2(to_int6126[4]), .A3(to_int6126[3]), 
      .A4(to_int6126[2]), .ZN(n_0));
   AND2_X1 i_1 (.A1(n_0), .A2(to_int6126[6]), .ZN(p_0));
endmodule

module datapath__1_13973(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   AND4_X1 i_0 (.A1(to_int6126[5]), .A2(to_int6126[4]), .A3(n_0), .A4(
      to_int6126[6]), .ZN(p_0));
   OR2_X1 i_1 (.A1(to_int6126[3]), .A2(to_int6126[2]), .ZN(n_0));
endmodule

module datapath__1_13941(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   AOI21_X1 i_0 (.A(to_int6126[4]), .B1(to_int6126[3]), .B2(to_int6126[2]), 
      .ZN(n_0));
   NAND2_X1 i_1 (.A1(to_int6126[6]), .A2(to_int6126[5]), .ZN(n_1));
   NOR2_X1 i_2 (.A1(n_1), .A2(n_0), .ZN(p_0));
endmodule

module datapath__1_13989(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NAND3_X1 i_0 (.A1(to_int6126[5]), .A2(to_int6126[4]), .A3(to_int6126[3]), 
      .ZN(n_0));
   INV_X1 i_1 (.A(to_int6126[6]), .ZN(n_1));
   NOR2_X1 i_2 (.A1(n_1), .A2(n_0), .ZN(p_0));
endmodule

module datapath__1_13957(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   AND3_X1 i_0 (.A1(to_int6126[6]), .A2(to_int6126[4]), .A3(to_int6126[5]), 
      .ZN(p_0));
endmodule

module datapath__1_13829(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   OAI21_X1 i_0 (.A(to_int6126[6]), .B1(to_int6126[5]), .B2(to_int6126[4]), 
      .ZN(n_0));
   INV_X1 i_1 (.A(n_0), .ZN(p_0));
endmodule

module datapath__1_13638(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   OR2_X1 i_0 (.A1(to_int6126[6]), .A2(to_int6126[5]), .ZN(p_0));
endmodule

module datapath__1_13765(to_int6128, p_0);
   input [7:0]to_int6128;
   output p_0;

   HA_X1 i_0 (.A(to_int6128[6]), .B(n_1), .CO(n_0), .S());
   NAND2_X1 i_1 (.A1(n_3), .A2(n_2), .ZN(n_1));
   NOR4_X1 i_2 (.A1(to_int6128[5]), .A2(to_int6128[4]), .A3(to_int6128[3]), 
      .A4(to_int6128[0]), .ZN(n_2));
   NOR2_X1 i_3 (.A1(to_int6128[2]), .A2(to_int6128[1]), .ZN(n_3));
   INV_X1 i_4 (.A(n_0), .ZN(p_0));
endmodule

module datapath__1_13509(\out_as[5] , \out_bs[5] , p_0);
   input [6:0]\out_as[5] ;
   input [6:0]\out_bs[5] ;
   output p_0;

   OAI21_X1 i_0 (.A(n_22), .B1(n_21), .B2(n_0), .ZN(p_0));
   INV_X1 i_1 (.A(n_1), .ZN(n_0));
   OAI21_X1 i_2 (.A(n_19), .B1(n_18), .B2(n_2), .ZN(n_1));
   NAND2_X1 i_3 (.A1(n_3), .A2(n_16), .ZN(n_2));
   OAI211_X1 i_4 (.A(n_15), .B(n_13), .C1(n_12), .C2(n_4), .ZN(n_3));
   OAI21_X1 i_5 (.A(n_5), .B1(n_11), .B2(\out_bs[5] [2]), .ZN(n_4));
   NAND3_X1 i_6 (.A1(n_10), .A2(n_8), .A3(n_6), .ZN(n_5));
   OAI22_X1 i_7 (.A1(\out_bs[5] [1]), .A2(n_9), .B1(n_7), .B2(\out_bs[5] [0]), 
      .ZN(n_6));
   INV_X1 i_8 (.A(\out_as[5] [0]), .ZN(n_7));
   NAND2_X1 i_9 (.A1(\out_bs[5] [1]), .A2(n_9), .ZN(n_8));
   INV_X1 i_10 (.A(\out_as[5] [1]), .ZN(n_9));
   NAND2_X1 i_11 (.A1(\out_bs[5] [2]), .A2(n_11), .ZN(n_10));
   INV_X1 i_12 (.A(\out_as[5] [2]), .ZN(n_11));
   NOR2_X1 i_13 (.A1(\out_bs[5] [3]), .A2(n_14), .ZN(n_12));
   NAND2_X1 i_14 (.A1(\out_bs[5] [3]), .A2(n_14), .ZN(n_13));
   INV_X1 i_15 (.A(\out_as[5] [3]), .ZN(n_14));
   NAND2_X1 i_16 (.A1(\out_bs[5] [4]), .A2(n_17), .ZN(n_15));
   OR2_X1 i_17 (.A1(\out_bs[5] [4]), .A2(n_17), .ZN(n_16));
   INV_X1 i_18 (.A(\out_as[5] [4]), .ZN(n_17));
   NOR2_X1 i_19 (.A1(\out_bs[5] [5]), .A2(n_20), .ZN(n_18));
   NAND2_X1 i_20 (.A1(\out_bs[5] [5]), .A2(n_20), .ZN(n_19));
   INV_X1 i_21 (.A(\out_as[5] [5]), .ZN(n_20));
   NOR2_X1 i_22 (.A1(\out_bs[5] [6]), .A2(n_23), .ZN(n_21));
   NAND2_X1 i_23 (.A1(\out_bs[5] [6]), .A2(n_23), .ZN(n_22));
   INV_X1 i_24 (.A(\out_as[5] [6]), .ZN(n_23));
endmodule

module half_adder__3_147(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   INV_X1 i_2 (.A(a), .ZN(f));
endmodule

module half_adder__3_144(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   AND2_X1 i_0_0 (.A1(b), .A2(a), .ZN(cout));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(b), .A2(a), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_4), .A2(n_1_3), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module half_adder__3_141(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_0_0;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   INV_X1 i_0_0 (.A(n_0_0), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(n_0_0));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_1), .A2(n_1_4), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(n_1_3), .A2(n_1_2), .ZN(n_1_1));
   INV_X1 i_1_3 (.A(a), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(b), .ZN(n_1_3));
   NAND2_X1 i_1_5 (.A1(b), .A2(a), .ZN(n_1_4));
endmodule

module half_adder__3_138(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;

   INV_X1 i_0_0 (.A(n_0_0), .ZN(f));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(n_0_4), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_3), .A2(n_0_2), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(a), .ZN(n_0_2));
   INV_X1 i_0_4 (.A(b), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(n_0_4), .ZN(cout));
   NAND2_X1 i_0_6 (.A1(b), .A2(a), .ZN(n_0_4));
endmodule

module half_adder__3_135(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   AND2_X1 i_0_0 (.A1(b), .A2(a), .ZN(cout));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(b), .A2(a), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_4), .A2(n_1_3), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module half_adder__3_132(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   AND2_X1 i_0_0 (.A1(b), .A2(a), .ZN(cout));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(b), .A2(a), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_4), .A2(n_1_3), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module half_adder__3_129(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(b), .A2(a), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_4), .A2(n_1_3), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module incrementor__3_148(a, enbl, c);
   input [6:0]a;
   input enbl;
   output [6:0]c;

   half_adder__3_147 half_adder_0_0_half_adder_0_i (.a(a[0]), .b(), .cout(), 
      .f(c[0]));
   half_adder__3_144 half_adder_0_1_half_adder_0_i (.a(a[1]), .b(a[0]), .cout(
      n_0), .f(c[1]));
   half_adder__3_141 half_adder_0_2_half_adder_0_i (.a(a[2]), .b(n_0), .cout(n_1), 
      .f(c[2]));
   half_adder__3_138 half_adder_0_3_half_adder_0_i (.a(a[3]), .b(n_1), .cout(n_2), 
      .f(c[3]));
   half_adder__3_135 half_adder_0_4_half_adder_0_i (.a(a[4]), .b(n_2), .cout(n_3), 
      .f(c[4]));
   half_adder__3_132 half_adder_0_5_half_adder_0_i (.a(a[5]), .b(n_3), .cout(n_4), 
      .f(c[5]));
   half_adder__3_129 half_adder_0_6_half_adder_0_i (.a(a[6]), .b(n_4), .cout(), 
      .f(c[6]));
endmodule

module full_adder__3_125(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;

   INV_X1 i_0_0 (.A(n_0_0), .ZN(f));
   NAND2_X1 i_0_1 (.A1(n_0_2), .A2(n_0_1), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(b), .A2(a), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(n_0_4), .A2(n_0_3), .ZN(n_0_2));
   INV_X1 i_0_4 (.A(a), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(b), .ZN(n_0_4));
   AND2_X1 i_1_0 (.A1(b), .A2(a), .ZN(cout));
endmodule

module full_adder__3_121(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_3;
   wire n_0_1;
   wire n_0_8;
   wire n_0_9;
   wire n_0_4;
   wire n_0_5;
   wire n_0_15;
   wire n_0_16;
   wire n_0_6;
   wire n_0_7;
   wire n_0_11;
   wire n_0_12;
   wire n_0_10;
   wire n_0_13;
   wire n_0_14;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(f));
   NAND2_X1 i_0_1 (.A1(n_0_16), .A2(cin), .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(n_0_3), .A2(n_0_9), .ZN(n_0_2));
   INV_X1 i_0_4 (.A(cin), .ZN(n_0_3));
   NAND2_X1 i_0_2 (.A1(n_0_7), .A2(n_0_1), .ZN(cout));
   NAND2_X1 i_0_5 (.A1(b), .A2(a), .ZN(n_0_1));
   INV_X1 i_0_6 (.A(b), .ZN(n_0_8));
   NAND2_X1 i_0_7 (.A1(n_0_4), .A2(n_0_13), .ZN(n_0_9));
   NAND2_X1 i_0_8 (.A1(n_0_8), .A2(a), .ZN(n_0_4));
   INV_X1 i_0_15 (.A(b), .ZN(n_0_5));
   NOR2_X1 i_0_9 (.A1(a), .A2(n_0_5), .ZN(n_0_15));
   OAI21_X1 i_0_10 (.A(n_0_14), .B1(n_0_15), .B2(n_0_8), .ZN(n_0_16));
   NAND2_X1 i_0_14 (.A1(n_0_10), .A2(n_0_4), .ZN(n_0_6));
   NAND2_X1 i_0_16 (.A1(n_0_6), .A2(cin), .ZN(n_0_7));
   INV_X1 i_0_11 (.A(a), .ZN(n_0_11));
   INV_X1 i_0_12 (.A(a), .ZN(n_0_12));
   NAND2_X1 i_0_13 (.A1(b), .A2(n_0_11), .ZN(n_0_10));
   NAND2_X1 i_0_17 (.A1(b), .A2(n_0_12), .ZN(n_0_13));
   NAND2_X1 i_0_18 (.A1(n_0_12), .A2(n_0_5), .ZN(n_0_14));
endmodule

module full_adder__3_117(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_1_1;
   wire n_1_2;
   wire n_1_4;
   wire n_1_5;
   wire n_1_6;
   wire n_1_0;
   wire n_1_3;

   NAND2_X1 i_0_0 (.A1(n_0), .A2(cin), .ZN(n_0_0));
   NAND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(n_0_1));
   NAND2_X1 i_0_2 (.A1(n_0_0), .A2(n_0_1), .ZN(cout));
   INV_X1 i_1_7 (.A(b), .ZN(n_1_1));
   INV_X1 i_1_6 (.A(n_1_1), .ZN(n_1_2));
   OAI21_X1 i_1_0 (.A(n_1_5), .B1(a), .B2(n_1_2), .ZN(n_1_4));
   OAI21_X1 i_1_1 (.A(n_1_3), .B1(cin), .B2(n_1_4), .ZN(f));
   NAND2_X1 i_1_2 (.A1(a), .A2(n_1_2), .ZN(n_1_5));
   INV_X1 i_1_5 (.A(n_1_2), .ZN(n_1_6));
   XNOR2_X1 i_1_8 (.A(n_1_6), .B(a), .ZN(n_0));
   XNOR2_X1 i_1_3 (.A(a), .B(b), .ZN(n_1_0));
   NAND2_X1 i_1_4 (.A1(n_1_0), .A2(cin), .ZN(n_1_3));
endmodule

module full_adder__3_113(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_1_0;

   INV_X1 i_0_4 (.A(a), .ZN(n_0_0));
   OAI21_X1 i_0_0 (.A(n_0_1), .B1(cin), .B2(n_0_2), .ZN(f));
   NAND2_X1 i_0_1 (.A1(cin), .A2(n_0_0), .ZN(n_0_1));
   INV_X1 i_0_2 (.A(a), .ZN(n_0_2));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(cout));
   NAND2_X1 i_1_1 (.A1(cin), .A2(a), .ZN(n_1_0));
endmodule

module full_adder__3_109(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_1_0;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(f));
   NAND2_X1 i_0_1 (.A1(a), .A2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(n_0_3), .A2(cin), .ZN(n_0_2));
   INV_X1 i_0_4 (.A(a), .ZN(n_0_3));
   NAND2_X1 i_1_0 (.A1(a), .A2(cin), .ZN(n_1_0));
   INV_X1 i_1_1 (.A(n_1_0), .ZN(cout));
endmodule

module full_adder__3_105(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_1_0;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_2), .ZN(f));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(a), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(cin), .A2(n_0_3), .ZN(n_0_2));
   INV_X1 i_0_4 (.A(a), .ZN(n_0_3));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(cout));
   NAND2_X1 i_1_1 (.A1(cin), .A2(a), .ZN(n_1_0));
endmodule

module full_adder__3_101(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(f));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(cin), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(a), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(n_0_3), .A2(a), .ZN(n_0_2));
   INV_X1 i_0_4 (.A(cin), .ZN(n_0_3));
endmodule

module int_adder__3_126(a, b, cin, enbl, c, cout);
   input [6:0]a;
   input [2:0]b;
   input cin;
   input enbl;
   output [6:0]c;
   output cout;

   full_adder__3_125 full_adder_0_0_full_adder_0_i (.a(a[0]), .b(b[0]), .cin(), 
      .f(c[0]), .cout(n_0));
   full_adder__3_121 full_adder_0_1_full_adder_0_i (.a(a[1]), .b(b[1]), .cin(n_0), 
      .f(c[1]), .cout(n_1));
   full_adder__3_117 full_adder_0_2_full_adder_0_i (.a(a[2]), .b(b[2]), .cin(n_1), 
      .f(c[2]), .cout(n_2));
   full_adder__3_113 full_adder_0_3_full_adder_0_i (.a(a[3]), .b(), .cin(n_2), 
      .f(c[3]), .cout(n_3));
   full_adder__3_109 full_adder_0_4_full_adder_0_i (.a(a[4]), .b(), .cin(n_3), 
      .f(c[4]), .cout(n_4));
   full_adder__3_105 full_adder_0_5_full_adder_0_i (.a(a[5]), .b(), .cin(n_4), 
      .f(c[5]), .cout(n_5));
   full_adder__3_101 full_adder_0_6_full_adder_0_i (.a(a[6]), .b(), .cin(n_5), 
      .f(c[6]), .cout());
endmodule

module range_extractor__3_149(in_a, in_size, out_a, out_b);
   input [6:0]in_a;
   input [2:0]in_size;
   output [6:0]out_a;
   output [6:0]out_b;

   incrementor__3_148 inc (.a(in_a), .enbl(), .c(out_a));
   int_adder__3_126 add (.a(out_a), .b(in_size), .cin(), .enbl(), .c(out_b), 
      .cout());
endmodule

module half_adder__3_199(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   INV_X1 i_2 (.A(a), .ZN(f));
endmodule

module half_adder__3_196(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_0_0;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   INV_X1 i_0_0 (.A(n_0_0), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(n_0_0));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(a), .A2(b), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_3), .A2(n_1_4), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module half_adder__3_193(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_0_0;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   INV_X1 i_0_0 (.A(n_0_0), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(n_0_0));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(b), .A2(a), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_4), .A2(n_1_3), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module half_adder__3_190(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_0_0;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   INV_X1 i_0_0 (.A(n_0_0), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(n_0_0));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(a), .A2(b), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_3), .A2(n_1_4), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module half_adder__3_187(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_0_0;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   INV_X1 i_0_0 (.A(n_0_0), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(n_0_0));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(a), .A2(b), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_3), .A2(n_1_4), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module half_adder__3_184(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   AND2_X1 i_0_0 (.A1(b), .A2(a), .ZN(cout));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(b), .A2(a), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_4), .A2(n_1_3), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module half_adder__3_181(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(b), .A2(a), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_4), .A2(n_1_3), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module incrementor__3_200(a, enbl, c);
   input [6:0]a;
   input enbl;
   output [6:0]c;

   half_adder__3_199 half_adder_0_0_half_adder_0_i (.a(a[0]), .b(), .cout(), 
      .f(c[0]));
   half_adder__3_196 half_adder_0_1_half_adder_0_i (.a(a[1]), .b(a[0]), .cout(
      n_0), .f(c[1]));
   half_adder__3_193 half_adder_0_2_half_adder_0_i (.a(a[2]), .b(n_0), .cout(n_1), 
      .f(c[2]));
   half_adder__3_190 half_adder_0_3_half_adder_0_i (.a(a[3]), .b(n_1), .cout(n_2), 
      .f(c[3]));
   half_adder__3_187 half_adder_0_4_half_adder_0_i (.a(a[4]), .b(n_2), .cout(n_3), 
      .f(c[4]));
   half_adder__3_184 half_adder_0_5_half_adder_0_i (.a(a[5]), .b(n_3), .cout(n_4), 
      .f(c[5]));
   half_adder__3_181 half_adder_0_6_half_adder_0_i (.a(a[6]), .b(n_4), .cout(), 
      .f(c[6]));
endmodule

module full_adder__3_177(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;

   INV_X1 i_0_0 (.A(n_0_0), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_3), .A2(n_0_1), .ZN(f));
   NAND2_X1 i_0_3 (.A1(a), .A2(n_0_2), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(b), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(n_0_4), .A2(b), .ZN(n_0_3));
   INV_X1 i_0_6 (.A(a), .ZN(n_0_4));
endmodule

module full_adder__3_173(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;
   wire n_1_5;
   wire n_1_6;
   wire n_1_7;
   wire n_1_8;
   wire n_1_9;

   NAND2_X1 i_0_0 (.A1(n_0_1), .A2(n_0_0), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(cin), .A2(b), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(a), .A2(n_0_2), .ZN(n_0_1));
   OR2_X1 i_0_3 (.A1(cin), .A2(b), .ZN(n_0_2));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_3), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(n_1_2), .A2(a), .ZN(n_1_1));
   INV_X1 i_1_3 (.A(n_1_4), .ZN(n_1_2));
   NAND2_X1 i_1_4 (.A1(n_1_9), .A2(n_1_4), .ZN(n_1_3));
   NAND2_X1 i_1_5 (.A1(n_1_6), .A2(n_1_5), .ZN(n_1_4));
   NAND2_X1 i_1_6 (.A1(cin), .A2(b), .ZN(n_1_5));
   NAND2_X1 i_1_7 (.A1(n_1_7), .A2(n_1_8), .ZN(n_1_6));
   INV_X1 i_1_8 (.A(cin), .ZN(n_1_7));
   INV_X1 i_1_9 (.A(b), .ZN(n_1_8));
   INV_X1 i_1_10 (.A(a), .ZN(n_1_9));
endmodule

module full_adder__3_169(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_5;
   wire n_0_6;
   wire n_0_2;
   wire n_0_8;
   wire n_0_4;
   wire n_0_3;
   wire n_0_7;
   wire n_0_9;
   wire n_0_10;

   NAND2_X1 i_0_0 (.A1(n_0_9), .A2(n_0_0), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(n_0_5), .A2(n_0_7), .ZN(f));
   NAND2_X1 i_0_2 (.A1(a), .A2(b), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(cin), .ZN(n_0_1));
   NAND3_X1 i_0_4 (.A1(n_0_8), .A2(cin), .A3(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_5 (.A1(a), .A2(n_0_2), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(b), .ZN(n_0_2));
   NAND2_X1 i_0_6 (.A1(n_0_4), .A2(b), .ZN(n_0_8));
   INV_X1 i_0_7 (.A(a), .ZN(n_0_4));
   NAND2_X1 i_0_8 (.A1(n_0_4), .A2(n_0_2), .ZN(n_0_3));
   NAND3_X1 i_0_10 (.A1(n_0_3), .A2(n_0_1), .A3(n_0_0), .ZN(n_0_7));
   NAND2_X1 i_0_11 (.A1(n_0_10), .A2(cin), .ZN(n_0_9));
   NAND2_X1 i_0_12 (.A1(n_0_4), .A2(n_0_2), .ZN(n_0_10));
endmodule

module full_adder__3_165(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_1_0;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_2), .ZN(f));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(a), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(cin), .A2(n_0_3), .ZN(n_0_2));
   INV_X1 i_0_4 (.A(a), .ZN(n_0_3));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(cout));
   NAND2_X1 i_1_1 (.A1(cin), .A2(a), .ZN(n_1_0));
endmodule

module full_adder__3_161(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_1_0;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_2), .ZN(f));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(a), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(cin), .A2(n_0_3), .ZN(n_0_2));
   INV_X1 i_0_4 (.A(a), .ZN(n_0_3));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(cout));
   NAND2_X1 i_1_1 (.A1(cin), .A2(a), .ZN(n_1_0));
endmodule

module full_adder__3_157(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_2), .ZN(f));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(a), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(cin), .A2(n_0_3), .ZN(n_0_2));
   INV_X1 i_0_4 (.A(a), .ZN(n_0_3));
   AND2_X1 i_1_0 (.A1(a), .A2(cin), .ZN(cout));
endmodule

module full_adder__3_153(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;

   NAND2_X1 i_0_0 (.A1(n_0_3), .A2(n_0_0), .ZN(f));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(cin), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(a), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(cin), .ZN(n_0_2));
   NAND2_X1 i_0_4 (.A1(a), .A2(n_0_2), .ZN(n_0_3));
endmodule

module int_adder__3_178(a, b, cin, enbl, c, cout);
   input [6:0]a;
   input [2:0]b;
   input cin;
   input enbl;
   output [6:0]c;
   output cout;

   full_adder__3_177 full_adder_0_0_full_adder_0_i (.a(a[0]), .b(b[0]), .cin(), 
      .f(c[0]), .cout(n_0));
   full_adder__3_173 full_adder_0_1_full_adder_0_i (.a(a[1]), .b(b[1]), .cin(n_0), 
      .f(c[1]), .cout(n_1));
   full_adder__3_169 full_adder_0_2_full_adder_0_i (.a(a[2]), .b(b[2]), .cin(n_1), 
      .f(c[2]), .cout(n_2));
   full_adder__3_165 full_adder_0_3_full_adder_0_i (.a(a[3]), .b(), .cin(n_2), 
      .f(c[3]), .cout(n_3));
   full_adder__3_161 full_adder_0_4_full_adder_0_i (.a(a[4]), .b(), .cin(n_3), 
      .f(c[4]), .cout(n_4));
   full_adder__3_157 full_adder_0_5_full_adder_0_i (.a(a[5]), .b(), .cin(n_4), 
      .f(c[5]), .cout(n_5));
   full_adder__3_153 full_adder_0_6_full_adder_0_i (.a(a[6]), .b(), .cin(n_5), 
      .f(c[6]), .cout());
endmodule

module range_extractor__3_201(in_a, in_size, out_a, out_b);
   input [6:0]in_a;
   input [2:0]in_size;
   output [6:0]out_a;
   output [6:0]out_b;

   incrementor__3_200 inc (.a(in_a), .enbl(), .c(out_a));
   int_adder__3_178 add (.a(out_a), .b(in_size), .cin(), .enbl(), .c(out_b), 
      .cout());
endmodule

module half_adder__3_251(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   INV_X1 i_2 (.A(a), .ZN(f));
endmodule

module half_adder__3_248(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_0_0;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   INV_X1 i_0_0 (.A(n_0_0), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(n_0_0));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(a), .A2(b), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_3), .A2(n_1_4), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module half_adder__3_245(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_0_0;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   NAND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(cout));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(a), .A2(b), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_3), .A2(n_1_4), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module half_adder__3_242(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_0_0;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   INV_X1 i_0_0 (.A(n_0_0), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(n_0_0));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(b), .A2(a), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_4), .A2(n_1_3), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module half_adder__3_239(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_0_0;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   INV_X1 i_0_0 (.A(n_0_0), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(n_0_0));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(b), .A2(a), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_4), .A2(n_1_3), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module half_adder__3_236(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   AND2_X1 i_0_0 (.A1(b), .A2(a), .ZN(cout));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(b), .A2(a), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_4), .A2(n_1_3), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module half_adder__3_233(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_4), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(b), .A2(a), .ZN(n_1_1));
   INV_X1 i_1_3 (.A(a), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(b), .ZN(n_1_3));
   NAND2_X1 i_1_5 (.A1(n_1_2), .A2(n_1_3), .ZN(n_1_4));
endmodule

module incrementor__3_252(a, enbl, c);
   input [6:0]a;
   input enbl;
   output [6:0]c;

   half_adder__3_251 half_adder_0_0_half_adder_0_i (.a(a[0]), .b(), .cout(), 
      .f(c[0]));
   half_adder__3_248 half_adder_0_1_half_adder_0_i (.a(a[1]), .b(a[0]), .cout(
      n_0), .f(c[1]));
   half_adder__3_245 half_adder_0_2_half_adder_0_i (.a(a[2]), .b(n_0), .cout(n_1), 
      .f(c[2]));
   half_adder__3_242 half_adder_0_3_half_adder_0_i (.a(a[3]), .b(n_1), .cout(n_2), 
      .f(c[3]));
   half_adder__3_239 half_adder_0_4_half_adder_0_i (.a(a[4]), .b(n_2), .cout(n_3), 
      .f(c[4]));
   half_adder__3_236 half_adder_0_5_half_adder_0_i (.a(a[5]), .b(n_3), .cout(n_4), 
      .f(c[5]));
   half_adder__3_233 half_adder_0_6_half_adder_0_i (.a(a[6]), .b(n_4), .cout(), 
      .f(c[6]));
endmodule

module full_adder__3_229(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(f));
   AND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(cout));
endmodule

module full_adder__3_225(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_2_0;
   wire n_2_1;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;

   NAND2_X1 i_2_0 (.A1(n_2_0), .A2(n_2_1), .ZN(cout));
   NAND2_X1 i_2_1 (.A1(n_0), .A2(cin), .ZN(n_2_0));
   NAND2_X1 i_2_2 (.A1(a), .A2(b), .ZN(n_2_1));
   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(f));
   NAND2_X1 i_0_1 (.A1(a), .A2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(n_0_5), .A2(n_0_3), .ZN(n_0_2));
   XNOR2_X1 i_0_4 (.A(cin), .B(n_0_4), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(b), .ZN(n_0_4));
   INV_X1 i_0_6 (.A(a), .ZN(n_0_5));
   NAND2_X1 i_1_0 (.A1(n_1_2), .A2(n_1_0), .ZN(n_0));
   NAND2_X1 i_1_1 (.A1(a), .A2(n_1_1), .ZN(n_1_0));
   INV_X1 i_1_2 (.A(b), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_3), .A2(b), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
endmodule

module full_adder__3_221(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_1_0;
   wire n_1_1;

   NAND2_X1 i_0_0 (.A1(n_0_1), .A2(n_0_0), .ZN(f));
   NAND3_X1 i_0_1 (.A1(n_0_5), .A2(n_0_3), .A3(cin), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(n_0_7), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(n_0_5), .A2(n_0_3), .ZN(n_0_2));
   NAND2_X1 i_0_4 (.A1(n_0_4), .A2(b), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(a), .ZN(n_0_4));
   NAND2_X1 i_0_6 (.A1(n_0_6), .A2(a), .ZN(n_0_5));
   INV_X1 i_0_7 (.A(b), .ZN(n_0_6));
   INV_X1 i_0_8 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_1_0 (.A1(n_1_1), .A2(n_1_0), .ZN(cout));
   NAND2_X1 i_1_1 (.A1(cin), .A2(b), .ZN(n_1_0));
   OAI21_X1 i_1_2 (.A(a), .B1(cin), .B2(b), .ZN(n_1_1));
endmodule

module full_adder__3_217(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_1_0;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_2), .ZN(f));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(a), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(cin), .A2(n_0_3), .ZN(n_0_2));
   INV_X1 i_0_4 (.A(a), .ZN(n_0_3));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(cout));
   NAND2_X1 i_1_1 (.A1(cin), .A2(a), .ZN(n_1_0));
endmodule

module full_adder__3_213(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_1_0;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(f));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(cin), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(a), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(n_0_3), .A2(a), .ZN(n_0_2));
   INV_X1 i_0_4 (.A(cin), .ZN(n_0_3));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(cout));
   NAND2_X1 i_1_1 (.A1(cin), .A2(a), .ZN(n_1_0));
endmodule

module full_adder__3_209(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(f));
   NAND2_X1 i_0_1 (.A1(a), .A2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(n_0_3), .A2(cin), .ZN(n_0_2));
   INV_X1 i_0_4 (.A(a), .ZN(n_0_3));
   AND2_X1 i_1_0 (.A1(a), .A2(cin), .ZN(cout));
endmodule

module full_adder__3_205(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;

   NAND2_X1 i_0_0 (.A1(n_0_3), .A2(n_0_0), .ZN(f));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(cin), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(a), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(cin), .ZN(n_0_2));
   NAND2_X1 i_0_4 (.A1(a), .A2(n_0_2), .ZN(n_0_3));
endmodule

module int_adder__3_230(a, b, cin, enbl, c, cout);
   input [6:0]a;
   input [2:0]b;
   input cin;
   input enbl;
   output [6:0]c;
   output cout;

   full_adder__3_229 full_adder_0_0_full_adder_0_i (.a(a[0]), .b(b[0]), .cin(), 
      .f(c[0]), .cout(n_0));
   full_adder__3_225 full_adder_0_1_full_adder_0_i (.a(a[1]), .b(b[1]), .cin(n_0), 
      .f(c[1]), .cout(n_1));
   full_adder__3_221 full_adder_0_2_full_adder_0_i (.a(a[2]), .b(b[2]), .cin(n_1), 
      .f(c[2]), .cout(n_2));
   full_adder__3_217 full_adder_0_3_full_adder_0_i (.a(a[3]), .b(), .cin(n_2), 
      .f(c[3]), .cout(n_3));
   full_adder__3_213 full_adder_0_4_full_adder_0_i (.a(a[4]), .b(), .cin(n_3), 
      .f(c[4]), .cout(n_4));
   full_adder__3_209 full_adder_0_5_full_adder_0_i (.a(a[5]), .b(), .cin(n_4), 
      .f(c[5]), .cout(n_5));
   full_adder__3_205 full_adder_0_6_full_adder_0_i (.a(a[6]), .b(), .cin(n_5), 
      .f(c[6]), .cout());
endmodule

module range_extractor__3_253(in_a, in_size, out_a, out_b);
   input [6:0]in_a;
   input [2:0]in_size;
   output [6:0]out_a;
   output [6:0]out_b;

   incrementor__3_252 inc (.a(in_a), .enbl(), .c(out_a));
   int_adder__3_230 add (.a(out_a), .b(in_size), .cin(), .enbl(), .c(out_b), 
      .cout());
endmodule

module half_adder__3_303(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   INV_X1 i_2 (.A(a), .ZN(f));
endmodule

module half_adder__3_300(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(b), .A2(a), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_4), .A2(n_1_3), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module half_adder__3_297(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_0_0;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   INV_X1 i_0_0 (.A(n_0_0), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(n_0_0));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(a), .A2(b), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_3), .A2(n_1_4), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module half_adder__3_294(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_0_0;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   INV_X1 i_0_0 (.A(n_0_0), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(a), .A2(b), .ZN(n_0_0));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(a), .A2(b), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_3), .A2(n_1_4), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module half_adder__3_291(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_0_0;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   INV_X1 i_0_0 (.A(n_0_0), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(n_0_0));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(b), .A2(a), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_4), .A2(n_1_3), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module half_adder__3_288(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;

   INV_X1 i_0_1 (.A(n_0_0), .ZN(f));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(n_0_1), .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(a), .A2(b), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_3), .A2(n_0_4), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(a), .ZN(n_0_3));
   INV_X1 i_0_6 (.A(b), .ZN(n_0_4));
   AND2_X1 i_0_0 (.A1(b), .A2(a), .ZN(cout));
endmodule

module half_adder__3_285(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(b), .A2(a), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_4), .A2(n_1_3), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module incrementor__3_304(a, enbl, c);
   input [6:0]a;
   input enbl;
   output [6:0]c;

   half_adder__3_303 half_adder_0_0_half_adder_0_i (.a(a[0]), .b(), .cout(), 
      .f(c[0]));
   half_adder__3_300 half_adder_0_1_half_adder_0_i (.a(a[1]), .b(a[0]), .cout(
      n_0), .f(c[1]));
   half_adder__3_297 half_adder_0_2_half_adder_0_i (.a(a[2]), .b(n_0), .cout(n_1), 
      .f(c[2]));
   half_adder__3_294 half_adder_0_3_half_adder_0_i (.a(a[3]), .b(n_1), .cout(n_2), 
      .f(c[3]));
   half_adder__3_291 half_adder_0_4_half_adder_0_i (.a(a[4]), .b(n_2), .cout(n_3), 
      .f(c[4]));
   half_adder__3_288 half_adder_0_5_half_adder_0_i (.a(a[5]), .b(n_3), .cout(n_4), 
      .f(c[5]));
   half_adder__3_285 half_adder_0_6_half_adder_0_i (.a(a[6]), .b(n_4), .cout(), 
      .f(c[6]));
endmodule

module full_adder__3_281(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(f));
   AND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(cout));
endmodule

module full_adder__3_277(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_2_0;
   wire n_2_1;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;

   NAND2_X1 i_2_0 (.A1(n_2_1), .A2(n_2_0), .ZN(cout));
   NAND2_X1 i_2_1 (.A1(a), .A2(b), .ZN(n_2_0));
   NAND2_X1 i_2_2 (.A1(n_0), .A2(cin), .ZN(n_2_1));
   INV_X1 i_0_8 (.A(b), .ZN(n_0_0));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_1));
   INV_X1 i_0_0 (.A(a), .ZN(n_0_2));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(b), .ZN(n_0_3));
   NAND2_X1 i_0_2 (.A1(cin), .A2(n_0_0), .ZN(n_0_4));
   NAND2_X1 i_0_3 (.A1(n_0_3), .A2(n_0_4), .ZN(n_0_5));
   NAND2_X1 i_0_4 (.A1(n_0_2), .A2(n_0_5), .ZN(n_0_6));
   NAND2_X1 i_0_5 (.A1(cin), .A2(b), .ZN(n_0_7));
   NAND2_X1 i_0_6 (.A1(n_0_10), .A2(n_0_7), .ZN(n_0_8));
   NAND2_X1 i_0_7 (.A1(n_0_8), .A2(a), .ZN(n_0_9));
   NAND2_X1 i_0_10 (.A1(n_0_6), .A2(n_0_9), .ZN(f));
   NAND2_X1 i_0_11 (.A1(n_0_1), .A2(n_0_0), .ZN(n_0_10));
   NAND2_X1 i_1_0 (.A1(n_1_2), .A2(n_1_0), .ZN(n_0));
   NAND2_X1 i_1_1 (.A1(a), .A2(n_1_1), .ZN(n_1_0));
   INV_X1 i_1_2 (.A(b), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_3), .A2(b), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
endmodule

module full_adder__3_273(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;

   INV_X1 i_0_0 (.A(n_0_0), .ZN(f));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(n_0_5), .ZN(n_0_0));
   NAND3_X1 i_0_2 (.A1(n_0_4), .A2(n_0_2), .A3(n_0_3), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(n_0_8), .A2(b), .ZN(n_0_2));
   NAND2_X1 i_0_4 (.A1(cin), .A2(n_0_9), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(a), .ZN(n_0_4));
   NAND3_X1 i_0_6 (.A1(n_0_7), .A2(a), .A3(n_0_6), .ZN(n_0_5));
   NAND2_X1 i_0_7 (.A1(cin), .A2(b), .ZN(n_0_6));
   NAND2_X1 i_0_8 (.A1(n_0_8), .A2(n_0_9), .ZN(n_0_7));
   INV_X1 i_0_9 (.A(cin), .ZN(n_0_8));
   INV_X1 i_0_10 (.A(b), .ZN(n_0_9));
   OAI21_X1 i_1_0 (.A(n_1_0), .B1(n_1_1), .B2(n_1_2), .ZN(cout));
   NAND2_X1 i_1_1 (.A1(cin), .A2(b), .ZN(n_1_0));
   NOR2_X1 i_1_2 (.A1(cin), .A2(b), .ZN(n_1_1));
   INV_X1 i_1_3 (.A(a), .ZN(n_1_2));
endmodule

module full_adder__3_269(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(f));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(a), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(n_0_3), .A2(cin), .ZN(n_0_2));
   INV_X1 i_0_4 (.A(a), .ZN(n_0_3));
   AND2_X1 i_1_0 (.A1(a), .A2(cin), .ZN(cout));
endmodule

module full_adder__3_265(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(f));
   NAND2_X1 i_0_1 (.A1(a), .A2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(n_0_3), .A2(cin), .ZN(n_0_2));
   INV_X1 i_0_4 (.A(a), .ZN(n_0_3));
   AND2_X1 i_1_0 (.A1(a), .A2(cin), .ZN(cout));
endmodule

module full_adder__3_261(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;

   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(f));
   NAND2_X1 i_0_2 (.A1(cin), .A2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_3), .A2(a), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(cin), .ZN(n_0_3));
endmodule

module full_adder__3_257(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(f));
   NAND2_X1 i_0_1 (.A1(a), .A2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(n_0_3), .A2(cin), .ZN(n_0_2));
   INV_X1 i_0_4 (.A(a), .ZN(n_0_3));
endmodule

module int_adder__3_282(a, b, cin, enbl, c, cout);
   input [6:0]a;
   input [2:0]b;
   input cin;
   input enbl;
   output [6:0]c;
   output cout;

   full_adder__3_281 full_adder_0_0_full_adder_0_i (.a(a[0]), .b(b[0]), .cin(), 
      .f(c[0]), .cout(n_0));
   full_adder__3_277 full_adder_0_1_full_adder_0_i (.a(a[1]), .b(b[1]), .cin(n_0), 
      .f(c[1]), .cout(n_1));
   full_adder__3_273 full_adder_0_2_full_adder_0_i (.a(a[2]), .b(b[2]), .cin(n_1), 
      .f(c[2]), .cout(n_2));
   full_adder__3_269 full_adder_0_3_full_adder_0_i (.a(a[3]), .b(), .cin(n_2), 
      .f(c[3]), .cout(n_3));
   full_adder__3_265 full_adder_0_4_full_adder_0_i (.a(a[4]), .b(), .cin(n_3), 
      .f(c[4]), .cout(n_4));
   full_adder__3_261 full_adder_0_5_full_adder_0_i (.a(a[5]), .b(), .cin(n_4), 
      .f(c[5]), .cout(n_5));
   full_adder__3_257 full_adder_0_6_full_adder_0_i (.a(a[6]), .b(), .cin(n_5), 
      .f(c[6]), .cout());
endmodule

module range_extractor__3_305(in_a, in_size, out_a, out_b);
   input [6:0]in_a;
   input [2:0]in_size;
   output [6:0]out_a;
   output [6:0]out_b;

   incrementor__3_304 inc (.a(in_a), .enbl(), .c(out_a));
   int_adder__3_282 add (.a(out_a), .b(in_size), .cin(), .enbl(), .c(out_b), 
      .cout());
endmodule

module half_adder__3_355(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   INV_X1 i_2 (.A(a), .ZN(f));
endmodule

module half_adder__3_352(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(a), .A2(b), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_3), .A2(n_1_4), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module half_adder__3_349(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_0_0;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   NAND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(cout));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(a), .A2(b), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_3), .A2(n_1_4), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module half_adder__3_346(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_0_0;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   INV_X1 i_0_0 (.A(n_0_0), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(n_0_0));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(b), .A2(a), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_4), .A2(n_1_3), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module half_adder__3_343(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   AND2_X1 i_0_0 (.A1(b), .A2(a), .ZN(cout));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(b), .A2(a), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_4), .A2(n_1_3), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module half_adder__3_340(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   AND2_X1 i_0_0 (.A1(b), .A2(a), .ZN(cout));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(b), .A2(a), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_4), .A2(n_1_3), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module half_adder__3_337(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_4), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(b), .A2(a), .ZN(n_1_1));
   INV_X1 i_1_3 (.A(a), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(b), .ZN(n_1_3));
   NAND2_X1 i_1_5 (.A1(n_1_2), .A2(n_1_3), .ZN(n_1_4));
endmodule

module incrementor__3_356(a, enbl, c);
   input [6:0]a;
   input enbl;
   output [6:0]c;

   half_adder__3_355 half_adder_0_0_half_adder_0_i (.a(a[0]), .b(), .cout(), 
      .f(c[0]));
   half_adder__3_352 half_adder_0_1_half_adder_0_i (.a(a[1]), .b(a[0]), .cout(
      n_0), .f(c[1]));
   half_adder__3_349 half_adder_0_2_half_adder_0_i (.a(a[2]), .b(n_0), .cout(n_1), 
      .f(c[2]));
   half_adder__3_346 half_adder_0_3_half_adder_0_i (.a(a[3]), .b(n_1), .cout(n_2), 
      .f(c[3]));
   half_adder__3_343 half_adder_0_4_half_adder_0_i (.a(a[4]), .b(n_2), .cout(n_3), 
      .f(c[4]));
   half_adder__3_340 half_adder_0_5_half_adder_0_i (.a(a[5]), .b(n_3), .cout(n_4), 
      .f(c[5]));
   half_adder__3_337 half_adder_0_6_half_adder_0_i (.a(a[6]), .b(n_4), .cout(), 
      .f(c[6]));
endmodule

module full_adder__3_333(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(f));
   AND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(cout));
endmodule

module full_adder__3_329(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_2_0;
   wire n_2_1;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(n_0));
   NAND2_X1 i_0_1 (.A1(a), .A2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(b), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(n_0_3), .A2(b), .ZN(n_0_2));
   INV_X1 i_0_4 (.A(a), .ZN(n_0_3));
   NAND2_X1 i_1_0 (.A1(n_1_2), .A2(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_0), .A2(n_1_1), .ZN(n_1_0));
   INV_X1 i_1_2 (.A(cin), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_3), .A2(cin), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(n_0), .ZN(n_1_3));
   NAND2_X1 i_2_0 (.A1(n_2_1), .A2(n_2_0), .ZN(cout));
   NAND2_X1 i_2_1 (.A1(a), .A2(b), .ZN(n_2_0));
   NAND2_X1 i_2_2 (.A1(n_0), .A2(cin), .ZN(n_2_1));
endmodule

module full_adder__3_325(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;
   wire n_1_5;
   wire n_1_6;
   wire n_1_7;

   OAI21_X1 i_0_0 (.A(a), .B1(cin), .B2(b), .ZN(n_0_0));
   NAND2_X1 i_0_1 (.A1(cin), .A2(b), .ZN(n_0_1));
   NAND2_X1 i_0_2 (.A1(n_0_0), .A2(n_0_1), .ZN(cout));
   NAND2_X1 i_1_0 (.A1(n_1_0), .A2(n_1_2), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_1), .A2(cin), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(n_1_4), .A2(n_1_3), .ZN(n_1_1));
   NAND3_X1 i_1_3 (.A1(n_1_4), .A2(n_1_7), .A3(n_1_3), .ZN(n_1_2));
   NAND2_X1 i_1_4 (.A1(a), .A2(b), .ZN(n_1_3));
   NAND2_X1 i_1_5 (.A1(n_1_6), .A2(n_1_5), .ZN(n_1_4));
   INV_X1 i_1_6 (.A(b), .ZN(n_1_5));
   INV_X1 i_1_7 (.A(a), .ZN(n_1_6));
   INV_X1 i_1_8 (.A(cin), .ZN(n_1_7));
endmodule

module full_adder__3_321(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_1_0;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_2), .ZN(f));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(a), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(cin), .A2(n_0_3), .ZN(n_0_2));
   INV_X1 i_0_4 (.A(a), .ZN(n_0_3));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(cout));
   NAND2_X1 i_1_1 (.A1(cin), .A2(a), .ZN(n_1_0));
endmodule

module full_adder__3_317(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;

   NAND2_X1 i_0_0 (.A1(n_0_0), .A2(n_0_2), .ZN(f));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(a), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(cin), .A2(n_0_3), .ZN(n_0_2));
   INV_X1 i_0_4 (.A(a), .ZN(n_0_3));
   AND2_X1 i_1_0 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__3_313(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;

   INV_X1 i_0_0 (.A(n_0_0), .ZN(f));
   NAND2_X1 i_0_1 (.A1(n_0_2), .A2(n_0_1), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(cin), .A2(a), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(n_0_4), .A2(n_0_3), .ZN(n_0_2));
   INV_X1 i_0_4 (.A(a), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(cin), .ZN(n_0_4));
   AND2_X1 i_1_0 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__3_309(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(f));
   NAND2_X1 i_0_1 (.A1(a), .A2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(n_0_3), .A2(cin), .ZN(n_0_2));
   INV_X1 i_0_4 (.A(a), .ZN(n_0_3));
endmodule

module int_adder__3_334(a, b, cin, enbl, c, cout);
   input [6:0]a;
   input [2:0]b;
   input cin;
   input enbl;
   output [6:0]c;
   output cout;

   full_adder__3_333 full_adder_0_0_full_adder_0_i (.a(a[0]), .b(b[0]), .cin(), 
      .f(c[0]), .cout(n_0));
   full_adder__3_329 full_adder_0_1_full_adder_0_i (.a(a[1]), .b(b[1]), .cin(n_0), 
      .f(c[1]), .cout(n_1));
   full_adder__3_325 full_adder_0_2_full_adder_0_i (.a(a[2]), .b(b[2]), .cin(n_1), 
      .f(c[2]), .cout(n_2));
   full_adder__3_321 full_adder_0_3_full_adder_0_i (.a(a[3]), .b(), .cin(n_2), 
      .f(c[3]), .cout(n_3));
   full_adder__3_317 full_adder_0_4_full_adder_0_i (.a(a[4]), .b(), .cin(n_3), 
      .f(c[4]), .cout(n_4));
   full_adder__3_313 full_adder_0_5_full_adder_0_i (.a(a[5]), .b(), .cin(n_4), 
      .f(c[5]), .cout(n_5));
   full_adder__3_309 full_adder_0_6_full_adder_0_i (.a(a[6]), .b(), .cin(n_5), 
      .f(c[6]), .cout());
endmodule

module range_extractor__3_357(in_a, in_size, out_a, out_b);
   input [6:0]in_a;
   input [2:0]in_size;
   output [6:0]out_a;
   output [6:0]out_b;

   incrementor__3_356 inc (.a(in_a), .enbl(), .c(out_a));
   int_adder__3_334 add (.a(out_a), .b(in_size), .cin(), .enbl(), .c(out_b), 
      .cout());
endmodule

module half_adder__3_407(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   INV_X1 i_2 (.A(a), .ZN(f));
endmodule

module half_adder__3_404(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(b), .A2(a), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_4), .A2(n_1_3), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module half_adder__3_401(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_0_0;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   NAND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(n_0_0));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(cout));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(a), .A2(b), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_3), .A2(n_1_4), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module half_adder__3_398(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_0_0;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   INV_X1 i_0_0 (.A(n_0_0), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(n_0_0));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(a), .A2(b), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_3), .A2(n_1_4), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module half_adder__3_395(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_0_0;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   INV_X1 i_0_0 (.A(n_0_0), .ZN(cout));
   NAND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(n_0_0));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(a), .A2(b), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_3), .A2(n_1_4), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module half_adder__3_392(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;
   wire n_1_4;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   INV_X1 i_1_0 (.A(n_1_0), .ZN(f));
   NAND2_X1 i_1_1 (.A1(n_1_2), .A2(n_1_1), .ZN(n_1_0));
   NAND2_X1 i_1_2 (.A1(a), .A2(b), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_3), .A2(n_1_4), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
   INV_X1 i_1_5 (.A(b), .ZN(n_1_4));
endmodule

module half_adder__3_389(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;

   INV_X1 i_1_0 (.A(b), .ZN(n_1_0));
   INV_X1 i_1_1 (.A(a), .ZN(n_1_1));
   NAND2_X1 i_1_2 (.A1(n_1_1), .A2(b), .ZN(n_1_2));
   NAND2_X1 i_1_3 (.A1(n_1_0), .A2(a), .ZN(n_1_3));
   NAND2_X1 i_1_4 (.A1(n_1_2), .A2(n_1_3), .ZN(f));
endmodule

module incrementor__3_408(a, enbl, c);
   input [6:0]a;
   input enbl;
   output [6:0]c;

   half_adder__3_407 half_adder_0_0_half_adder_0_i (.a(a[0]), .b(), .cout(), 
      .f(c[0]));
   half_adder__3_404 half_adder_0_1_half_adder_0_i (.a(a[1]), .b(a[0]), .cout(
      n_0), .f(c[1]));
   half_adder__3_401 half_adder_0_2_half_adder_0_i (.a(a[2]), .b(n_0), .cout(n_1), 
      .f(c[2]));
   half_adder__3_398 half_adder_0_3_half_adder_0_i (.a(a[3]), .b(n_1), .cout(n_2), 
      .f(c[3]));
   half_adder__3_395 half_adder_0_4_half_adder_0_i (.a(a[4]), .b(n_2), .cout(n_3), 
      .f(c[4]));
   half_adder__3_392 half_adder_0_5_half_adder_0_i (.a(a[5]), .b(n_3), .cout(n_4), 
      .f(c[5]));
   half_adder__3_389 half_adder_0_6_half_adder_0_i (.a(a[6]), .b(n_4), .cout(), 
      .f(c[6]));
endmodule

module full_adder__3_385(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(f));
   AND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(cout));
endmodule

module full_adder__3_381(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_2_0;
   wire n_2_1;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;

   NAND2_X1 i_2_0 (.A1(n_2_0), .A2(n_2_1), .ZN(cout));
   NAND2_X1 i_2_1 (.A1(cin), .A2(n_0), .ZN(n_2_0));
   NAND2_X1 i_2_2 (.A1(a), .A2(b), .ZN(n_2_1));
   NAND2_X1 i_0_0 (.A1(n_0_1), .A2(n_0_0), .ZN(f));
   NAND2_X1 i_0_1 (.A1(a), .A2(n_0_3), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_4), .A2(n_0_2), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(n_0_3), .ZN(n_0_2));
   XNOR2_X1 i_0_4 (.A(cin), .B(b), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(a), .ZN(n_0_4));
   NAND2_X1 i_1_0 (.A1(n_1_2), .A2(n_1_0), .ZN(n_0));
   NAND2_X1 i_1_1 (.A1(a), .A2(n_1_1), .ZN(n_1_0));
   INV_X1 i_1_2 (.A(b), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_3), .A2(b), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
endmodule

module full_adder__3_377(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_2_0;
   wire n_2_1;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_1_0;
   wire n_1_1;
   wire n_1_2;
   wire n_1_3;

   NAND2_X1 i_2_0 (.A1(n_2_0), .A2(n_2_1), .ZN(cout));
   NAND2_X1 i_2_1 (.A1(n_0), .A2(cin), .ZN(n_2_0));
   NAND2_X1 i_2_2 (.A1(a), .A2(b), .ZN(n_2_1));
   NAND2_X1 i_0_0 (.A1(n_0_1), .A2(n_0_0), .ZN(f));
   NAND3_X1 i_0_1 (.A1(n_0_5), .A2(n_0_3), .A3(cin), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(n_0_7), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(n_0_5), .A2(n_0_3), .ZN(n_0_2));
   NAND2_X1 i_0_4 (.A1(n_0_4), .A2(b), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(a), .ZN(n_0_4));
   NAND2_X1 i_0_6 (.A1(n_0_6), .A2(a), .ZN(n_0_5));
   INV_X1 i_0_7 (.A(b), .ZN(n_0_6));
   INV_X1 i_0_8 (.A(cin), .ZN(n_0_7));
   NAND2_X1 i_1_0 (.A1(n_1_2), .A2(n_1_0), .ZN(n_0));
   NAND2_X1 i_1_1 (.A1(a), .A2(n_1_1), .ZN(n_1_0));
   INV_X1 i_1_2 (.A(b), .ZN(n_1_1));
   NAND2_X1 i_1_3 (.A1(n_1_3), .A2(b), .ZN(n_1_2));
   INV_X1 i_1_4 (.A(a), .ZN(n_1_3));
endmodule

module full_adder__3_373(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;

   INV_X1 i_0_0 (.A(n_0_0), .ZN(f));
   NAND2_X1 i_0_1 (.A1(n_0_2), .A2(n_0_1), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(cin), .A2(a), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(n_0_4), .A2(n_0_3), .ZN(n_0_2));
   INV_X1 i_0_4 (.A(a), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(cin), .ZN(n_0_4));
   AND2_X1 i_1_0 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__3_369(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;

   INV_X1 i_0_0 (.A(n_0_0), .ZN(f));
   NAND2_X1 i_0_1 (.A1(n_0_2), .A2(n_0_1), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(cin), .A2(a), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(n_0_4), .A2(n_0_3), .ZN(n_0_2));
   INV_X1 i_0_4 (.A(a), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(cin), .ZN(n_0_4));
   AND2_X1 i_1_0 (.A1(a), .A2(cin), .ZN(cout));
endmodule

module full_adder__3_365(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;

   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
   INV_X1 i_0_0 (.A(n_0_0), .ZN(f));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(n_0_1), .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(cin), .A2(a), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_3), .A2(n_0_4), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(cin), .ZN(n_0_3));
   INV_X1 i_0_6 (.A(a), .ZN(n_0_4));
endmodule

module full_adder__3_361(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_0), .ZN(f));
   NAND2_X1 i_0_1 (.A1(a), .A2(n_0_1), .ZN(n_0_0));
   INV_X1 i_0_2 (.A(cin), .ZN(n_0_1));
   NAND2_X1 i_0_3 (.A1(n_0_3), .A2(cin), .ZN(n_0_2));
   INV_X1 i_0_4 (.A(a), .ZN(n_0_3));
endmodule

module int_adder__3_386(a, b, cin, enbl, c, cout);
   input [6:0]a;
   input [2:0]b;
   input cin;
   input enbl;
   output [6:0]c;
   output cout;

   full_adder__3_385 full_adder_0_0_full_adder_0_i (.a(a[0]), .b(b[0]), .cin(), 
      .f(c[0]), .cout(n_0));
   full_adder__3_381 full_adder_0_1_full_adder_0_i (.a(a[1]), .b(b[1]), .cin(n_0), 
      .f(c[1]), .cout(n_1));
   full_adder__3_377 full_adder_0_2_full_adder_0_i (.a(a[2]), .b(b[2]), .cin(n_1), 
      .f(c[2]), .cout(n_2));
   full_adder__3_373 full_adder_0_3_full_adder_0_i (.a(a[3]), .b(), .cin(n_2), 
      .f(c[3]), .cout(n_3));
   full_adder__3_369 full_adder_0_4_full_adder_0_i (.a(a[4]), .b(), .cin(n_3), 
      .f(c[4]), .cout(n_4));
   full_adder__3_365 full_adder_0_5_full_adder_0_i (.a(a[5]), .b(), .cin(n_4), 
      .f(c[5]), .cout(n_5));
   full_adder__3_361 full_adder_0_6_full_adder_0_i (.a(a[6]), .b(), .cin(n_5), 
      .f(c[6]), .cout());
endmodule

module range_extractor__3_409(in_a, in_size, out_a, out_b);
   input [6:0]in_a;
   input [2:0]in_size;
   output [6:0]out_a;
   output [6:0]out_b;

   incrementor__3_408 inc (.a(in_a), .enbl(), .c(out_a));
   int_adder__3_386 add (.a(out_a), .b(in_size), .cin(), .enbl(), .c(out_b), 
      .cout());
endmodule

module datapath__1_14044(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   NAND2_X1 i_0 (.A1(n_1), .A2(n_0), .ZN(p_0));
   NOR4_X1 i_1 (.A1(to_int5359[6]), .A2(to_int5359[5]), .A3(to_int5359[4]), 
      .A4(to_int5359[1]), .ZN(n_0));
   NOR2_X1 i_2 (.A1(to_int5359[3]), .A2(to_int5359[2]), .ZN(n_1));
endmodule

module datapath__1_14076(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   NAND2_X1 i_0 (.A1(n_1), .A2(n_0), .ZN(p_0));
   NOR4_X1 i_1 (.A1(to_int5359[6]), .A2(to_int5359[5]), .A3(to_int5359[4]), 
      .A4(to_int5359[2]), .ZN(n_0));
   AOI21_X1 i_2 (.A(to_int5359[3]), .B1(to_int5359[1]), .B2(to_int5359[0]), 
      .ZN(n_1));
endmodule

module datapath__1_14108(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   OR4_X1 i_0 (.A1(to_int5359[4]), .A2(to_int5359[3]), .A3(to_int5359[2]), 
      .A4(to_int5359[5]), .ZN(n_0));
   OR2_X1 i_1 (.A1(n_0), .A2(to_int5359[6]), .ZN(p_0));
endmodule

module datapath__1_14300(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   NAND2_X1 i_0 (.A1(n_1), .A2(n_0), .ZN(p_0));
   NOR3_X1 i_1 (.A1(to_int5359[5]), .A2(to_int5359[4]), .A3(to_int5359[6]), 
      .ZN(n_0));
   OAI21_X1 i_2 (.A(to_int5359[3]), .B1(to_int5359[2]), .B2(to_int5359[1]), 
      .ZN(n_1));
endmodule

module datapath__1_14364(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   OR4_X1 i_0 (.A1(to_int5359[4]), .A2(n_0), .A3(to_int5359[5]), .A4(
      to_int5359[6]), .ZN(p_0));
   AND2_X1 i_1 (.A1(to_int5359[3]), .A2(to_int5359[2]), .ZN(n_0));
endmodule

module datapath__1_14396(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   NAND2_X1 i_0 (.A1(n_1), .A2(n_0), .ZN(p_0));
   NOR3_X1 i_1 (.A1(to_int5359[5]), .A2(to_int5359[4]), .A3(to_int5359[6]), 
      .ZN(n_0));
   OAI211_X1 i_2 (.A(to_int5359[2]), .B(to_int5359[3]), .C1(to_int5359[1]), 
      .C2(to_int5359[0]), .ZN(n_1));
endmodule

module datapath__1_14524(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   NAND2_X1 i_0 (.A1(n_1), .A2(n_0), .ZN(p_0));
   NOR2_X1 i_1 (.A1(to_int5359[6]), .A2(to_int5359[5]), .ZN(n_0));
   OAI21_X1 i_2 (.A(to_int5359[4]), .B1(to_int5359[3]), .B2(n_2), .ZN(n_1));
   OR3_X1 i_3 (.A1(to_int5359[1]), .A2(to_int5359[0]), .A3(to_int5359[2]), 
      .ZN(n_2));
endmodule

module datapath__1_14652(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   NAND2_X1 i_0 (.A1(n_1), .A2(n_0), .ZN(p_0));
   NOR2_X1 i_1 (.A1(to_int5359[6]), .A2(to_int5359[5]), .ZN(n_0));
   OAI21_X1 i_2 (.A(to_int5359[4]), .B1(to_int5359[3]), .B2(n_2), .ZN(n_1));
   INV_X1 i_3 (.A(n_3), .ZN(n_2));
   OAI21_X1 i_4 (.A(to_int5359[2]), .B1(to_int5359[1]), .B2(to_int5359[0]), 
      .ZN(n_3));
endmodule

module datapath__1_14780(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   OR3_X1 i_0 (.A1(to_int5359[5]), .A2(n_0), .A3(to_int5359[6]), .ZN(p_0));
   AND3_X1 i_1 (.A1(to_int5359[3]), .A2(n_1), .A3(to_int5359[4]), .ZN(n_0));
   OR3_X1 i_2 (.A1(to_int5359[1]), .A2(to_int5359[0]), .A3(to_int5359[2]), 
      .ZN(n_1));
endmodule

module datapath__1_14812(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   NAND2_X1 i_0 (.A1(n_1), .A2(n_0), .ZN(p_0));
   NOR2_X1 i_1 (.A1(to_int5359[6]), .A2(to_int5359[5]), .ZN(n_0));
   OAI211_X1 i_2 (.A(to_int5359[3]), .B(to_int5359[4]), .C1(to_int5359[2]), 
      .C2(to_int5359[1]), .ZN(n_1));
endmodule

module datapath__1_14844(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   OAI21_X1 i_0 (.A(n_0), .B1(n_2), .B2(n_1), .ZN(p_0));
   NOR2_X1 i_1 (.A1(to_int5359[6]), .A2(to_int5359[5]), .ZN(n_0));
   NAND2_X1 i_2 (.A1(to_int5359[4]), .A2(to_int5359[3]), .ZN(n_1));
   AOI21_X1 i_3 (.A(to_int5359[2]), .B1(to_int5359[1]), .B2(to_int5359[0]), 
      .ZN(n_2));
endmodule

module datapath__1_14908(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   OR3_X1 i_0 (.A1(to_int5359[5]), .A2(n_0), .A3(to_int5359[6]), .ZN(p_0));
   AND4_X1 i_1 (.A1(to_int5359[2]), .A2(n_1), .A3(to_int5359[3]), .A4(
      to_int5359[4]), .ZN(n_0));
   OR2_X1 i_2 (.A1(to_int5359[1]), .A2(to_int5359[0]), .ZN(n_1));
endmodule

module datapath__1_15420(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   OAI21_X1 i_0 (.A(n_4), .B1(n_3), .B2(n_0), .ZN(p_0));
   AOI21_X1 i_1 (.A(to_int5359[4]), .B1(to_int5359[3]), .B2(n_1), .ZN(n_0));
   INV_X1 i_2 (.A(n_2), .ZN(n_1));
   OAI21_X1 i_3 (.A(to_int5359[2]), .B1(to_int5359[1]), .B2(to_int5359[0]), 
      .ZN(n_2));
   INV_X1 i_4 (.A(to_int5359[5]), .ZN(n_3));
   INV_X1 i_5 (.A(to_int5359[6]), .ZN(n_4));
endmodule

module datapath__1_15452(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   NAND2_X1 i_0 (.A1(n_2), .A2(n_0), .ZN(p_0));
   OAI21_X1 i_1 (.A(to_int5359[5]), .B1(to_int5359[4]), .B2(n_1), .ZN(n_0));
   AND3_X1 i_2 (.A1(to_int5359[2]), .A2(to_int5359[1]), .A3(to_int5359[3]), 
      .ZN(n_1));
   INV_X1 i_3 (.A(to_int5359[6]), .ZN(n_2));
endmodule

module datapath__1_15484(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   OAI21_X1 i_0 (.A(n_3), .B1(n_2), .B2(n_0), .ZN(p_0));
   AOI21_X1 i_1 (.A(to_int5359[4]), .B1(to_int5359[3]), .B2(n_1), .ZN(n_0));
   AND3_X1 i_2 (.A1(to_int5359[1]), .A2(to_int5359[0]), .A3(to_int5359[2]), 
      .ZN(n_1));
   INV_X1 i_3 (.A(to_int5359[5]), .ZN(n_2));
   INV_X1 i_4 (.A(to_int5359[6]), .ZN(n_3));
endmodule

module datapath__1_15516(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0));
   AOI21_X1 i_1 (.A(to_int5359[6]), .B1(to_int5359[5]), .B2(to_int5359[4]), 
      .ZN(n_0));
endmodule

module datapath__1_15676(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   NAND2_X1 i_0 (.A1(n_3), .A2(n_0), .ZN(p_0));
   OAI211_X1 i_1 (.A(to_int5359[4]), .B(to_int5359[5]), .C1(to_int5359[3]), 
      .C2(n_1), .ZN(n_0));
   INV_X1 i_2 (.A(n_2), .ZN(n_1));
   OAI21_X1 i_3 (.A(to_int5359[2]), .B1(to_int5359[1]), .B2(to_int5359[0]), 
      .ZN(n_2));
   INV_X1 i_4 (.A(to_int5359[6]), .ZN(n_3));
endmodule

module datapath__1_15740(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   NAND2_X1 i_0 (.A1(n_2), .A2(n_0), .ZN(p_0));
   OAI211_X1 i_1 (.A(to_int5359[4]), .B(to_int5359[5]), .C1(to_int5359[3]), 
      .C2(n_1), .ZN(n_0));
   AND3_X1 i_2 (.A1(to_int5359[1]), .A2(to_int5359[0]), .A3(to_int5359[2]), 
      .ZN(n_1));
   INV_X1 i_3 (.A(to_int5359[6]), .ZN(n_2));
endmodule

module datapath__1_16117(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   INV_X1 i_0 (.A(to_int5359[6]), .ZN(n_0));
   NOR4_X1 i_1 (.A1(to_int5359[4]), .A2(to_int5359[3]), .A3(to_int5359[5]), 
      .A4(to_int5359[2]), .ZN(n_1));
   NAND2_X1 i_2 (.A1(to_int5359[1]), .A2(to_int5359[0]), .ZN(n_2));
   AOI21_X1 i_3 (.A(n_0), .B1(n_1), .B2(n_2), .ZN(p_0));
endmodule

module datapath__1_16149(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0));
   OAI21_X1 i_1 (.A(to_int5359[6]), .B1(to_int5359[5]), .B2(n_1), .ZN(n_0));
   OR3_X1 i_2 (.A1(to_int5359[3]), .A2(to_int5359[2]), .A3(to_int5359[4]), 
      .ZN(n_1));
endmodule

module datapath__1_16309(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   NOR2_X1 i_0 (.A1(n_2), .A2(n_0), .ZN(p_0));
   AOI211_X1 i_1 (.A(to_int5359[4]), .B(to_int5359[5]), .C1(to_int5359[3]), 
      .C2(n_1), .ZN(n_0));
   OR3_X1 i_2 (.A1(to_int5359[1]), .A2(to_int5359[0]), .A3(to_int5359[2]), 
      .ZN(n_1));
   INV_X1 i_3 (.A(to_int5359[6]), .ZN(n_2));
endmodule

module datapath__1_16437(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   AOI21_X1 i_0 (.A(n_2), .B1(n_1), .B2(n_0), .ZN(p_0));
   NOR2_X1 i_1 (.A1(to_int5359[5]), .A2(to_int5359[4]), .ZN(n_0));
   OAI211_X1 i_2 (.A(to_int5359[2]), .B(to_int5359[3]), .C1(to_int5359[1]), 
      .C2(to_int5359[0]), .ZN(n_1));
   INV_X1 i_3 (.A(to_int5359[6]), .ZN(n_2));
endmodule

module datapath__1_16725(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   NOR2_X1 i_0 (.A1(n_3), .A2(n_0), .ZN(p_0));
   AOI21_X1 i_1 (.A(to_int5359[5]), .B1(to_int5359[4]), .B2(n_1), .ZN(n_0));
   INV_X1 i_2 (.A(n_2), .ZN(n_1));
   AOI21_X1 i_3 (.A(to_int5359[3]), .B1(to_int5359[2]), .B2(to_int5359[1]), 
      .ZN(n_2));
   INV_X1 i_4 (.A(to_int5359[6]), .ZN(n_3));
endmodule

module datapath__1_16757(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0));
   OAI21_X1 i_1 (.A(to_int5359[6]), .B1(to_int5359[5]), .B2(n_1), .ZN(n_0));
   INV_X1 i_2 (.A(n_2), .ZN(n_1));
   OAI21_X1 i_3 (.A(to_int5359[4]), .B1(to_int5359[3]), .B2(n_3), .ZN(n_2));
   AND3_X1 i_4 (.A1(to_int5359[1]), .A2(to_int5359[0]), .A3(to_int5359[2]), 
      .ZN(n_3));
endmodule

module datapath__1_16821(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0));
   OAI21_X1 i_1 (.A(to_int5359[6]), .B1(to_int5359[5]), .B2(n_1), .ZN(n_0));
   AND3_X1 i_2 (.A1(to_int5359[3]), .A2(n_2), .A3(to_int5359[4]), .ZN(n_1));
   OR3_X1 i_3 (.A1(to_int5359[1]), .A2(to_int5359[0]), .A3(to_int5359[2]), 
      .ZN(n_2));
endmodule

module datapath__1_16885(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0));
   OAI21_X1 i_1 (.A(to_int5359[6]), .B1(to_int5359[5]), .B2(n_1), .ZN(n_0));
   NOR2_X1 i_2 (.A1(n_3), .A2(n_2), .ZN(n_1));
   NAND2_X1 i_3 (.A1(to_int5359[4]), .A2(to_int5359[3]), .ZN(n_2));
   AOI21_X1 i_4 (.A(to_int5359[2]), .B1(to_int5359[1]), .B2(to_int5359[0]), 
      .ZN(n_3));
endmodule

module datapath__1_17109(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   AND3_X1 i_0 (.A1(to_int5359[5]), .A2(n_0), .A3(to_int5359[6]), .ZN(p_0));
   OR4_X1 i_1 (.A1(to_int5359[2]), .A2(to_int5359[1]), .A3(to_int5359[3]), 
      .A4(to_int5359[4]), .ZN(n_0));
endmodule

module datapath__1_17397(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0));
   OAI211_X1 i_1 (.A(to_int5359[5]), .B(to_int5359[6]), .C1(to_int5359[4]), 
      .C2(n_1), .ZN(n_0));
   NOR2_X1 i_2 (.A1(n_3), .A2(n_2), .ZN(n_1));
   AOI21_X1 i_3 (.A(to_int5359[2]), .B1(to_int5359[1]), .B2(to_int5359[0]), 
      .ZN(n_2));
   INV_X1 i_4 (.A(to_int5359[3]), .ZN(n_3));
endmodule

module datapath__1_17461(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   AOI21_X1 i_0 (.A(n_0), .B1(n_2), .B2(n_1), .ZN(p_0));
   NAND2_X1 i_1 (.A1(to_int5359[6]), .A2(to_int5359[5]), .ZN(n_0));
   OAI211_X1 i_2 (.A(to_int5359[2]), .B(to_int5359[3]), .C1(to_int5359[1]), 
      .C2(to_int5359[0]), .ZN(n_1));
   INV_X1 i_3 (.A(to_int5359[4]), .ZN(n_2));
endmodule

module datapath__1_17493(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0));
   OAI211_X1 i_1 (.A(to_int5359[5]), .B(to_int5359[6]), .C1(to_int5359[4]), 
      .C2(n_1), .ZN(n_0));
   AND3_X1 i_2 (.A1(to_int5359[2]), .A2(to_int5359[1]), .A3(to_int5359[3]), 
      .ZN(n_1));
endmodule

module datapath__1_17525(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0));
   OAI211_X1 i_1 (.A(to_int5359[5]), .B(to_int5359[6]), .C1(to_int5359[4]), 
      .C2(n_1), .ZN(n_0));
   AND4_X1 i_2 (.A1(to_int5359[1]), .A2(to_int5359[0]), .A3(to_int5359[2]), 
      .A4(to_int5359[3]), .ZN(n_1));
endmodule

module datapath__1_17781(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   AND4_X1 i_0 (.A1(to_int5359[4]), .A2(n_0), .A3(to_int5359[5]), .A4(
      to_int5359[6]), .ZN(p_0));
   OR2_X1 i_1 (.A1(to_int5359[3]), .A2(n_1), .ZN(n_0));
   AND3_X1 i_2 (.A1(to_int5359[1]), .A2(to_int5359[0]), .A3(to_int5359[2]), 
      .ZN(n_1));
endmodule

module datapath__1_17877(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   NOR2_X1 i_0 (.A1(n_1), .A2(n_0), .ZN(p_0));
   OAI211_X1 i_1 (.A(to_int5359[5]), .B(to_int5359[4]), .C1(to_int5359[2]), 
      .C2(to_int5359[1]), .ZN(n_0));
   NAND2_X1 i_2 (.A1(to_int5359[6]), .A2(to_int5359[3]), .ZN(n_1));
endmodule

module datapath__1_17909(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   NOR2_X1 i_0 (.A1(n_1), .A2(n_0), .ZN(p_0));
   NAND4_X1 i_1 (.A1(to_int5359[5]), .A2(to_int5359[4]), .A3(to_int5359[6]), 
      .A4(to_int5359[3]), .ZN(n_0));
   AOI21_X1 i_2 (.A(to_int5359[2]), .B1(to_int5359[1]), .B2(to_int5359[0]), 
      .ZN(n_1));
endmodule

module datapath__1_17973(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   NOR2_X1 i_0 (.A1(n_1), .A2(n_0), .ZN(p_0));
   OAI21_X1 i_1 (.A(to_int5359[3]), .B1(to_int5359[1]), .B2(to_int5359[0]), 
      .ZN(n_0));
   NAND4_X1 i_2 (.A1(to_int5359[6]), .A2(to_int5359[5]), .A3(to_int5359[4]), 
      .A4(to_int5359[2]), .ZN(n_1));
endmodule

module datapath__1_13530(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NAND2_X1 i_0 (.A1(n_3), .A2(n_0), .ZN(p_0));
   NOR4_X1 i_1 (.A1(to_int6126[5]), .A2(to_int6126[4]), .A3(to_int6126[3]), 
      .A4(n_1), .ZN(n_0));
   INV_X1 i_2 (.A(n_2), .ZN(n_1));
   OAI21_X1 i_3 (.A(to_int6126[2]), .B1(to_int6126[1]), .B2(to_int6126[0]), 
      .ZN(n_2));
   INV_X1 i_4 (.A(to_int6126[6]), .ZN(n_3));
endmodule

module datapath__1_13546(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NAND2_X1 i_0 (.A1(n_2), .A2(n_0), .ZN(p_0));
   AOI211_X1 i_1 (.A(to_int6126[4]), .B(to_int6126[5]), .C1(to_int6126[3]), 
      .C2(n_1), .ZN(n_0));
   OR3_X1 i_2 (.A1(to_int6126[2]), .A2(to_int6126[1]), .A3(to_int6126[0]), 
      .ZN(n_1));
   INV_X1 i_3 (.A(to_int6126[6]), .ZN(n_2));
endmodule

module datapath__1_13554(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NAND2_X1 i_0 (.A1(n_4), .A2(n_0), .ZN(p_0));
   AOI211_X1 i_1 (.A(to_int6126[4]), .B(to_int6126[5]), .C1(to_int6126[3]), 
      .C2(n_1), .ZN(n_0));
   NAND2_X1 i_2 (.A1(n_2), .A2(n_3), .ZN(n_1));
   NAND2_X1 i_3 (.A1(to_int6126[1]), .A2(to_int6126[0]), .ZN(n_2));
   INV_X1 i_4 (.A(to_int6126[2]), .ZN(n_3));
   INV_X1 i_5 (.A(to_int6126[6]), .ZN(n_4));
endmodule

module datapath__1_13630(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NAND2_X1 i_0 (.A1(n_3), .A2(n_0), .ZN(p_0));
   AOI21_X1 i_1 (.A(to_int6126[5]), .B1(to_int6126[4]), .B2(n_1), .ZN(n_0));
   INV_X1 i_2 (.A(n_2), .ZN(n_1));
   NAND3_X1 i_3 (.A1(to_int6126[3]), .A2(to_int6126[2]), .A3(to_int6126[1]), 
      .ZN(n_2));
   INV_X1 i_4 (.A(to_int6126[6]), .ZN(n_3));
endmodule

module full_adder__3_51(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XNOR2_X1 i_0_0 (.A(b), .B(a), .ZN(f));
   OR2_X1 i_0_1 (.A1(b), .A2(a), .ZN(cout));
endmodule

module full_adder__3_55(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(cin), .Z(f));
endmodule

module int_adder__parameterized1(a, b, cin, enbl, c, cout);
   input [6:0]a;
   input [6:0]b;
   input cin;
   input enbl;
   output [6:0]c;
   output cout;

   full_adder__3_51 full_adder_0_5_full_adder_0_i (.a(a[5]), .b(b[5]), .cin(), 
      .f(c[5]), .cout(n_0));
   full_adder__3_55 full_adder_0_6_full_adder_0_i (.a(a[6]), .b(b[6]), .cin(n_0), 
      .f(c[6]), .cout());
endmodule

module datapath__1_13570(to_int6126, p_0);
   input [7:0]to_int6126;
   output p_0;

   NAND2_X1 i_0 (.A1(n_3), .A2(n_0), .ZN(p_0));
   NOR3_X1 i_1 (.A1(to_int6126[5]), .A2(to_int6126[4]), .A3(n_1), .ZN(n_0));
   INV_X1 i_2 (.A(n_2), .ZN(n_1));
   NAND4_X1 i_3 (.A1(to_int6126[3]), .A2(to_int6126[2]), .A3(to_int6126[1]), 
      .A4(to_int6126[0]), .ZN(n_2));
   INV_X1 i_4 (.A(to_int6126[6]), .ZN(n_3));
endmodule

module datapath__1_14204(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   NAND2_X1 i_0 (.A1(n_1), .A2(n_0), .ZN(p_0));
   NOR4_X1 i_1 (.A1(to_int5359[5]), .A2(to_int5359[4]), .A3(to_int5359[6]), 
      .A4(to_int5359[3]), .ZN(n_0));
   NAND3_X1 i_2 (.A1(to_int5359[1]), .A2(to_int5359[0]), .A3(to_int5359[2]), 
      .ZN(n_1));
endmodule

module datapath__1_14236(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   OR4_X1 i_0 (.A1(to_int5359[4]), .A2(to_int5359[3]), .A3(to_int5359[5]), 
      .A4(to_int5359[6]), .ZN(p_0));
endmodule

module datapath__1_14588(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   NAND2_X1 i_0 (.A1(n_1), .A2(n_0), .ZN(p_0));
   NOR2_X1 i_1 (.A1(to_int5359[6]), .A2(to_int5359[5]), .ZN(n_0));
   OAI21_X1 i_2 (.A(to_int5359[4]), .B1(to_int5359[3]), .B2(n_2), .ZN(n_1));
   INV_X1 i_3 (.A(n_3), .ZN(n_2));
   AOI21_X1 i_4 (.A(to_int5359[2]), .B1(to_int5359[1]), .B2(to_int5359[0]), 
      .ZN(n_3));
endmodule

module datapath__1_14620(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   NAND2_X1 i_0 (.A1(n_1), .A2(n_0), .ZN(p_0));
   NOR2_X1 i_1 (.A1(to_int5359[6]), .A2(to_int5359[5]), .ZN(n_0));
   OAI21_X1 i_2 (.A(to_int5359[4]), .B1(to_int5359[3]), .B2(to_int5359[2]), 
      .ZN(n_1));
endmodule

module datapath__1_14684(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   OAI21_X1 i_0 (.A(n_0), .B1(n_2), .B2(n_1), .ZN(p_0));
   NOR2_X1 i_1 (.A1(to_int5359[6]), .A2(to_int5359[5]), .ZN(n_0));
   AOI21_X1 i_2 (.A(to_int5359[3]), .B1(to_int5359[2]), .B2(to_int5359[1]), 
      .ZN(n_1));
   INV_X1 i_3 (.A(to_int5359[4]), .ZN(n_2));
endmodule

module datapath__1_14716(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   NAND2_X1 i_0 (.A1(n_1), .A2(n_0), .ZN(p_0));
   NOR2_X1 i_1 (.A1(to_int5359[6]), .A2(to_int5359[5]), .ZN(n_0));
   OAI21_X1 i_2 (.A(to_int5359[4]), .B1(to_int5359[3]), .B2(n_2), .ZN(n_1));
   AND3_X1 i_3 (.A1(to_int5359[1]), .A2(to_int5359[0]), .A3(to_int5359[2]), 
      .ZN(n_2));
endmodule

module datapath__1_14972(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   OAI21_X1 i_0 (.A(n_0), .B1(n_2), .B2(n_1), .ZN(p_0));
   NOR2_X1 i_1 (.A1(to_int5359[6]), .A2(to_int5359[5]), .ZN(n_0));
   NAND4_X1 i_2 (.A1(to_int5359[2]), .A2(to_int5359[1]), .A3(to_int5359[0]), 
      .A4(to_int5359[3]), .ZN(n_1));
   INV_X1 i_3 (.A(to_int5359[4]), .ZN(n_2));
endmodule

module datapath__1_16053(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   INV_X1 i_0 (.A(to_int5359[6]), .ZN(n_0));
   NOR4_X1 i_1 (.A1(to_int5359[1]), .A2(to_int5359[0]), .A3(to_int5359[2]), 
      .A4(to_int5359[3]), .ZN(n_1));
   NOR2_X1 i_2 (.A1(to_int5359[5]), .A2(to_int5359[4]), .ZN(n_2));
   AOI21_X1 i_3 (.A(n_0), .B1(n_1), .B2(n_2), .ZN(p_0));
endmodule

module datapath__1_16469(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   AND3_X1 i_0 (.A1(to_int5359[2]), .A2(to_int5359[1]), .A3(to_int5359[3]), 
      .ZN(n_0));
   OR3_X1 i_1 (.A1(n_0), .A2(to_int5359[4]), .A3(to_int5359[5]), .ZN(n_1));
   AND2_X1 i_2 (.A1(n_1), .A2(to_int5359[6]), .ZN(p_0));
endmodule

module datapath__1_16501(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   AND4_X1 i_0 (.A1(to_int5359[1]), .A2(to_int5359[0]), .A3(to_int5359[2]), 
      .A4(to_int5359[3]), .ZN(n_0));
   OR3_X1 i_1 (.A1(n_0), .A2(to_int5359[4]), .A3(to_int5359[5]), .ZN(n_1));
   AND2_X1 i_2 (.A1(n_1), .A2(to_int5359[6]), .ZN(p_0));
endmodule

module datapath__1_16565(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0));
   OAI21_X1 i_1 (.A(to_int5359[6]), .B1(to_int5359[5]), .B2(n_1), .ZN(n_0));
   INV_X1 i_2 (.A(n_2), .ZN(n_1));
   OAI21_X1 i_3 (.A(to_int5359[4]), .B1(to_int5359[3]), .B2(n_3), .ZN(n_2));
   OR3_X1 i_4 (.A1(to_int5359[1]), .A2(to_int5359[0]), .A3(to_int5359[2]), 
      .ZN(n_3));
endmodule

module datapath__1_16629(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0));
   OAI21_X1 i_1 (.A(to_int5359[6]), .B1(to_int5359[5]), .B2(n_1), .ZN(n_0));
   INV_X1 i_2 (.A(n_2), .ZN(n_1));
   OAI21_X1 i_3 (.A(to_int5359[4]), .B1(to_int5359[3]), .B2(n_3), .ZN(n_2));
   INV_X1 i_4 (.A(n_4), .ZN(n_3));
   AOI21_X1 i_5 (.A(to_int5359[2]), .B1(to_int5359[1]), .B2(to_int5359[0]), 
      .ZN(n_4));
endmodule

module datapath__1_16693(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0));
   OAI21_X1 i_1 (.A(to_int5359[6]), .B1(to_int5359[5]), .B2(n_1), .ZN(n_0));
   INV_X1 i_2 (.A(n_2), .ZN(n_1));
   OAI21_X1 i_3 (.A(to_int5359[4]), .B1(to_int5359[3]), .B2(n_3), .ZN(n_2));
   INV_X1 i_4 (.A(n_4), .ZN(n_3));
   OAI21_X1 i_5 (.A(to_int5359[2]), .B1(to_int5359[1]), .B2(to_int5359[0]), 
      .ZN(n_4));
endmodule

module datapath__1_17301(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0));
   OAI211_X1 i_1 (.A(to_int5359[5]), .B(to_int5359[6]), .C1(to_int5359[4]), 
      .C2(to_int5359[3]), .ZN(n_0));
endmodule

module datapath__1_17045(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   AND2_X1 i_0 (.A1(to_int5359[6]), .A2(to_int5359[5]), .ZN(p_0));
endmodule

module datapath__1_14748(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   INV_X1 i_0 (.A(n_0), .ZN(p_0));
   AOI211_X1 i_1 (.A(to_int5359[5]), .B(to_int5359[6]), .C1(to_int5359[4]), 
      .C2(to_int5359[3]), .ZN(n_0));
endmodule

module datapath__1_14940(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   OR3_X1 i_0 (.A1(to_int5359[5]), .A2(n_0), .A3(to_int5359[6]), .ZN(p_0));
   AND4_X1 i_1 (.A1(to_int5359[2]), .A2(to_int5359[1]), .A3(to_int5359[3]), 
      .A4(to_int5359[4]), .ZN(n_0));
endmodule

module datapath__1_14460(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   OR4_X1 i_0 (.A1(to_int5359[4]), .A2(n_0), .A3(to_int5359[5]), .A4(
      to_int5359[6]), .ZN(p_0));
   AND4_X1 i_1 (.A1(to_int5359[1]), .A2(to_int5359[0]), .A3(to_int5359[2]), 
      .A4(to_int5359[3]), .ZN(n_0));
endmodule

module datapath__1_14428(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   OR4_X1 i_0 (.A1(to_int5359[4]), .A2(n_0), .A3(to_int5359[5]), .A4(
      to_int5359[6]), .ZN(p_0));
   AND3_X1 i_1 (.A1(to_int5359[2]), .A2(to_int5359[1]), .A3(to_int5359[3]), 
      .ZN(n_0));
endmodule

module datapath__1_14332(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   OAI21_X1 i_0 (.A(n_0), .B1(n_2), .B2(n_1), .ZN(p_0));
   NOR3_X1 i_1 (.A1(to_int5359[5]), .A2(to_int5359[4]), .A3(to_int5359[6]), 
      .ZN(n_0));
   AOI21_X1 i_2 (.A(to_int5359[2]), .B1(to_int5359[1]), .B2(to_int5359[0]), 
      .ZN(n_1));
   INV_X1 i_3 (.A(to_int5359[3]), .ZN(n_2));
endmodule

module datapath__1_14268(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   OAI21_X1 i_0 (.A(n_0), .B1(n_2), .B2(n_1), .ZN(p_0));
   NOR3_X1 i_1 (.A1(to_int5359[5]), .A2(to_int5359[4]), .A3(to_int5359[6]), 
      .ZN(n_0));
   NOR3_X1 i_2 (.A1(to_int5359[1]), .A2(to_int5359[0]), .A3(to_int5359[2]), 
      .ZN(n_1));
   INV_X1 i_3 (.A(to_int5359[3]), .ZN(n_2));
endmodule

module datapath__1_14140(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   NAND2_X1 i_0 (.A1(n_1), .A2(n_0), .ZN(p_0));
   NOR4_X1 i_1 (.A1(to_int5359[5]), .A2(to_int5359[4]), .A3(to_int5359[6]), 
      .A4(to_int5359[3]), .ZN(n_0));
   OAI21_X1 i_2 (.A(to_int5359[2]), .B1(to_int5359[1]), .B2(to_int5359[0]), 
      .ZN(n_1));
endmodule

module datapath__1_14876(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   OR3_X1 i_0 (.A1(to_int5359[5]), .A2(n_0), .A3(to_int5359[6]), .ZN(p_0));
   AND3_X1 i_1 (.A1(to_int5359[3]), .A2(to_int5359[2]), .A3(to_int5359[4]), 
      .ZN(n_0));
endmodule

module datapath__1_14492(to_int5359, p_0);
   input [7:0]to_int5359;
   output p_0;

   OR3_X1 i_0 (.A1(to_int5359[5]), .A2(to_int5359[4]), .A3(to_int5359[6]), 
      .ZN(p_0));
endmodule

module full_adder__3_79(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   INV_X1 i_3 (.A(a), .ZN(f));
endmodule

module full_adder(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
endmodule

module int_adder__parameterized0(a, b, cin, enbl, c, cout);
   input [6:0]a;
   input [5:0]b;
   input cin;
   input enbl;
   output [6:0]c;
   output cout;

   full_adder__3_79 full_adder_0_5_full_adder_0_i (.a(a[5]), .b(), .cin(), 
      .f(c[5]), .cout());
   full_adder full_adder_0_6_full_adder_0_i (.a(a[6]), .b(), .cin(a[5]), 
      .f(c[6]), .cout());
endmodule

module decompressor(in_data, rst, enbl_in, clk, state_wait, out_ready, out_data, 
      error_success, buf_test);
   input [31:0]in_data;
   input rst;
   input enbl_in;
   input clk;
   input state_wait;
   output out_ready;
   output [31:0]out_data;
   output error_success;
   output [127:0]buf_test;

   wire [6:0]\out_bs[6] ;
   wire [6:0]\out_as[6] ;
   wire n_1_737_0;
   wire n_1_737_1;
   wire n_1_737_2;
   wire n_1_737_3;
   wire n_1_737_4;
   wire n_1_737_5;
   wire n_1_737_6;
   wire n_1_737_7;
   wire n_1_737_8;
   wire n_1_737_9;
   wire n_1_737_10;
   wire n_1_737_11;
   wire n_1_737_12;
   wire n_1_737_13;
   wire n_1_737_14;
   wire n_1_737_15;
   wire n_1_737_16;
   wire n_1_737_17;
   wire n_1_737_18;
   wire n_1_737_19;
   wire n_1_737_20;
   wire n_1_737_21;
   wire n_1_737_22;
   wire n_1_737_23;
   wire n_1_737_24;
   wire n_1_737_25;
   wire n_1_737_26;
   wire n_1_737_27;
   wire n_1_737_28;
   wire n_1_737_29;
   wire n_1_737_30;
   wire n_1_737_31;
   wire n_1_737_32;
   wire n_1_737_33;
   wire n_1_737_34;
   wire n_1_737_35;
   wire n_1_737_36;
   wire n_1_737_37;
   wire n_1_737_38;
   wire n_1_737_39;
   wire n_1_737_40;
   wire n_1_737_41;
   wire n_1_737_42;
   wire n_1_737_43;
   wire n_1_737_44;
   wire n_1_737_45;
   wire n_1_737_46;
   wire n_1_737_47;
   wire n_1_737_48;
   wire n_1_737_49;
   wire n_1_737_50;
   wire n_1_737_51;
   wire n_1_737_52;
   wire n_1_737_53;
   wire n_1_737_54;
   wire n_1_737_55;
   wire n_1_737_56;
   wire n_1_737_57;
   wire n_1_737_58;
   wire n_1_737_59;
   wire n_1_737_60;
   wire n_1_737_61;
   wire n_1_737_62;
   wire n_1_737_63;
   wire n_1_737_64;
   wire n_1_737_65;
   wire n_1_737_66;
   wire n_1_737_67;
   wire n_1_737_68;
   wire n_1_737_69;
   wire n_1_737_70;
   wire n_1_737_71;
   wire n_1_737_72;
   wire n_1_737_73;
   wire n_1_737_74;
   wire n_1_737_75;
   wire n_1_737_76;
   wire n_1_737_77;
   wire n_1_737_78;
   wire n_1_737_79;
   wire n_1_737_80;
   wire n_1_737_81;
   wire n_1_737_82;
   wire n_1_737_83;
   wire n_1_737_84;
   wire n_1_737_85;
   wire n_1_737_86;
   wire n_1_737_87;
   wire n_1_737_88;
   wire n_1_737_89;
   wire n_1_737_90;
   wire n_1_737_91;
   wire n_1_737_92;
   wire n_1_737_93;
   wire n_1_737_94;
   wire n_1_737_95;
   wire n_1_737_96;
   wire n_1_737_97;
   wire n_1_737_98;
   wire n_1_737_99;
   wire n_1_737_100;
   wire n_1_737_101;
   wire n_1_737_102;
   wire n_1_737_103;
   wire n_1_737_104;
   wire n_1_737_105;
   wire n_1_737_106;
   wire n_1_737_107;
   wire n_1_737_108;
   wire n_1_737_109;
   wire n_1_737_110;
   wire n_1_737_111;
   wire n_1_737_112;
   wire n_1_737_113;
   wire n_1_737_114;
   wire n_1_737_115;
   wire n_1_737_116;
   wire n_1_737_117;
   wire n_1_737_118;
   wire n_1_737_119;
   wire n_1_737_120;
   wire n_1_737_121;
   wire n_1_737_122;
   wire n_1_737_123;
   wire n_1_737_124;
   wire n_1_737_125;
   wire n_1_737_126;
   wire n_1_737_127;
   wire n_1_737_128;
   wire n_1_737_129;
   wire n_1_737_130;
   wire n_1_737_131;
   wire n_1_737_132;
   wire n_1_737_133;
   wire n_1_737_134;
   wire n_1_737_135;
   wire n_1_737_136;
   wire n_1_737_137;
   wire n_1_737_138;
   wire n_1_737_139;
   wire n_1_737_140;
   wire n_1_737_141;
   wire n_1_737_142;
   wire n_1_737_143;
   wire n_1_737_144;
   wire n_1_737_145;
   wire n_1_737_146;
   wire n_1_737_147;
   wire n_1_737_148;
   wire n_1_737_149;
   wire n_1_737_150;
   wire n_1_737_151;
   wire n_1_737_152;
   wire n_1_737_153;
   wire n_1_737_154;
   wire n_1_737_155;
   wire n_1_737_156;
   wire n_1_737_157;
   wire n_1_737_158;
   wire n_1_737_159;
   wire n_1_737_160;
   wire n_1_737_161;
   wire n_1_737_162;
   wire n_1_737_163;
   wire n_1_737_164;
   wire n_1_737_165;
   wire n_1_737_166;
   wire n_1_737_167;
   wire n_1_737_168;
   wire n_1_737_169;
   wire n_1_737_170;
   wire n_1_737_171;
   wire n_1_737_172;
   wire n_1_737_173;
   wire n_1_737_174;
   wire n_1_737_175;
   wire n_1_737_176;
   wire n_1_737_177;
   wire n_1_737_178;
   wire n_1_737_179;
   wire n_1_737_180;
   wire n_1_737_181;
   wire n_1_737_182;
   wire n_1_737_183;
   wire n_1_737_184;
   wire n_1_737_185;
   wire n_1_737_186;
   wire n_1_737_187;
   wire n_1_737_188;
   wire n_1_737_189;
   wire n_1_737_190;
   wire n_1_737_191;
   wire n_1_737_192;
   wire n_1_737_193;
   wire n_1_737_194;
   wire n_1_737_195;
   wire n_1_737_196;
   wire n_1_737_197;
   wire n_1_737_198;
   wire n_1_737_199;
   wire n_1_737_200;
   wire n_1_737_201;
   wire n_1_737_202;
   wire n_1_737_203;
   wire n_1_737_204;
   wire n_1_737_205;
   wire n_1_737_206;
   wire n_1_737_207;
   wire n_1_737_208;
   wire n_1_737_209;
   wire n_1_737_210;
   wire n_1_737_211;
   wire n_1_737_212;
   wire n_1_737_213;
   wire n_1_737_214;
   wire n_1_737_215;
   wire n_1_737_216;
   wire n_1_737_217;
   wire n_1_737_218;
   wire n_1_737_219;
   wire n_1_737_220;
   wire n_1_737_221;
   wire n_1_737_222;
   wire n_1_737_223;
   wire n_1_737_224;
   wire n_1_737_225;
   wire n_1_737_226;
   wire n_1_737_227;
   wire n_1_737_228;
   wire n_1_737_229;
   wire n_1_737_230;
   wire n_1_737_231;
   wire n_1_737_232;
   wire n_1_737_233;
   wire n_1_737_234;
   wire n_1_737_235;
   wire n_1_737_236;
   wire n_1_737_237;
   wire n_1_737_238;
   wire n_1_737_239;
   wire n_1_737_240;
   wire n_1_737_241;
   wire n_1_737_242;
   wire n_1_737_243;
   wire n_1_737_244;
   wire n_1_737_245;
   wire n_1_737_246;
   wire n_1_737_247;
   wire n_1_737_248;
   wire n_1_737_249;
   wire n_1_737_250;
   wire n_1_737_251;
   wire n_1_737_252;
   wire n_1_737_253;
   wire n_1_737_254;
   wire n_1_737_255;
   wire n_1_737_256;
   wire n_1_737_257;
   wire n_1_737_258;
   wire n_1_737_259;
   wire n_1_737_260;
   wire n_1_737_261;
   wire n_1_737_262;
   wire n_1_737_263;
   wire n_1_737_264;
   wire n_1_737_265;
   wire n_1_737_266;
   wire n_1_737_267;
   wire n_1_737_268;
   wire n_1_737_269;
   wire n_1_737_270;
   wire n_1_737_271;
   wire n_1_737_272;
   wire n_1_737_273;
   wire n_1_737_274;
   wire n_1_737_275;
   wire n_1_737_276;
   wire n_1_737_277;
   wire n_1_737_278;
   wire n_1_737_279;
   wire n_1_737_280;
   wire n_1_737_281;
   wire n_1_737_282;
   wire n_1_737_283;
   wire n_1_737_284;
   wire n_1_737_285;
   wire n_1_737_286;
   wire n_1_737_287;
   wire n_1_737_288;
   wire n_1_737_289;
   wire n_1_737_290;
   wire n_1_737_291;
   wire n_1_737_292;
   wire n_1_737_293;
   wire n_1_737_294;
   wire n_1_737_295;
   wire n_1_737_296;
   wire n_1_737_297;
   wire n_1_737_298;
   wire n_1_737_299;
   wire n_1_737_300;
   wire n_1_737_301;
   wire n_1_737_302;
   wire n_1_737_303;
   wire n_1_737_304;
   wire n_1_737_305;
   wire n_1_737_306;
   wire n_1_737_307;
   wire n_1_737_308;
   wire n_1_737_309;
   wire n_1_737_310;
   wire n_1_737_311;
   wire n_1_737_312;
   wire n_1_737_313;
   wire n_1_737_314;
   wire n_1_737_315;
   wire n_1_737_316;
   wire n_1_737_317;
   wire n_1_737_318;
   wire n_1_737_319;
   wire n_1_737_320;
   wire n_1_737_321;
   wire n_1_737_322;
   wire n_1_737_323;
   wire n_1_737_324;
   wire n_1_737_325;
   wire n_1_737_326;
   wire n_1_737_327;
   wire n_1_737_328;
   wire n_1_737_329;
   wire n_1_737_330;
   wire n_1_737_331;
   wire n_1_737_332;
   wire n_1_737_333;
   wire n_1_737_334;
   wire n_1_737_335;
   wire n_1_737_336;
   wire n_1_737_337;
   wire n_1_737_338;
   wire n_1_737_339;
   wire n_1_737_340;
   wire n_1_737_341;
   wire n_1_737_342;
   wire n_1_737_343;
   wire n_1_737_344;
   wire n_1_737_345;
   wire n_1_737_346;
   wire n_1_737_347;
   wire n_1_737_348;
   wire n_1_737_349;
   wire n_1_737_350;
   wire n_1_737_351;
   wire n_1_737_352;
   wire n_1_737_353;
   wire n_1_737_354;
   wire n_1_737_355;
   wire n_1_737_356;
   wire n_1_737_357;
   wire n_1_737_358;
   wire n_1_737_359;
   wire n_1_737_360;
   wire n_1_737_361;
   wire n_1_737_362;
   wire n_1_737_363;
   wire n_1_737_364;
   wire n_1_737_365;
   wire n_1_737_366;
   wire n_1_737_367;
   wire n_1_737_368;
   wire n_1_737_369;
   wire n_1_737_370;
   wire n_1_737_371;
   wire n_1_737_372;
   wire n_1_737_373;
   wire n_1_737_374;
   wire n_1_737_375;
   wire n_1_737_376;
   wire n_1_737_377;
   wire n_1_737_378;
   wire n_1_737_379;
   wire n_1_737_380;
   wire n_1_737_381;
   wire n_1_737_382;
   wire n_1_737_383;
   wire n_1_737_384;
   wire n_1_737_385;
   wire n_1_737_386;
   wire n_1_737_387;
   wire n_1_737_388;
   wire n_1_737_389;
   wire n_1_737_390;
   wire n_1_737_391;
   wire n_1_737_392;
   wire n_1_737_393;
   wire n_1_737_394;
   wire n_1_737_395;
   wire n_1_737_396;
   wire n_1_737_397;
   wire n_1_737_398;
   wire n_1_737_399;
   wire n_1_737_400;
   wire n_1_737_401;
   wire n_1_737_402;
   wire n_1_737_403;
   wire n_1_737_404;
   wire n_1_737_405;
   wire n_1_737_406;
   wire n_1_737_407;
   wire n_1_737_408;
   wire n_1_737_409;
   wire n_1_737_410;
   wire n_1_737_411;
   wire n_1_737_412;
   wire n_1_737_413;
   wire n_1_737_414;
   wire n_1_737_415;
   wire n_1_737_416;
   wire n_1_737_417;
   wire n_1_737_418;
   wire n_1_737_419;
   wire n_1_737_420;
   wire n_1_737_421;
   wire n_1_737_422;
   wire n_1_737_423;
   wire n_1_737_424;
   wire n_1_737_425;
   wire n_1_737_426;
   wire n_1_737_427;
   wire n_1_737_428;
   wire n_1_737_429;
   wire n_1_737_430;
   wire n_1_737_431;
   wire n_1_737_432;
   wire n_1_737_433;
   wire n_1_737_434;
   wire n_1_737_435;
   wire n_1_737_436;
   wire n_1_737_437;
   wire n_1_737_438;
   wire n_1_737_439;
   wire n_1_737_440;
   wire n_1_737_441;
   wire n_1_737_442;
   wire n_1_737_443;
   wire n_1_737_444;
   wire n_1_737_445;
   wire n_1_737_446;
   wire n_1_737_447;
   wire n_1_737_448;
   wire n_1_737_449;
   wire n_1_737_450;
   wire n_1_737_451;
   wire n_1_737_452;
   wire n_1_737_453;
   wire n_1_737_454;
   wire n_1_737_455;
   wire n_1_737_456;
   wire n_1_737_457;
   wire n_1_737_458;
   wire n_1_737_459;
   wire n_1_737_460;
   wire n_1_737_461;
   wire n_1_737_462;
   wire n_1_737_463;
   wire n_1_737_464;
   wire n_1_737_465;
   wire n_1_737_466;
   wire n_1_737_467;
   wire n_1_737_468;
   wire n_1_737_469;
   wire n_1_737_470;
   wire n_1_737_471;
   wire n_1_737_472;
   wire n_1_737_473;
   wire n_1_737_474;
   wire n_1_737_475;
   wire n_1_737_476;
   wire n_1_737_477;
   wire n_1_737_478;
   wire n_1_737_479;
   wire n_1_737_480;
   wire n_1_737_481;
   wire n_1_737_482;
   wire n_1_737_483;
   wire n_1_737_484;
   wire n_1_737_485;
   wire n_1_737_486;
   wire n_1_737_487;
   wire n_1_737_488;
   wire n_1_737_489;
   wire n_1_737_490;
   wire n_1_737_491;
   wire n_1_737_492;
   wire n_1_737_493;
   wire n_1_737_494;
   wire n_1_737_495;
   wire n_1_737_496;
   wire n_1_737_497;
   wire n_1_737_498;
   wire n_1_737_499;
   wire n_1_737_500;
   wire n_1_737_501;
   wire n_1_737_502;
   wire n_1_737_503;
   wire n_1_737_504;
   wire n_1_737_505;
   wire n_1_737_506;
   wire n_1_737_507;
   wire n_1_737_508;
   wire n_1_737_509;
   wire n_1_737_510;
   wire n_1_737_511;
   wire n_1_737_512;
   wire n_1_737_513;
   wire n_1_737_514;
   wire n_1_737_515;
   wire n_1_737_516;
   wire n_1_737_517;
   wire n_1_737_518;
   wire n_1_737_519;
   wire n_1_737_520;
   wire n_1_737_521;
   wire n_1_737_522;
   wire n_1_737_523;
   wire n_1_737_524;
   wire n_1_737_525;
   wire n_1_737_526;
   wire n_1_737_527;
   wire n_1_737_528;
   wire n_1_737_529;
   wire n_1_737_530;
   wire n_1_737_531;
   wire n_1_737_532;
   wire n_1_737_533;
   wire n_1_737_534;
   wire n_1_737_535;
   wire n_1_737_536;
   wire n_1_737_537;
   wire n_1_737_538;
   wire n_1_737_539;
   wire n_1_737_540;
   wire n_1_737_541;
   wire n_1_737_542;
   wire n_1_737_543;
   wire n_1_737_544;
   wire n_1_737_545;
   wire n_1_737_546;
   wire n_1_737_547;
   wire n_1_737_548;
   wire n_1_737_549;
   wire n_1_737_550;
   wire n_1_737_551;
   wire n_1_737_552;
   wire n_1_737_553;
   wire n_1_737_554;
   wire n_1_737_555;
   wire n_1_737_556;
   wire n_1_737_557;
   wire n_1_737_558;
   wire n_1_737_559;
   wire n_1_737_560;
   wire n_1_737_561;
   wire n_1_737_562;
   wire n_1_737_563;
   wire n_1_737_564;
   wire n_1_737_565;
   wire n_1_737_566;
   wire n_1_737_567;
   wire n_1_737_568;
   wire n_1_737_569;
   wire n_1_737_570;
   wire n_1_737_571;
   wire n_1_737_572;
   wire n_1_737_573;
   wire n_1_737_574;
   wire n_1_737_575;
   wire n_1_737_576;
   wire n_1_737_577;
   wire n_1_737_578;
   wire n_1_737_579;
   wire n_1_737_580;
   wire n_1_737_581;
   wire n_1_737_582;
   wire n_1_737_583;
   wire n_1_737_584;
   wire n_1_737_585;
   wire n_1_737_586;
   wire n_1_737_587;
   wire n_1_737_588;
   wire n_1_737_589;
   wire n_1_737_590;
   wire n_1_737_591;
   wire n_1_737_592;
   wire n_1_737_593;
   wire n_1_737_594;
   wire n_1_737_595;
   wire n_1_737_596;
   wire n_1_737_597;
   wire n_1_737_598;
   wire n_1_737_599;
   wire n_1_737_600;
   wire n_1_737_601;
   wire n_1_737_602;
   wire n_1_737_603;
   wire n_1_737_604;
   wire n_1_737_605;
   wire n_1_737_606;
   wire n_1_737_607;
   wire n_1_737_608;
   wire n_1_737_609;
   wire n_1_737_610;
   wire n_1_737_611;
   wire n_1_737_612;
   wire n_1_737_613;
   wire n_1_737_614;
   wire n_1_737_615;
   wire n_1_737_616;
   wire n_1_737_617;
   wire n_1_737_618;
   wire n_1_737_619;
   wire n_1_737_620;
   wire n_1_737_621;
   wire n_1_737_622;
   wire n_1_737_623;
   wire n_1_737_624;
   wire n_1_737_625;
   wire n_1_737_626;
   wire n_1_737_627;
   wire n_1_737_628;
   wire n_1_737_629;
   wire n_1_737_630;
   wire n_1_737_631;
   wire n_1_737_632;
   wire n_1_737_633;
   wire n_1_737_634;
   wire n_1_737_635;
   wire n_1_737_636;
   wire n_1_737_637;
   wire n_1_737_638;
   wire n_1_737_639;
   wire n_1_737_640;
   wire n_1_737_641;
   wire n_1_737_642;
   wire n_1_737_643;
   wire n_1_737_644;
   wire n_1_737_645;
   wire n_1_737_646;
   wire n_1_737_647;
   wire n_1_737_648;
   wire n_1_737_649;
   wire n_1_737_650;
   wire n_1_737_651;
   wire n_1_737_652;
   wire n_1_737_653;
   wire n_1_737_654;
   wire n_1_737_655;
   wire n_1_737_656;
   wire n_1_737_657;
   wire n_1_737_658;
   wire n_1_737_659;
   wire n_1_737_660;
   wire n_1_737_661;
   wire n_1_737_662;
   wire n_1_737_663;
   wire n_1_737_664;
   wire n_1_737_665;
   wire n_1_737_666;
   wire n_1_737_667;
   wire n_1_737_668;
   wire n_1_737_669;
   wire n_1_737_670;
   wire n_1_737_671;
   wire n_1_737_672;
   wire n_1_737_673;
   wire n_1_737_674;
   wire n_1_737_675;
   wire n_1_737_676;
   wire n_1_737_677;
   wire n_1_737_678;
   wire n_1_737_679;
   wire n_1_737_680;
   wire n_1_737_681;
   wire n_1_737_682;
   wire n_1_737_683;
   wire n_1_737_684;
   wire n_1_737_685;
   wire n_1_737_686;
   wire n_1_737_687;
   wire n_1_737_688;
   wire n_1_737_689;
   wire n_1_737_690;
   wire n_1_737_691;
   wire n_1_737_692;
   wire n_1_737_693;
   wire n_1_737_694;
   wire n_1_737_695;
   wire n_1_737_696;
   wire n_1_737_697;
   wire n_1_737_698;
   wire n_1_737_699;
   wire n_1_737_700;
   wire n_1_737_701;
   wire n_1_737_702;
   wire n_1_737_703;
   wire n_1_737_704;
   wire n_1_737_705;
   wire n_1_737_706;
   wire n_1_737_707;
   wire n_1_737_708;
   wire n_1_737_709;
   wire n_1_737_710;
   wire n_1_737_711;
   wire n_1_737_712;
   wire n_1_737_713;
   wire n_1_737_714;
   wire n_1_737_715;
   wire n_1_737_716;
   wire n_1_737_717;
   wire n_1_737_718;
   wire n_1_737_719;
   wire n_1_737_720;
   wire n_1_737_721;
   wire n_1_737_722;
   wire n_1_737_723;
   wire n_1_737_724;
   wire n_1_737_725;
   wire n_1_737_726;
   wire n_1_737_727;
   wire n_1_737_728;
   wire n_1_737_729;
   wire n_1_737_730;
   wire n_1_737_731;
   wire n_1_737_732;
   wire n_1_737_733;
   wire n_1_737_734;
   wire n_1_737_735;
   wire n_1_737_736;
   wire n_1_737_737;
   wire n_1_737_738;
   wire n_1_737_739;
   wire n_1_737_740;
   wire n_1_737_741;
   wire n_1_737_742;
   wire n_1_737_743;
   wire n_1_737_744;
   wire n_1_737_745;
   wire n_1_737_746;
   wire n_1_737_747;
   wire n_1_737_748;
   wire n_1_737_749;
   wire n_1_737_750;
   wire n_1_737_751;
   wire n_1_737_752;
   wire n_1_737_753;
   wire n_1_737_754;
   wire n_1_737_755;
   wire n_1_737_756;
   wire n_1_737_757;
   wire n_1_737_758;
   wire n_1_737_759;
   wire n_1_737_760;
   wire n_1_737_761;
   wire n_1_737_762;
   wire n_1_737_763;
   wire n_1_737_764;
   wire n_1_737_765;
   wire n_1_737_766;
   wire n_1_737_767;
   wire n_1_737_768;
   wire n_1_737_769;
   wire n_1_737_770;
   wire n_1_737_771;
   wire n_1_737_772;
   wire n_1_737_773;
   wire n_1_737_774;
   wire n_1_737_775;
   wire n_1_737_776;
   wire n_1_737_777;
   wire n_1_737_778;
   wire n_1_737_779;
   wire n_1_737_780;
   wire n_1_737_781;
   wire n_1_737_782;
   wire n_1_737_783;
   wire n_1_737_784;
   wire n_1_737_785;
   wire n_1_737_786;
   wire n_1_737_787;
   wire n_1_737_788;
   wire n_1_737_789;
   wire n_1_737_790;
   wire n_1_737_791;
   wire n_1_737_792;
   wire n_1_737_793;
   wire n_1_737_794;
   wire n_1_737_795;
   wire n_1_737_796;
   wire n_1_737_797;
   wire n_1_737_798;
   wire n_1_737_799;
   wire n_1_737_800;
   wire n_1_737_801;
   wire n_1_737_802;
   wire n_1_737_803;
   wire n_1_737_804;
   wire n_1_737_805;
   wire n_1_737_806;
   wire n_1_737_807;
   wire n_1_737_808;
   wire n_1_737_809;
   wire n_1_737_810;
   wire n_1_737_811;
   wire n_1_737_812;
   wire n_1_737_813;
   wire n_1_737_814;
   wire n_1_737_815;
   wire n_1_737_816;
   wire n_1_737_817;
   wire n_1_737_818;
   wire n_1_737_819;
   wire n_1_737_820;
   wire n_1_737_821;
   wire n_1_737_822;
   wire n_1_737_823;
   wire n_1_737_824;
   wire n_1_737_825;
   wire n_1_737_826;
   wire n_1_737_827;
   wire n_1_737_828;
   wire n_1_737_829;
   wire n_1_737_830;
   wire n_1_737_831;
   wire n_1_737_832;
   wire n_1_737_833;
   wire n_1_737_834;
   wire n_1_737_835;
   wire n_1_737_836;
   wire n_1_737_837;
   wire n_1_737_838;
   wire n_1_737_839;
   wire n_1_737_840;
   wire n_1_737_841;
   wire n_1_737_842;
   wire n_1_737_843;
   wire n_1_737_844;
   wire n_1_737_845;
   wire n_1_737_846;
   wire n_1_737_847;
   wire n_1_737_848;
   wire n_1_737_849;
   wire n_1_737_850;
   wire n_1_737_851;
   wire n_1_737_852;
   wire n_1_737_853;
   wire n_1_737_854;
   wire n_1_737_855;
   wire n_1_737_856;
   wire n_1_737_857;
   wire n_1_737_858;
   wire n_1_737_859;
   wire n_1_737_860;
   wire n_1_737_861;
   wire n_1_737_862;
   wire n_1_737_863;
   wire n_1_737_864;
   wire n_1_737_865;
   wire n_1_737_866;
   wire n_1_737_867;
   wire n_1_737_868;
   wire n_1_737_869;
   wire n_1_737_870;
   wire n_1_737_871;
   wire n_1_737_872;
   wire n_1_737_873;
   wire n_1_737_874;
   wire n_1_737_875;
   wire n_1_737_876;
   wire n_1_737_877;
   wire n_1_737_878;
   wire n_1_737_879;
   wire n_1_737_880;
   wire n_1_737_881;
   wire n_1_737_882;
   wire n_1_737_883;
   wire n_1_737_884;
   wire n_1_737_885;
   wire n_1_737_886;
   wire n_1_737_887;
   wire n_1_737_888;
   wire n_1_737_889;
   wire n_1_737_890;
   wire n_1_737_891;
   wire n_1_737_892;
   wire n_1_737_893;
   wire n_1_737_894;
   wire n_1_737_895;
   wire n_1_737_896;
   wire n_1_737_897;
   wire n_1_737_898;
   wire n_1_737_899;
   wire n_1_737_900;
   wire n_1_737_901;
   wire n_1_737_902;
   wire n_1_737_903;
   wire n_1_737_904;
   wire n_1_737_905;
   wire n_1_737_906;
   wire n_1_737_907;
   wire n_1_737_908;
   wire n_1_737_909;
   wire n_1_737_910;
   wire n_1_737_911;
   wire n_1_737_912;
   wire n_1_737_913;
   wire n_1_737_914;
   wire n_1_737_915;
   wire n_1_737_916;
   wire n_1_737_917;
   wire n_1_737_918;
   wire n_1_737_919;
   wire n_1_737_920;
   wire n_1_737_921;
   wire n_1_737_922;
   wire n_1_737_923;
   wire n_1_737_924;
   wire n_1_737_925;
   wire n_1_737_926;
   wire n_1_737_927;
   wire n_1_737_928;
   wire n_1_737_929;
   wire n_1_737_930;
   wire n_1_737_931;
   wire n_1_737_932;
   wire n_1_737_933;
   wire n_1_737_934;
   wire n_1_737_935;
   wire n_1_737_936;
   wire n_1_737_937;
   wire n_1_737_938;
   wire n_1_737_939;
   wire n_1_737_940;
   wire n_1_737_941;
   wire n_1_737_942;
   wire n_1_737_943;
   wire n_1_737_944;
   wire n_1_737_945;
   wire n_1_737_946;
   wire n_1_737_947;
   wire n_1_737_948;
   wire n_1_737_949;
   wire n_1_737_950;
   wire n_1_737_951;
   wire n_1_737_952;
   wire n_1_737_953;
   wire n_1_737_954;
   wire n_1_737_955;
   wire n_1_737_956;
   wire n_1_737_957;
   wire n_1_737_958;
   wire n_1_737_959;
   wire n_1_737_960;
   wire n_1_737_961;
   wire n_1_737_962;
   wire n_1_737_963;
   wire n_1_737_964;
   wire n_1_737_965;
   wire n_1_737_966;
   wire n_1_737_967;
   wire n_1_737_968;
   wire n_1_737_969;
   wire n_1_737_970;
   wire n_1_737_971;
   wire n_1_737_972;
   wire n_1_737_973;
   wire n_1_737_974;
   wire n_1_737_975;
   wire n_1_737_976;
   wire n_1_737_977;
   wire n_1_737_978;
   wire n_1_737_979;
   wire n_1_737_980;
   wire n_1_737_981;
   wire n_1_737_982;
   wire n_1_737_983;
   wire n_1_737_984;
   wire n_1_737_985;
   wire n_1_737_986;
   wire n_1_737_987;
   wire n_1_737_988;
   wire n_1_737_989;
   wire n_1_737_990;
   wire n_1_737_991;
   wire n_1_737_992;
   wire n_1_737_993;
   wire n_1_737_994;
   wire n_1_737_995;
   wire n_1_737_996;
   wire n_1_737_997;
   wire n_1_737_998;
   wire n_1_737_999;
   wire n_1_737_1000;
   wire n_1_737_1001;
   wire n_1_737_1002;
   wire n_1_737_1003;
   wire n_1_737_1004;
   wire n_1_737_1005;
   wire n_1_737_1006;
   wire n_1_737_1007;
   wire n_1_737_1008;
   wire n_1_737_1009;
   wire n_1_737_1010;
   wire n_1_737_1011;
   wire n_1_737_1012;
   wire n_1_737_1013;
   wire n_1_737_1014;
   wire n_1_737_1015;
   wire n_1_737_1016;
   wire n_1_737_1017;
   wire n_1_737_1018;
   wire n_1_737_1019;
   wire n_1_737_1020;
   wire n_1_737_1021;
   wire n_1_737_1022;
   wire n_1_737_1023;
   wire n_1_737_1024;
   wire n_1_737_1025;
   wire n_1_737_1026;
   wire n_1_737_1027;
   wire n_1_737_1028;
   wire n_1_737_1029;
   wire n_1_737_1030;
   wire n_1_737_1031;
   wire n_1_737_1032;
   wire n_1_737_1033;
   wire n_1_737_1034;
   wire n_1_737_1035;
   wire n_1_737_1036;
   wire n_1_737_1037;
   wire n_1_737_1038;
   wire n_1_737_1039;
   wire n_1_737_1040;
   wire n_1_737_1041;
   wire n_1_737_1042;
   wire n_1_737_1043;
   wire n_1_737_1044;
   wire n_1_737_1045;
   wire n_1_737_1046;
   wire n_1_737_1047;
   wire n_1_737_1048;
   wire n_1_737_1049;
   wire n_1_737_1050;
   wire n_1_737_1051;
   wire n_1_737_1052;
   wire n_1_737_1053;
   wire n_1_737_1054;
   wire n_1_737_1055;
   wire n_1_737_1056;
   wire n_1_737_1057;
   wire n_1_737_1058;
   wire n_1_737_1059;
   wire n_1_737_1060;
   wire n_1_737_1061;
   wire n_1_737_1062;
   wire n_1_737_1063;
   wire n_1_737_1064;
   wire n_1_737_1065;
   wire n_1_737_1066;
   wire n_1_737_1067;
   wire n_1_737_1068;
   wire n_1_737_1069;
   wire n_1_737_1070;
   wire n_1_737_1071;
   wire n_1_737_1072;
   wire n_1_737_1073;
   wire n_1_737_1074;
   wire n_1_737_1075;
   wire n_1_737_1076;
   wire n_1_737_1077;
   wire n_1_737_1078;
   wire n_1_737_1079;
   wire n_1_737_1080;
   wire n_1_737_1081;
   wire n_1_737_1082;
   wire n_1_737_1083;
   wire n_1_737_1084;
   wire n_1_737_1085;
   wire n_1_737_1086;
   wire n_1_737_1087;
   wire n_1_737_1088;
   wire n_1_737_1089;
   wire n_1_737_1090;
   wire n_1_737_1091;
   wire n_1_737_1092;
   wire n_1_737_1093;
   wire n_1_737_1094;
   wire n_1_737_1095;
   wire n_1_737_1096;
   wire n_1_737_1097;
   wire n_1_737_1098;
   wire n_1_737_1099;
   wire n_1_737_1100;
   wire n_1_737_1101;
   wire n_1_737_1102;
   wire n_1_737_1103;
   wire n_1_737_1104;
   wire n_1_737_1105;
   wire n_1_737_1106;
   wire n_1_737_1107;
   wire n_1_737_1108;
   wire n_1_737_1109;
   wire n_1_737_1110;
   wire n_1_737_1111;
   wire n_1_737_1112;
   wire n_1_737_1113;
   wire n_1_737_1114;
   wire n_1_737_1115;
   wire n_1_737_1116;
   wire n_1_737_1117;
   wire n_1_737_1118;
   wire n_1_737_1119;
   wire n_1_737_1120;
   wire n_1_737_1121;
   wire n_1_737_1122;
   wire n_1_737_1123;
   wire n_1_737_1124;
   wire n_1_737_1125;
   wire n_1_737_1126;
   wire n_1_737_1127;
   wire n_1_737_1128;
   wire n_1_737_1129;
   wire n_1_737_1130;
   wire n_1_737_1131;
   wire n_1_737_1132;
   wire n_1_737_1133;
   wire n_1_737_1134;
   wire n_1_737_1135;
   wire n_1_737_1136;
   wire n_1_737_1137;
   wire n_1_737_1138;
   wire n_1_737_1139;
   wire n_1_737_1140;
   wire n_1_737_1141;
   wire n_1_737_1142;
   wire n_1_737_1143;
   wire n_1_737_1144;
   wire n_1_737_1145;
   wire n_1_737_1146;
   wire n_1_737_1147;
   wire n_1_737_1148;
   wire n_1_737_1149;
   wire n_1_737_1150;
   wire n_1_737_1151;
   wire n_1_737_1152;
   wire n_1_737_1153;
   wire n_1_737_1154;
   wire n_1_737_1155;
   wire n_1_737_1156;
   wire n_1_737_1157;
   wire n_1_737_1158;
   wire n_1_737_1159;
   wire n_1_737_1160;
   wire n_1_737_1161;
   wire n_1_737_1162;
   wire n_1_737_1163;
   wire n_1_737_1164;
   wire n_1_737_1165;
   wire n_1_737_1166;
   wire n_1_737_1167;
   wire n_1_737_1168;
   wire n_1_737_1169;
   wire n_1_737_1170;
   wire n_1_737_1171;
   wire n_1_737_1172;
   wire n_1_737_1173;
   wire n_1_737_1174;
   wire n_1_737_1175;
   wire n_1_737_1176;
   wire n_1_737_1177;
   wire n_1_737_1178;
   wire n_1_737_1179;
   wire n_1_737_1180;
   wire n_1_737_1181;
   wire n_1_737_1182;
   wire n_1_737_1183;
   wire n_1_737_1184;
   wire n_1_737_1185;
   wire n_1_737_1186;
   wire n_1_737_1187;
   wire n_1_737_1188;
   wire n_1_737_1189;
   wire n_1_737_1190;
   wire n_1_737_1191;
   wire n_1_737_1192;
   wire n_1_737_1193;
   wire n_1_737_1194;
   wire n_1_737_1195;
   wire n_1_737_1196;
   wire n_1_737_1197;
   wire n_1_737_1198;
   wire n_1_737_1199;
   wire n_1_737_1200;
   wire n_1_737_1201;
   wire n_1_737_1202;
   wire n_1_737_1203;
   wire n_1_737_1204;
   wire n_1_737_1205;
   wire n_1_737_1206;
   wire n_1_737_1207;
   wire n_1_737_1208;
   wire n_1_737_1209;
   wire n_1_737_1210;
   wire n_1_737_1211;
   wire n_1_737_1212;
   wire n_1_737_1213;
   wire n_1_737_1214;
   wire n_1_737_1215;
   wire n_1_737_1216;
   wire n_1_737_1217;
   wire n_1_737_1218;
   wire n_1_737_1219;
   wire n_1_737_1220;
   wire n_1_737_1221;
   wire n_1_737_1222;
   wire n_1_737_1223;
   wire n_1_737_1224;
   wire n_1_737_1225;
   wire n_1_737_1226;
   wire n_1_737_1227;
   wire n_1_737_1228;
   wire n_1_737_1229;
   wire n_1_737_1230;
   wire n_1_737_1231;
   wire n_1_737_1232;
   wire n_1_737_1233;
   wire n_1_737_1234;
   wire n_1_737_1235;
   wire n_1_737_1236;
   wire n_1_737_1237;
   wire n_1_737_1238;
   wire n_1_737_1239;
   wire n_1_737_1240;
   wire n_1_737_1241;
   wire n_1_737_1242;
   wire n_1_737_1243;
   wire n_1_737_1244;
   wire n_1_737_1245;
   wire n_1_737_1246;
   wire n_1_737_1247;
   wire n_1_737_1248;
   wire n_1_737_1249;
   wire n_1_737_1250;
   wire n_1_737_1251;
   wire n_1_737_1252;
   wire n_1_737_1253;
   wire n_1_737_1254;
   wire n_1_737_1255;
   wire n_1_737_1256;
   wire n_1_737_1257;
   wire n_1_737_1258;
   wire n_1_737_1259;
   wire n_1_737_1260;
   wire n_1_737_1261;
   wire n_1_737_1262;
   wire n_1_737_1263;
   wire n_1_737_1264;
   wire n_1_737_1265;
   wire n_1_737_1266;
   wire n_1_737_1267;
   wire n_1_737_1268;
   wire n_1_737_1269;
   wire n_1_737_1270;
   wire n_1_737_1271;
   wire n_1_737_1272;
   wire n_1_737_1273;
   wire n_1_737_1274;
   wire n_1_737_1275;
   wire n_1_737_1276;
   wire n_1_737_1277;
   wire n_1_737_1278;
   wire n_1_737_1279;
   wire n_1_737_1280;
   wire n_1_737_1281;
   wire n_1_737_1282;
   wire n_1_737_1283;
   wire n_1_737_1284;
   wire n_1_737_1285;
   wire n_1_737_1286;
   wire n_1_737_1287;
   wire n_1_737_1288;
   wire n_1_737_1289;
   wire n_1_737_1290;
   wire n_1_737_1291;
   wire n_1_737_1292;
   wire n_1_737_1293;
   wire n_1_737_1294;
   wire n_1_737_1295;
   wire n_1_737_1296;
   wire n_1_737_1297;
   wire n_1_737_1298;
   wire n_1_737_1299;
   wire n_1_737_1300;
   wire n_1_737_1301;
   wire n_1_737_1302;
   wire n_1_737_1303;
   wire n_1_737_1304;
   wire n_1_737_1305;
   wire n_1_737_1306;
   wire n_1_737_1307;
   wire n_1_737_1308;
   wire n_1_737_1309;
   wire n_1_737_1310;
   wire n_1_737_1311;
   wire n_1_737_1312;
   wire n_1_737_1313;
   wire n_1_737_1314;
   wire n_1_737_1315;
   wire n_1_737_1316;
   wire n_1_737_1317;
   wire n_1_737_1318;
   wire n_1_737_1319;
   wire n_1_737_1320;
   wire n_1_737_1321;
   wire n_1_737_1322;
   wire n_1_737_1323;
   wire n_1_737_1324;
   wire n_1_737_1325;
   wire n_1_737_1326;
   wire n_1_737_1327;
   wire n_1_737_1328;
   wire n_1_737_1329;
   wire n_1_737_1330;
   wire n_1_737_1331;
   wire n_1_737_1332;
   wire n_1_737_1333;
   wire n_1_737_1334;
   wire n_1_737_1335;
   wire n_1_737_1336;
   wire n_1_737_1337;
   wire n_1_737_1338;
   wire n_1_737_1339;
   wire n_1_737_1340;
   wire n_1_737_1341;
   wire n_1_737_1342;
   wire n_1_737_1343;
   wire n_1_737_1344;
   wire n_1_737_1345;
   wire n_1_737_1346;
   wire n_1_737_1347;
   wire n_1_737_1348;
   wire n_1_737_1349;
   wire n_1_737_1350;
   wire n_1_737_1351;
   wire n_1_737_1352;
   wire n_1_737_1353;
   wire n_1_737_1354;
   wire n_1_737_1355;
   wire n_1_737_1356;
   wire n_1_737_1357;
   wire n_1_737_1358;
   wire n_1_737_1359;
   wire n_1_737_1360;
   wire n_1_737_1361;
   wire n_1_737_1362;
   wire n_1_737_1363;
   wire n_1_737_1364;
   wire n_1_737_1365;
   wire n_1_737_1366;
   wire n_1_737_1367;
   wire n_1_737_1368;
   wire n_1_737_1369;
   wire n_1_737_1370;
   wire n_1_737_1371;
   wire n_1_737_1372;
   wire n_1_737_1373;
   wire n_1_737_1374;
   wire n_1_737_1375;
   wire n_1_737_1376;
   wire n_1_737_1377;
   wire n_1_737_1378;
   wire n_1_737_1379;
   wire n_1_737_1380;
   wire n_1_737_1381;
   wire n_1_737_1382;
   wire n_1_737_1383;
   wire n_1_737_1384;
   wire n_1_737_1385;
   wire n_1_737_1386;
   wire n_1_737_1387;
   wire n_1_737_1388;
   wire n_1_737_1389;
   wire n_1_737_1390;
   wire n_1_737_1391;
   wire n_1_737_1392;
   wire n_1_737_1393;
   wire n_1_737_1394;
   wire n_1_737_1395;
   wire n_1_737_1396;
   wire n_1_737_1397;
   wire n_1_737_1398;
   wire n_1_737_1399;
   wire n_1_737_1400;
   wire n_1_737_1401;
   wire n_1_737_1402;
   wire n_1_737_1403;
   wire n_1_737_1404;
   wire n_1_737_1405;
   wire n_1_737_1406;
   wire n_1_737_1407;
   wire n_1_737_1408;
   wire n_1_737_1409;
   wire n_1_737_1410;
   wire n_1_737_1411;
   wire n_1_737_1412;
   wire n_1_737_1413;
   wire n_1_737_1414;
   wire n_1_737_1415;
   wire n_1_737_1416;
   wire n_1_737_1417;
   wire n_1_737_1418;
   wire n_1_737_1419;
   wire n_1_737_1420;
   wire n_1_737_1421;
   wire n_1_737_1422;
   wire n_1_737_1423;
   wire n_1_737_1424;
   wire n_1_737_1425;
   wire n_1_737_1426;
   wire n_1_737_1427;
   wire n_1_737_1428;
   wire n_1_737_1429;
   wire n_1_737_1430;
   wire n_1_737_1431;
   wire n_1_737_1432;
   wire n_1_737_1433;
   wire n_1_737_1434;
   wire n_1_737_1435;
   wire n_1_737_1436;
   wire n_1_737_1437;
   wire n_1_737_1438;
   wire n_1_737_1439;
   wire n_1_737_1440;
   wire n_1_737_1441;
   wire n_1_737_1442;
   wire n_1_737_1443;
   wire n_1_737_1444;
   wire n_1_737_1445;
   wire n_1_737_1446;
   wire n_1_737_1447;
   wire n_1_737_1448;
   wire n_1_737_1449;
   wire n_1_737_1450;
   wire n_1_737_1451;
   wire n_1_737_1452;
   wire n_1_737_1453;
   wire n_1_737_1454;
   wire n_1_737_1455;
   wire n_1_737_1456;
   wire n_1_737_1457;
   wire n_1_737_1458;
   wire n_1_737_1459;
   wire n_1_737_1460;
   wire n_1_737_1461;
   wire n_1_737_1462;
   wire n_1_737_1463;
   wire n_1_737_1464;
   wire n_1_737_1465;
   wire n_1_737_1466;
   wire n_1_737_1467;
   wire n_1_737_1468;
   wire n_1_737_1469;
   wire n_1_737_1470;
   wire n_1_737_1471;
   wire n_1_737_1472;
   wire n_1_737_1473;
   wire n_1_737_1474;
   wire n_1_737_1475;
   wire n_1_737_1476;
   wire n_1_737_1477;
   wire n_1_737_1478;
   wire n_1_737_1479;
   wire n_1_737_1480;
   wire n_1_737_1481;
   wire n_1_737_1482;
   wire n_1_737_1483;
   wire n_1_737_1484;
   wire n_1_737_1485;
   wire n_1_737_1486;
   wire n_1_737_1487;
   wire n_1_737_1488;
   wire n_1_737_1489;
   wire n_1_737_1490;
   wire n_1_737_1491;
   wire n_1_737_1492;
   wire n_1_737_1493;
   wire n_1_737_1494;
   wire n_1_737_1495;
   wire n_1_737_1496;
   wire n_1_737_1497;
   wire n_1_737_1498;
   wire n_1_737_1499;
   wire n_1_737_1500;
   wire n_1_737_1501;
   wire n_1_737_1502;
   wire n_1_737_1503;
   wire n_1_737_1504;
   wire n_1_737_1505;
   wire n_1_737_1506;
   wire n_1_737_1507;
   wire n_1_737_1508;
   wire n_1_737_1509;
   wire n_1_737_1510;
   wire n_1_737_1511;
   wire n_1_737_1512;
   wire n_1_737_1513;
   wire n_1_737_1514;
   wire n_1_737_1515;
   wire n_1_737_1516;
   wire n_1_737_1517;
   wire n_1_737_1518;
   wire n_1_737_1519;
   wire n_1_737_1520;
   wire n_1_737_1521;
   wire n_1_737_1522;
   wire n_1_737_1523;
   wire n_1_737_1524;
   wire n_1_737_1525;
   wire n_1_737_1526;
   wire n_1_737_1527;
   wire n_1_737_1528;
   wire n_1_737_1529;
   wire n_1_737_1530;
   wire n_1_737_1531;
   wire n_1_737_1532;
   wire n_1_737_1533;
   wire n_1_737_1534;
   wire n_1_737_1535;
   wire n_1_737_1536;
   wire n_1_737_1537;
   wire n_1_737_1538;
   wire n_1_737_1539;
   wire n_1_737_1540;
   wire n_1_737_1541;
   wire n_1_737_1542;
   wire n_1_737_1543;
   wire n_1_737_1544;
   wire n_1_737_1545;
   wire n_1_737_1546;
   wire n_1_737_1547;
   wire n_1_737_1548;
   wire n_1_737_1549;
   wire n_1_737_1550;
   wire n_1_737_1551;
   wire n_1_737_1552;
   wire n_1_737_1553;
   wire n_1_737_1554;
   wire n_1_737_1555;
   wire n_1_737_1556;
   wire n_1_737_1557;
   wire n_1_737_1558;
   wire n_1_737_1559;
   wire n_1_737_1560;
   wire n_1_737_1561;
   wire n_1_737_1562;
   wire n_1_737_1563;
   wire n_1_737_1564;
   wire n_1_737_1565;
   wire n_1_737_1566;
   wire n_1_737_1567;
   wire n_1_737_1568;
   wire n_1_737_1569;
   wire n_1_737_1570;
   wire n_1_737_1571;
   wire n_1_737_1572;
   wire n_1_737_1573;
   wire n_1_737_1574;
   wire n_1_737_1575;
   wire n_1_737_1576;
   wire n_1_737_1577;
   wire n_1_737_1578;
   wire n_1_737_1579;
   wire n_1_737_1580;
   wire n_1_737_1581;
   wire n_1_737_1582;
   wire n_1_737_1583;
   wire n_1_737_1584;
   wire n_1_737_1585;
   wire n_1_737_1586;
   wire n_1_737_1587;
   wire n_1_737_1588;
   wire n_1_737_1589;
   wire n_1_737_1590;
   wire n_1_737_1591;
   wire n_1_737_1592;
   wire n_1_737_1593;
   wire n_1_737_1594;
   wire n_1_737_1595;
   wire n_1_737_1596;
   wire n_1_737_1597;
   wire n_1_737_1598;
   wire n_1_737_1599;
   wire n_1_737_1600;
   wire n_1_737_1601;
   wire n_1_737_1602;
   wire n_1_737_1603;
   wire n_1_737_1604;
   wire n_1_737_1605;
   wire n_1_737_1606;
   wire n_1_737_1607;
   wire n_1_737_1608;
   wire n_1_737_1609;
   wire n_1_737_1610;
   wire n_1_737_1611;
   wire n_1_737_1612;
   wire n_1_737_1613;
   wire n_1_737_1614;
   wire n_1_737_1615;
   wire n_1_737_1616;
   wire n_1_737_1617;
   wire n_1_737_1618;
   wire n_1_737_1619;
   wire n_1_737_1620;
   wire n_1_737_1621;
   wire n_1_737_1622;
   wire n_1_737_1623;
   wire n_1_737_1624;
   wire n_1_737_1625;
   wire n_1_737_1626;
   wire n_1_737_1627;
   wire n_1_737_1628;
   wire n_1_737_1629;
   wire n_1_737_1630;
   wire n_1_737_1631;
   wire n_1_737_1632;
   wire n_1_737_1633;
   wire n_1_737_1634;
   wire n_1_737_1635;
   wire n_1_737_1636;
   wire n_1_737_1637;
   wire n_1_737_1638;
   wire n_1_737_1639;
   wire n_1_737_1640;
   wire n_1_737_1641;
   wire n_1_737_1642;
   wire n_1_737_1643;
   wire n_1_737_1644;
   wire n_1_737_1645;
   wire n_1_737_1646;
   wire n_1_737_1647;
   wire n_1_737_1648;
   wire n_1_737_1649;
   wire n_1_737_1650;
   wire n_1_737_1651;
   wire n_1_737_1652;
   wire n_1_737_1653;
   wire n_1_737_1654;
   wire n_1_737_1655;
   wire n_1_737_1656;
   wire n_1_737_1657;
   wire n_1_737_1658;
   wire n_1_737_1659;
   wire n_1_737_1660;
   wire n_1_737_1661;
   wire n_1_737_1662;
   wire n_1_737_1663;
   wire n_1_737_1664;
   wire n_1_737_1665;
   wire n_1_737_1666;
   wire n_1_737_1667;
   wire n_1_737_1668;
   wire n_1_737_1669;
   wire n_1_737_1670;
   wire n_1_737_1671;
   wire n_1_737_1672;
   wire n_1_737_1673;
   wire n_1_737_1674;
   wire n_1_737_1675;
   wire n_1_737_1676;
   wire n_1_737_1677;
   wire n_1_737_1678;
   wire n_1_737_1679;
   wire n_1_737_1680;
   wire n_1_737_1681;
   wire n_1_737_1682;
   wire n_1_737_1683;
   wire n_1_737_1684;
   wire n_1_737_1685;
   wire n_1_737_1686;
   wire n_1_737_1687;
   wire n_1_737_1688;
   wire n_1_737_1689;
   wire n_1_737_1690;
   wire n_1_737_1691;
   wire n_1_737_1692;
   wire n_1_737_1693;
   wire n_1_737_1694;
   wire n_1_737_1695;
   wire n_1_737_1696;
   wire n_1_737_1697;
   wire n_1_737_1698;
   wire n_1_737_1699;
   wire n_1_737_1700;
   wire n_1_737_1701;
   wire n_1_737_1702;
   wire n_1_737_1703;
   wire n_1_737_1704;
   wire n_1_737_1705;
   wire n_1_737_1706;
   wire n_1_737_1707;
   wire n_1_737_1708;
   wire n_1_737_1709;
   wire n_1_737_1710;
   wire n_1_737_1711;
   wire n_1_737_1712;
   wire n_1_737_1713;
   wire n_1_737_1714;
   wire n_1_737_1715;
   wire n_1_737_1716;
   wire n_1_737_1717;
   wire n_1_737_1718;
   wire n_1_737_1719;
   wire n_1_737_1720;
   wire n_1_737_1721;
   wire n_1_737_1722;
   wire n_1_737_1723;
   wire n_1_737_1724;
   wire n_1_737_1725;
   wire n_1_737_1726;
   wire n_1_737_1727;
   wire n_1_737_1728;
   wire n_1_737_1729;
   wire n_1_737_1730;
   wire n_1_737_1731;
   wire n_1_737_1732;
   wire n_1_737_1733;
   wire n_1_737_1734;
   wire n_1_737_1735;
   wire n_1_737_1736;
   wire n_1_737_1737;
   wire n_1_737_1738;
   wire n_1_737_1739;
   wire n_1_737_1740;
   wire n_1_737_1741;
   wire n_1_737_1742;
   wire n_1_737_1743;
   wire n_1_737_1744;
   wire n_1_737_1745;
   wire n_1_737_1746;
   wire n_1_737_1747;
   wire n_1_737_1748;
   wire n_1_737_1749;
   wire n_1_737_1750;
   wire n_1_737_1751;
   wire n_1_737_1752;
   wire n_1_737_1753;
   wire n_1_737_1754;
   wire n_1_737_1755;
   wire n_1_737_1756;
   wire n_1_737_1757;
   wire n_1_737_1758;
   wire n_1_737_1759;
   wire n_1_737_1760;
   wire n_1_737_1761;
   wire n_1_737_1762;
   wire n_1_737_1763;
   wire n_1_737_1764;
   wire n_1_737_1765;
   wire n_1_737_1766;
   wire n_1_737_1767;
   wire n_1_737_1768;
   wire n_1_737_1769;
   wire n_1_737_1770;
   wire n_1_737_1771;
   wire n_1_737_1772;
   wire n_1_737_1773;
   wire n_1_737_1774;
   wire n_1_737_1775;
   wire n_1_737_1776;
   wire n_1_737_1777;
   wire n_1_737_1778;
   wire n_1_737_1779;
   wire n_1_737_1780;
   wire n_1_737_1781;
   wire n_1_737_1782;
   wire n_1_737_1783;
   wire n_1_737_1784;
   wire n_1_737_1785;
   wire n_1_737_1786;
   wire n_1_737_1787;
   wire n_1_737_1788;
   wire n_1_737_1789;
   wire n_1_737_1790;
   wire n_1_737_1791;
   wire n_1_737_1792;
   wire n_1_737_1793;
   wire n_1_737_1794;
   wire n_1_737_1795;
   wire n_1_737_1796;
   wire n_1_737_1797;
   wire n_1_737_1798;
   wire n_1_737_1799;
   wire n_1_737_1800;
   wire n_1_737_1801;
   wire n_1_737_1802;
   wire n_1_737_1803;
   wire n_1_737_1804;
   wire n_1_737_1805;
   wire n_1_737_1806;
   wire n_1_737_1807;
   wire n_1_737_1808;
   wire n_1_737_1809;
   wire n_1_737_1810;
   wire n_1_737_1811;
   wire n_1_737_1812;
   wire n_1_737_1813;
   wire n_1_737_1814;
   wire n_1_737_1815;
   wire n_1_737_1816;
   wire n_1_737_1817;
   wire n_1_737_1818;
   wire n_1_737_1819;
   wire n_1_737_1820;
   wire n_1_737_1821;
   wire n_1_737_1822;
   wire n_1_737_1823;
   wire n_1_737_1824;
   wire n_1_737_1825;
   wire n_1_737_1826;
   wire n_1_737_1827;
   wire n_1_737_1828;
   wire n_1_737_1829;
   wire n_1_737_1830;
   wire n_1_737_1831;
   wire n_1_737_1832;
   wire n_1_737_1833;
   wire n_1_737_1834;
   wire n_1_737_1835;
   wire n_1_737_1836;
   wire n_1_737_1837;
   wire n_1_737_1838;
   wire n_1_737_1839;
   wire n_1_737_1840;
   wire n_1_737_1841;
   wire n_1_737_1842;
   wire n_1_737_1843;
   wire n_1_737_1844;
   wire n_1_737_1845;
   wire n_1_737_1846;
   wire n_1_737_1847;
   wire n_1_737_1848;
   wire n_1_737_1849;
   wire n_1_737_1850;
   wire n_1_737_1851;
   wire n_1_737_1852;
   wire n_1_737_1853;
   wire n_1_737_1854;
   wire n_1_737_1855;
   wire n_1_737_1856;
   wire n_1_737_1857;
   wire n_1_737_1858;
   wire n_1_737_1859;
   wire n_1_737_1860;
   wire n_1_737_1861;
   wire n_1_737_1862;
   wire n_1_737_1863;
   wire n_1_737_1864;
   wire n_1_737_1865;
   wire n_1_737_1866;
   wire n_1_737_1867;
   wire n_1_737_1868;
   wire n_1_737_1869;
   wire n_1_737_1872;
   wire n_1_737_1873;
   wire n_1_737_1876;
   wire n_1_737_1877;
   wire n_1_737_1878;
   wire n_1_737_1879;
   wire n_1_737_1880;
   wire n_1_737_1881;
   wire n_1_737_1882;
   wire n_1_737_1883;
   wire n_1_737_1884;
   wire n_1_737_1885;
   wire n_1_737_1886;
   wire n_1_737_1887;
   wire n_1_737_1888;
   wire n_1_737_1889;
   wire n_1_737_1890;
   wire n_1_737_1891;
   wire n_1_737_1892;
   wire n_1_737_1893;
   wire n_1_737_1894;
   wire n_1_737_1895;
   wire n_1_737_1896;
   wire n_1_737_1897;
   wire n_1_737_1898;
   wire n_1_737_1899;
   wire n_1_737_1900;
   wire n_1_737_1901;
   wire n_1_737_1902;
   wire n_1_737_1903;
   wire n_1_737_1904;
   wire n_1_737_1905;
   wire n_1_737_1906;
   wire n_1_737_1907;
   wire n_1_737_1908;
   wire n_1_737_1909;
   wire n_1_737_1910;
   wire n_1_737_1911;
   wire n_1_737_1912;
   wire n_1_737_1913;
   wire n_1_737_1914;
   wire n_1_737_1915;
   wire n_1_737_1916;
   wire n_1_737_1917;
   wire n_1_737_1918;
   wire n_1_737_1919;
   wire n_1_737_1920;
   wire n_1_737_1921;
   wire n_1_737_1922;
   wire n_1_737_1923;
   wire n_1_737_1924;
   wire n_1_737_1925;
   wire n_1_737_1926;
   wire n_1_737_1927;
   wire n_1_737_1928;
   wire n_1_737_1929;
   wire n_1_737_1930;
   wire n_1_737_1931;
   wire n_1_737_1932;
   wire n_1_737_1933;
   wire n_1_737_1934;
   wire n_1_737_1935;
   wire n_1_737_1936;
   wire n_1_737_1937;
   wire n_1_737_1938;
   wire n_1_737_1939;
   wire n_1_737_1940;
   wire n_1_737_1941;
   wire n_1_737_1942;
   wire n_1_737_1943;
   wire n_1_737_1944;
   wire n_1_737_1945;
   wire n_1_737_1946;
   wire n_1_737_1947;
   wire n_1_737_1948;
   wire n_1_737_1949;
   wire n_1_737_1950;
   wire n_1_737_1951;
   wire n_1_737_1952;
   wire n_1_737_1953;
   wire n_1_737_1954;
   wire n_1_737_1955;
   wire n_1_737_1956;
   wire n_1_737_1957;
   wire n_1_737_1958;
   wire n_1_737_1959;
   wire n_1_737_1960;
   wire n_1_737_1961;
   wire n_1_737_1962;
   wire n_1_737_1963;
   wire n_1_737_1964;
   wire n_1_737_1965;
   wire n_1_737_1966;
   wire n_1_737_1967;
   wire n_1_737_1968;
   wire n_1_737_1972;
   wire n_1_737_1974;
   wire n_1_737_1975;
   wire n_1_737_1977;
   wire n_1_737_1980;
   wire n_1_737_1981;
   wire n_1_737_1982;
   wire n_1_737_1983;
   wire n_1_737_1984;
   wire n_1_737_1985;
   wire n_1_737_1986;
   wire n_1_737_1987;
   wire n_1_737_1988;
   wire n_1_737_1989;
   wire n_1_737_1990;
   wire n_1_737_1991;
   wire n_1_737_1992;
   wire n_1_737_1993;
   wire n_1_737_1994;
   wire n_1_737_1995;
   wire n_1_737_1996;
   wire n_1_737_1997;
   wire n_1_737_1998;
   wire n_1_737_1999;
   wire n_1_737_2000;
   wire n_1_737_2001;
   wire n_1_737_2002;
   wire n_1_737_2003;
   wire n_1_737_2004;
   wire n_1_737_2005;
   wire n_1_737_2006;
   wire n_1_737_2007;
   wire n_1_737_2008;
   wire n_1_737_2009;
   wire n_1_737_2010;
   wire n_1_737_2011;
   wire n_1_737_2012;
   wire n_1_737_2013;
   wire n_1_737_2014;
   wire n_1_737_2015;
   wire n_1_737_2016;
   wire n_1_737_2017;
   wire n_1_737_2018;
   wire n_1_737_2019;
   wire n_1_737_2020;
   wire n_1_737_2021;
   wire n_1_737_2022;
   wire n_1_737_2023;
   wire n_1_737_2024;
   wire n_1_737_2025;
   wire n_1_737_2026;
   wire n_1_737_2027;
   wire n_1_737_2028;
   wire n_1_737_2029;
   wire n_1_737_2030;
   wire n_1_737_2031;
   wire n_1_737_2032;
   wire n_1_737_2033;
   wire n_1_737_2034;
   wire n_1_737_2035;
   wire n_1_737_2036;
   wire n_1_737_2037;
   wire n_1_737_2038;
   wire n_1_737_2039;
   wire n_1_737_2040;
   wire n_1_737_2041;
   wire n_1_737_2042;
   wire n_1_737_2043;
   wire n_1_737_2044;
   wire n_1_737_2045;
   wire n_1_737_2046;
   wire n_1_737_2047;
   wire n_1_737_2048;
   wire n_1_737_2049;
   wire n_1_737_2050;
   wire n_1_737_2051;
   wire n_1_737_2052;
   wire n_1_737_2053;
   wire n_1_737_2054;
   wire n_1_737_2055;
   wire n_1_737_2056;
   wire n_1_737_2057;
   wire n_1_737_2058;
   wire n_1_737_2059;
   wire n_1_737_2060;
   wire n_1_737_2061;
   wire n_1_737_2062;
   wire n_1_737_2063;
   wire n_1_737_2064;
   wire n_1_737_2065;
   wire n_1_737_2066;
   wire n_1_737_2067;
   wire n_1_737_2068;
   wire n_1_737_2069;
   wire n_1_737_2070;
   wire n_1_737_2071;
   wire n_1_737_2072;
   wire n_1_737_2073;
   wire n_1_737_2074;
   wire n_1_737_2075;
   wire n_1_737_2076;
   wire n_1_737_2077;
   wire n_1_737_2078;
   wire n_1_737_2079;
   wire n_1_737_2080;
   wire n_1_737_2081;
   wire n_1_737_2082;
   wire n_1_737_2083;
   wire n_1_737_2084;
   wire n_1_737_2085;
   wire n_1_737_2086;
   wire n_1_737_2087;
   wire n_1_737_2088;
   wire n_1_737_2089;
   wire n_1_737_2090;
   wire n_1_737_2091;
   wire n_1_737_2092;
   wire n_1_737_2093;
   wire n_1_737_2094;
   wire n_1_737_2095;
   wire n_1_737_2096;
   wire n_1_737_2097;
   wire n_1_737_2098;
   wire n_1_737_2099;
   wire n_1_737_2100;
   wire n_1_737_2101;
   wire n_1_737_2102;
   wire n_1_737_2103;
   wire n_1_737_2104;
   wire n_1_737_2105;
   wire n_1_737_2106;
   wire n_1_737_2107;
   wire n_1_737_2108;
   wire n_1_737_2109;
   wire n_1_737_2110;
   wire n_1_737_2111;
   wire n_1_737_2112;
   wire n_1_737_2113;
   wire n_1_737_2114;
   wire n_1_737_2115;
   wire n_1_737_2116;
   wire n_1_737_2117;
   wire n_1_737_2118;
   wire n_1_737_2119;
   wire n_1_737_2120;
   wire n_1_737_2121;
   wire n_1_737_2122;
   wire n_1_737_2123;
   wire n_1_737_2124;
   wire n_1_737_2125;
   wire n_1_737_2126;
   wire n_1_737_2127;
   wire n_1_737_2128;
   wire n_1_737_2129;
   wire n_1_737_2130;
   wire n_1_737_2131;
   wire n_1_737_2132;
   wire n_1_737_2133;
   wire n_1_737_2134;
   wire n_1_737_2135;
   wire n_1_737_2136;
   wire n_1_737_2137;
   wire n_1_737_2138;
   wire n_1_737_2139;
   wire n_1_737_2140;
   wire n_1_737_2141;
   wire n_1_737_2142;
   wire n_1_737_2143;
   wire n_1_737_2144;
   wire n_1_737_2145;
   wire n_1_737_2146;
   wire n_1_737_2147;
   wire n_1_737_2148;
   wire n_1_737_2149;
   wire n_1_737_2150;
   wire n_1_737_2151;
   wire n_1_737_2152;
   wire n_1_737_2153;
   wire n_1_737_2154;
   wire n_1_737_2155;
   wire n_1_737_2156;
   wire n_1_737_2157;
   wire n_1_737_2158;
   wire n_1_737_2159;
   wire n_1_737_2160;
   wire n_1_737_2161;
   wire n_1_737_2162;
   wire n_1_737_2163;
   wire n_1_737_2164;
   wire n_1_737_2165;
   wire n_1_737_2166;
   wire n_1_737_2167;
   wire n_1_737_2168;
   wire n_1_737_2169;
   wire n_1_737_2170;
   wire n_1_737_2171;
   wire n_1_737_2172;
   wire n_1_737_2173;
   wire n_1_737_2174;
   wire n_1_737_2175;
   wire n_1_737_2176;
   wire n_1_737_2177;
   wire n_1_737_2178;
   wire n_1_737_2179;
   wire n_1_737_2180;
   wire n_1_737_2181;
   wire n_1_737_2182;
   wire n_1_737_2183;
   wire n_1_737_2184;
   wire n_1_737_2185;
   wire n_1_737_2186;
   wire n_1_737_2187;
   wire n_1_737_2188;
   wire n_1_737_2189;
   wire n_1_737_2190;
   wire n_1_737_2191;
   wire n_1_737_2192;
   wire n_1_737_2193;
   wire n_1_737_2194;
   wire n_1_737_2195;
   wire n_1_737_2196;
   wire n_1_737_2197;
   wire n_1_737_2198;
   wire n_1_737_2199;
   wire n_1_737_2200;
   wire n_1_737_2201;
   wire n_1_737_2202;
   wire n_1_737_2203;
   wire n_1_737_2204;
   wire n_1_737_2205;
   wire n_1_737_2206;
   wire n_1_737_2207;
   wire n_1_737_2208;
   wire n_1_737_2209;
   wire n_1_737_2210;
   wire n_1_737_2211;
   wire n_1_737_2212;
   wire n_1_737_2213;
   wire n_1_737_2214;
   wire n_1_737_2215;
   wire n_1_737_2216;
   wire n_1_737_2217;
   wire n_1_737_2218;
   wire n_1_737_2219;
   wire n_1_737_2220;
   wire n_1_737_2221;
   wire n_1_737_2222;
   wire n_1_737_2223;
   wire n_1_737_2224;
   wire n_1_737_2225;
   wire n_1_737_2226;
   wire n_1_737_2227;
   wire n_1_737_2228;
   wire n_1_737_2229;
   wire n_1_737_2230;
   wire n_1_737_2231;
   wire n_1_737_2232;
   wire n_1_737_2233;
   wire n_1_737_2234;
   wire n_1_737_2235;
   wire n_1_737_2236;
   wire n_1_737_2237;
   wire n_1_737_2238;
   wire n_1_737_2239;
   wire n_1_737_2240;
   wire n_1_737_2241;
   wire n_1_737_2242;
   wire n_1_737_2243;
   wire n_1_737_2244;
   wire n_1_737_2245;
   wire n_1_737_2246;
   wire n_1_737_2247;
   wire n_1_737_2248;
   wire n_1_737_2249;
   wire n_1_737_2250;
   wire n_1_737_2251;
   wire n_1_737_2252;
   wire n_1_737_2253;
   wire n_1_737_2254;
   wire n_1_737_2255;
   wire n_1_737_2256;
   wire n_1_737_2257;
   wire n_1_737_2258;
   wire n_1_737_2259;
   wire n_1_737_2260;
   wire n_1_737_2261;
   wire n_1_737_2262;
   wire n_1_737_2263;
   wire n_1_737_2264;
   wire n_1_737_2265;
   wire n_1_737_2266;
   wire n_1_737_2267;
   wire n_1_737_2268;
   wire n_1_737_2269;
   wire n_1_737_2270;
   wire n_1_737_2271;
   wire n_1_737_2272;
   wire n_1_737_2273;
   wire n_1_737_2274;
   wire n_1_737_2275;
   wire n_1_737_2276;
   wire n_1_737_2277;
   wire n_1_737_2278;
   wire n_1_737_2279;
   wire n_1_737_2280;
   wire n_1_737_2281;
   wire n_1_737_2282;
   wire n_1_737_2283;
   wire n_1_737_2284;
   wire n_1_737_2285;
   wire n_1_737_2286;
   wire n_1_737_2287;
   wire n_1_737_2288;
   wire n_1_737_2289;
   wire n_1_737_2290;
   wire n_1_737_2291;
   wire n_1_737_2292;
   wire n_1_737_2293;
   wire n_1_737_2294;
   wire n_1_737_2295;
   wire n_1_737_2296;
   wire n_1_737_2297;
   wire n_1_737_2298;
   wire n_1_737_2299;
   wire n_1_737_2300;
   wire n_1_737_2301;
   wire n_1_737_2302;
   wire n_1_737_2303;
   wire n_1_737_2304;
   wire n_1_737_2305;
   wire n_1_737_2306;
   wire n_1_737_2307;
   wire n_1_737_2308;
   wire n_1_737_2309;
   wire n_1_737_2310;
   wire n_1_737_2311;
   wire n_1_737_2312;
   wire n_1_737_2313;
   wire n_1_737_2314;
   wire n_1_737_2315;
   wire n_1_737_2316;
   wire n_1_737_2317;
   wire n_1_737_2318;
   wire n_1_737_2319;
   wire n_1_737_2320;
   wire n_1_737_2321;
   wire n_1_737_2322;
   wire n_1_737_2323;
   wire n_1_737_2324;
   wire n_1_737_2325;
   wire n_1_737_2326;
   wire n_1_737_2327;
   wire n_1_737_2328;
   wire n_1_737_2329;
   wire n_1_737_2330;
   wire n_1_737_2331;
   wire n_1_737_2332;
   wire n_1_737_2333;
   wire n_1_737_2334;
   wire n_1_737_2335;
   wire n_1_737_2336;
   wire n_1_737_2337;
   wire n_1_737_2338;
   wire n_1_737_2339;
   wire n_1_737_2340;
   wire n_1_737_2341;
   wire n_1_737_2342;
   wire n_1_737_2343;
   wire n_1_737_2344;
   wire n_1_737_2345;
   wire n_1_737_2346;
   wire n_1_737_2347;
   wire n_1_737_2348;
   wire n_1_737_2349;
   wire n_1_737_2350;
   wire n_1_737_2351;
   wire n_1_737_2352;
   wire n_1_737_2353;
   wire n_1_737_2354;
   wire n_1_737_2355;
   wire n_1_737_2356;
   wire n_1_737_2357;
   wire n_1_737_2358;
   wire n_1_737_2359;
   wire n_1_737_2360;
   wire n_1_737_2361;
   wire n_1_737_2362;
   wire n_1_737_2363;
   wire n_1_737_2364;
   wire n_1_737_2365;
   wire n_1_737_2366;
   wire n_1_737_2367;
   wire n_1_737_2368;
   wire n_1_737_2369;
   wire n_1_737_2370;
   wire n_1_737_2371;
   wire n_1_737_2372;
   wire n_1_737_2373;
   wire n_1_737_2374;
   wire n_1_737_2375;
   wire n_1_737_2376;
   wire n_1_737_2377;
   wire n_1_737_2378;
   wire n_1_737_2379;
   wire n_1_737_2380;
   wire n_1_737_2381;
   wire n_1_737_2382;
   wire n_1_737_2383;
   wire n_1_737_2384;
   wire n_1_737_2385;
   wire n_1_737_2386;
   wire n_1_737_2387;
   wire n_1_737_2388;
   wire n_1_737_2389;
   wire n_1_737_2390;
   wire n_1_737_2391;
   wire n_1_737_2392;
   wire n_1_737_2393;
   wire n_1_737_2394;
   wire n_1_737_2395;
   wire n_1_737_2396;
   wire n_1_737_2397;
   wire n_1_737_2398;
   wire n_1_737_2399;
   wire n_1_737_2400;
   wire n_1_737_2401;
   wire n_1_737_2402;
   wire n_1_737_2403;
   wire n_1_737_2404;
   wire n_1_737_2405;
   wire n_1_737_2406;
   wire n_1_737_2407;
   wire n_1_737_2408;
   wire n_1_737_2409;
   wire n_1_737_2410;
   wire n_1_737_2411;
   wire n_1_737_2412;
   wire n_1_737_2413;
   wire n_1_737_2414;
   wire n_1_737_2415;
   wire n_1_737_2416;
   wire n_1_737_2417;
   wire n_1_737_2418;
   wire n_1_737_2419;
   wire n_1_737_2420;
   wire n_1_737_2421;
   wire n_1_737_2422;
   wire n_1_737_2423;
   wire n_1_737_2424;
   wire n_1_737_2425;
   wire n_1_737_2426;
   wire n_1_737_2427;
   wire n_1_737_2428;
   wire n_1_737_2429;
   wire n_1_737_2430;
   wire n_1_737_2431;
   wire n_1_737_2432;
   wire n_1_737_2433;
   wire n_1_737_2434;
   wire n_1_737_2435;
   wire n_1_737_2436;
   wire n_1_737_2437;
   wire n_1_737_2438;
   wire n_1_737_2439;
   wire n_1_737_2440;
   wire n_1_737_2441;
   wire n_1_737_2442;
   wire n_1_737_2443;
   wire n_1_737_2444;
   wire n_1_737_2445;
   wire n_1_737_2446;
   wire n_1_737_2447;
   wire n_1_737_2448;
   wire n_1_737_2449;
   wire n_1_737_2450;
   wire n_1_737_2451;
   wire n_1_737_2452;
   wire n_1_737_2453;
   wire n_1_737_2454;
   wire n_1_737_2455;
   wire n_1_737_2456;
   wire n_1_737_2457;
   wire n_1_737_2458;
   wire n_1_737_2459;
   wire n_1_737_2460;
   wire n_1_737_2461;
   wire n_1_737_2462;
   wire n_1_737_2463;
   wire n_1_737_2464;
   wire n_1_737_2465;
   wire n_1_737_2466;
   wire n_1_737_2467;
   wire n_1_737_2468;
   wire n_1_737_2469;
   wire n_1_737_2470;
   wire n_1_737_2471;
   wire n_1_737_2472;
   wire n_1_737_2473;
   wire n_1_737_2474;
   wire n_1_737_2475;
   wire n_1_737_2476;
   wire n_1_737_2477;
   wire n_1_737_2478;
   wire n_1_737_2479;
   wire n_1_737_2480;
   wire n_1_737_2481;
   wire n_1_737_2482;
   wire n_1_737_2483;
   wire n_1_737_2484;
   wire n_1_737_2485;
   wire n_1_737_2486;
   wire n_1_737_2487;
   wire n_1_737_2488;
   wire n_1_737_2489;
   wire n_1_737_2490;
   wire n_1_737_2491;
   wire n_1_737_2492;
   wire n_1_737_2493;
   wire n_1_737_2494;
   wire n_1_737_2495;
   wire n_1_737_2496;
   wire n_1_737_2497;
   wire n_1_737_2498;
   wire n_1_737_2499;
   wire n_1_737_2500;
   wire n_1_737_2501;
   wire n_1_737_2502;
   wire n_1_737_2503;
   wire n_1_737_2504;
   wire n_1_737_2505;
   wire n_1_737_2506;
   wire n_1_737_2507;
   wire n_1_737_2508;
   wire n_1_737_2509;
   wire n_1_737_2510;
   wire n_1_737_2511;
   wire n_1_737_2512;
   wire n_1_737_2513;
   wire n_1_737_2514;
   wire n_1_737_2515;
   wire n_1_737_2516;
   wire n_1_737_2517;
   wire n_1_737_2518;
   wire n_1_737_2519;
   wire n_1_737_2520;
   wire n_1_737_2521;
   wire n_1_737_2522;
   wire n_1_737_2523;
   wire n_1_737_2524;
   wire n_1_737_2525;
   wire n_1_737_2526;
   wire n_1_737_2527;
   wire n_1_737_2528;
   wire n_1_737_2529;
   wire n_1_737_2530;
   wire n_1_737_2531;
   wire n_1_737_2532;
   wire n_1_737_2533;
   wire n_1_737_2534;
   wire n_1_737_2535;
   wire n_1_737_2536;
   wire n_1_737_2537;
   wire n_1_737_2538;
   wire n_1_737_2539;
   wire n_1_737_2540;
   wire n_1_737_2541;
   wire n_1_737_2542;
   wire n_1_737_2543;
   wire n_1_737_2544;
   wire n_1_737_2545;
   wire n_1_737_2546;
   wire n_1_737_2547;
   wire n_1_737_2548;
   wire n_1_737_2549;
   wire n_1_737_2550;
   wire n_1_737_2551;
   wire n_1_737_2552;
   wire n_1_737_2553;
   wire n_1_737_2554;
   wire n_1_737_2555;
   wire n_1_737_2556;
   wire n_1_737_2557;
   wire n_1_737_2558;
   wire n_1_737_2559;
   wire n_1_737_2560;
   wire n_1_737_2561;
   wire n_1_737_2562;
   wire n_1_737_2563;
   wire n_1_737_2564;
   wire n_1_737_2565;
   wire n_1_737_2566;
   wire n_1_737_2567;
   wire n_1_737_2568;
   wire n_1_737_2569;
   wire n_1_737_2570;
   wire n_1_737_2571;
   wire n_1_737_2572;
   wire n_1_737_2573;
   wire n_1_737_2574;
   wire n_1_737_2575;
   wire n_1_737_2576;
   wire n_1_737_2577;
   wire n_1_737_2578;
   wire n_1_737_2579;
   wire n_1_737_2580;
   wire n_1_737_2581;
   wire n_1_737_2582;
   wire n_1_737_2583;
   wire n_1_737_2584;
   wire n_1_737_2585;
   wire n_1_737_2586;
   wire n_1_737_2587;
   wire n_1_737_2588;
   wire n_1_737_2589;
   wire n_1_737_2590;
   wire n_1_737_2591;
   wire n_1_737_2592;
   wire n_1_737_2593;
   wire n_1_737_2594;
   wire n_1_737_2595;
   wire n_1_737_2596;
   wire n_1_737_2597;
   wire n_1_737_2598;
   wire n_1_737_2599;
   wire n_1_737_2600;
   wire n_1_737_2601;
   wire n_1_737_2602;
   wire n_1_737_2603;
   wire n_1_737_2604;
   wire n_1_737_2605;
   wire n_1_737_2606;
   wire n_1_737_2607;
   wire n_1_737_2608;
   wire n_1_737_2609;
   wire n_1_737_2610;
   wire n_1_737_2611;
   wire n_1_737_2612;
   wire n_1_737_2613;
   wire n_1_737_2614;
   wire n_1_737_2615;
   wire n_1_737_2616;
   wire n_1_737_2617;
   wire n_1_737_2618;
   wire n_1_737_2619;
   wire n_1_737_2620;
   wire n_1_737_2621;
   wire n_1_737_2622;
   wire n_1_737_2623;
   wire n_1_737_2624;
   wire n_1_737_2625;
   wire n_1_737_2626;
   wire n_1_737_2627;
   wire n_1_737_2628;
   wire n_1_737_2629;
   wire n_1_737_2630;
   wire n_1_737_2631;
   wire n_1_737_2632;
   wire n_1_737_2633;
   wire n_1_737_2634;
   wire n_1_737_2635;
   wire n_1_737_2636;
   wire n_1_737_2637;
   wire n_1_737_2638;
   wire n_1_737_2639;
   wire n_1_737_2640;
   wire n_1_737_2641;
   wire n_1_737_2642;
   wire n_1_737_2643;
   wire n_1_737_2644;
   wire n_1_737_2645;
   wire n_1_737_2646;
   wire n_1_737_2647;
   wire n_1_737_2648;
   wire n_1_737_2649;
   wire n_1_737_2650;
   wire n_1_737_2651;
   wire n_1_737_2652;
   wire n_1_737_2653;
   wire n_1_737_2654;
   wire n_1_737_2655;
   wire n_1_737_2656;
   wire n_1_737_2657;
   wire n_1_737_2658;
   wire n_1_737_2659;
   wire n_1_737_2660;
   wire n_1_737_2661;
   wire n_1_737_2662;
   wire n_1_737_2663;
   wire n_1_737_2664;
   wire n_1_737_2665;
   wire n_1_737_2666;
   wire n_1_737_2667;
   wire n_1_737_2668;
   wire n_1_737_2669;
   wire n_1_737_2670;
   wire n_1_737_2671;
   wire n_1_737_2672;
   wire n_1_737_2673;
   wire n_1_737_2674;
   wire n_1_737_2675;
   wire n_1_737_2676;
   wire n_1_737_2677;
   wire n_1_737_2678;
   wire n_1_737_2679;
   wire n_1_737_2680;
   wire n_1_737_2681;
   wire n_1_737_2682;
   wire n_1_737_2683;
   wire n_1_737_2684;
   wire n_1_737_2685;
   wire n_1_737_2686;
   wire n_1_737_2687;
   wire n_1_737_2688;
   wire n_1_737_2689;
   wire n_1_737_2690;
   wire n_1_737_2691;
   wire n_1_737_2692;
   wire n_1_737_2693;
   wire n_1_737_2694;
   wire n_1_737_2695;
   wire n_1_737_2696;
   wire n_1_737_2697;
   wire n_1_737_2698;
   wire n_1_737_2699;
   wire n_1_737_2700;
   wire n_1_737_2701;
   wire n_1_737_2702;
   wire n_1_737_2703;
   wire n_1_737_2704;
   wire n_1_737_2705;
   wire n_1_737_2706;
   wire n_1_737_2707;
   wire n_1_737_2708;
   wire n_1_737_2709;
   wire n_1_737_2710;
   wire n_1_737_2711;
   wire n_1_737_2712;
   wire n_1_737_2713;
   wire n_1_737_2714;
   wire n_1_737_2715;
   wire n_1_737_2716;
   wire n_1_737_2717;
   wire n_1_737_2718;
   wire n_1_737_2719;
   wire n_1_737_2720;
   wire n_1_737_2721;
   wire n_1_737_2722;
   wire n_1_737_2723;
   wire n_1_737_2724;
   wire n_1_737_2725;
   wire n_1_737_2726;
   wire n_1_737_2727;
   wire n_1_737_2728;
   wire n_1_737_2729;
   wire n_1_737_2730;
   wire n_1_737_2731;
   wire n_1_737_2732;
   wire n_1_737_2733;
   wire n_1_737_2734;
   wire n_1_737_2735;
   wire n_1_737_2736;
   wire n_1_737_2737;
   wire n_1_737_2738;
   wire n_1_737_2739;
   wire n_1_737_2740;
   wire n_1_737_2741;
   wire n_1_737_2742;
   wire n_1_737_2743;
   wire n_1_737_2744;
   wire n_1_737_2745;
   wire n_1_737_2746;
   wire n_1_737_2747;
   wire n_1_737_2748;
   wire n_1_737_2749;
   wire n_1_737_2750;
   wire n_1_737_2751;
   wire n_1_737_2752;
   wire n_1_737_2753;
   wire n_1_737_2754;
   wire n_1_737_2755;
   wire n_1_737_2756;
   wire n_1_737_2757;
   wire n_1_737_2758;
   wire n_1_737_2759;
   wire n_1_737_2760;
   wire n_1_737_2761;
   wire n_1_737_2762;
   wire n_1_737_2763;
   wire n_1_737_2764;
   wire n_1_737_2765;
   wire n_1_737_2766;
   wire n_1_737_2767;
   wire n_1_737_2768;
   wire n_1_737_2769;
   wire n_1_737_2770;
   wire n_1_737_2771;
   wire n_1_737_2772;
   wire n_1_737_2773;
   wire n_1_737_2774;
   wire n_1_737_2775;
   wire n_1_737_2776;
   wire n_1_737_2777;
   wire n_1_737_2778;
   wire n_1_737_2779;
   wire n_1_737_2780;
   wire n_1_737_2781;
   wire n_1_737_2782;
   wire n_1_737_2783;
   wire n_1_737_2784;
   wire n_1_737_2785;
   wire n_1_737_2786;
   wire n_1_737_2787;
   wire n_1_737_2788;
   wire n_1_737_2789;
   wire n_1_737_2790;
   wire n_1_737_2791;
   wire n_1_737_2792;
   wire n_1_737_2793;
   wire n_1_737_2794;
   wire n_1_737_2795;
   wire n_1_737_2796;
   wire n_1_737_2797;
   wire n_1_737_2798;
   wire n_1_737_2799;
   wire n_1_737_2800;
   wire n_1_737_2801;
   wire n_1_737_2802;
   wire n_1_737_2803;
   wire n_1_737_2804;
   wire n_1_737_2805;
   wire n_1_737_2806;
   wire n_1_737_2807;
   wire n_1_737_2808;
   wire n_1_737_2809;
   wire n_1_737_2810;
   wire n_1_737_2811;
   wire n_1_737_2812;
   wire n_1_737_2813;
   wire n_1_737_2814;
   wire n_1_737_2815;
   wire n_1_737_2816;
   wire n_1_737_2817;
   wire n_1_737_2818;
   wire n_1_737_2819;
   wire n_1_737_2820;
   wire n_1_737_2821;
   wire n_1_737_2822;
   wire n_1_737_2823;
   wire n_1_737_2824;
   wire n_1_737_2825;
   wire n_1_737_2826;
   wire n_1_737_2827;
   wire n_1_737_2828;
   wire n_1_737_2829;
   wire n_1_737_2830;
   wire n_1_737_2831;
   wire n_1_737_2832;
   wire n_1_737_2833;
   wire n_1_737_2834;
   wire n_1_737_2835;
   wire n_1_737_2836;
   wire n_1_737_2837;
   wire n_1_737_2838;
   wire n_1_737_2839;
   wire n_1_737_2840;
   wire n_1_737_2841;
   wire n_1_737_2842;
   wire n_1_737_2843;
   wire n_1_737_2844;
   wire n_1_737_2845;
   wire n_1_737_2846;
   wire n_1_737_2847;
   wire n_1_737_2848;
   wire n_1_737_2849;
   wire n_1_737_2850;
   wire n_1_737_2851;
   wire n_1_737_2852;
   wire n_1_737_2853;
   wire n_1_737_2854;
   wire n_1_737_2855;
   wire n_1_737_2856;
   wire n_1_737_2857;
   wire n_1_737_2858;
   wire n_1_737_2859;
   wire n_1_737_2860;
   wire n_1_737_2861;
   wire n_1_737_2862;
   wire n_1_737_2863;
   wire n_1_737_2864;
   wire n_1_737_2865;
   wire n_1_737_2866;
   wire n_1_737_2867;
   wire n_1_737_2868;
   wire n_1_737_2869;
   wire n_1_737_2870;
   wire n_1_737_2871;
   wire n_1_737_2872;
   wire n_1_737_2873;
   wire n_1_737_2874;
   wire n_1_737_2875;
   wire n_1_737_2876;
   wire n_1_737_2877;
   wire n_1_737_2878;
   wire n_1_737_2879;
   wire n_1_737_2880;
   wire n_1_737_2881;
   wire n_1_737_2882;
   wire n_1_737_2883;
   wire n_1_737_2884;
   wire n_1_737_2885;
   wire n_1_737_2886;
   wire n_1_737_2887;
   wire n_1_737_2888;
   wire n_1_737_2889;
   wire n_1_737_2890;
   wire n_1_737_2891;
   wire n_1_737_2892;
   wire n_1_737_2893;
   wire n_1_737_2894;
   wire n_1_737_2895;
   wire n_1_737_2896;
   wire n_1_737_2897;
   wire n_1_737_2898;
   wire n_1_737_2899;
   wire n_1_737_2900;
   wire n_1_737_2901;
   wire n_1_737_2902;
   wire n_1_737_2903;
   wire n_1_737_2904;
   wire n_1_737_2905;
   wire n_1_737_2906;
   wire n_1_737_2907;
   wire n_1_737_2908;
   wire n_1_737_2909;
   wire n_1_737_2910;
   wire n_1_737_2911;
   wire n_1_737_2912;
   wire n_1_737_2913;
   wire n_1_737_2914;
   wire n_1_737_2915;
   wire n_1_737_2916;
   wire n_1_737_2917;
   wire n_1_737_2918;
   wire n_1_737_2919;
   wire n_1_737_2920;
   wire n_1_737_2921;
   wire n_1_737_2922;
   wire n_1_737_2923;
   wire n_1_737_2924;
   wire n_1_737_2925;
   wire n_1_737_2926;
   wire n_1_737_2927;
   wire n_1_737_2928;
   wire n_1_737_2929;
   wire n_1_737_2930;
   wire n_1_737_2931;
   wire n_1_737_2932;
   wire n_1_737_2933;
   wire n_1_737_2934;
   wire n_1_737_2935;
   wire n_1_737_2936;
   wire n_1_737_2937;
   wire n_1_737_2938;
   wire n_1_737_2939;
   wire n_1_737_2940;
   wire n_1_737_2941;
   wire n_1_737_2942;
   wire n_1_737_2943;
   wire n_1_737_2944;
   wire n_1_737_2945;
   wire n_1_737_2946;
   wire n_1_737_2947;
   wire n_1_737_2948;
   wire n_1_737_2949;
   wire n_1_737_2950;
   wire n_1_737_2951;
   wire n_1_737_2952;
   wire n_1_737_2953;
   wire n_1_737_2954;
   wire n_1_737_2955;
   wire n_1_737_2956;
   wire n_1_737_2957;
   wire n_1_737_2958;
   wire n_1_737_2959;
   wire n_1_737_2960;
   wire n_1_737_2961;
   wire n_1_737_2962;
   wire n_1_737_2963;
   wire n_1_737_2964;
   wire n_1_737_2965;
   wire n_1_737_2966;
   wire n_1_737_2967;
   wire n_1_737_2968;
   wire n_1_737_2969;
   wire n_1_737_2970;
   wire n_1_737_2971;
   wire n_1_737_2972;
   wire n_1_737_2973;
   wire n_1_737_2974;
   wire n_1_737_2975;
   wire n_1_737_2976;
   wire n_1_737_2977;
   wire n_1_737_2978;
   wire n_1_737_2979;
   wire n_1_737_2980;
   wire n_1_737_2981;
   wire n_1_737_2982;
   wire n_1_737_2983;
   wire n_1_737_2984;
   wire n_1_737_2985;
   wire n_1_737_2986;
   wire n_1_737_2987;
   wire n_1_737_2988;
   wire n_1_737_2989;
   wire n_1_737_2990;
   wire n_1_737_2991;
   wire n_1_737_2992;
   wire n_1_737_2993;
   wire n_1_737_2994;
   wire n_1_737_2995;
   wire n_1_737_2996;
   wire n_1_737_2997;
   wire n_1_737_2998;
   wire n_1_737_2999;
   wire n_1_737_3000;
   wire n_1_737_3001;
   wire n_1_737_3002;
   wire n_1_737_3003;
   wire n_1_737_3004;
   wire n_1_737_3005;
   wire n_1_737_3006;
   wire n_1_737_3007;
   wire n_1_737_3008;
   wire n_1_737_3009;
   wire n_1_737_3010;
   wire n_1_737_3011;
   wire n_1_737_3012;
   wire n_1_737_3013;
   wire n_1_737_3014;
   wire n_1_737_3015;
   wire n_1_737_3016;
   wire n_1_737_3017;
   wire n_1_737_3018;
   wire n_1_737_3019;
   wire n_1_737_3020;
   wire n_1_737_3021;
   wire n_1_737_3022;
   wire n_1_737_3023;
   wire n_1_737_3024;
   wire n_1_737_3025;
   wire n_1_737_3026;
   wire n_1_737_3027;
   wire n_1_737_3028;
   wire n_1_737_3029;
   wire n_1_737_3030;
   wire n_1_737_3031;
   wire n_1_737_3032;
   wire n_1_737_3033;
   wire n_1_737_3034;
   wire n_1_737_3035;
   wire n_1_737_3036;
   wire n_1_737_3037;
   wire n_1_737_3038;
   wire n_1_737_3039;
   wire n_1_737_3040;
   wire n_1_737_3041;
   wire n_1_737_3042;
   wire n_1_737_3043;
   wire n_1_737_3044;
   wire n_1_737_3045;
   wire n_1_737_3046;
   wire n_1_737_3047;
   wire n_1_737_3048;
   wire n_1_737_3049;
   wire n_1_737_3050;
   wire n_1_737_3051;
   wire n_1_737_3052;
   wire n_1_737_3053;
   wire n_1_737_3054;
   wire n_1_737_3055;
   wire n_1_737_3056;
   wire n_1_737_3057;
   wire n_1_737_3058;
   wire n_1_737_3059;
   wire n_1_737_3060;
   wire n_1_737_3061;
   wire n_1_737_3062;
   wire n_1_737_3063;
   wire n_1_737_3064;
   wire n_1_737_3065;
   wire n_1_737_3066;
   wire n_1_737_3067;
   wire n_1_737_3068;
   wire n_1_737_3069;
   wire n_1_737_3070;
   wire n_1_737_3071;
   wire n_1_737_3072;
   wire n_1_737_3073;
   wire n_1_737_3074;
   wire n_1_737_3075;
   wire n_1_737_3076;
   wire n_1_737_3077;
   wire n_1_737_3078;
   wire n_1_737_3079;
   wire n_1_737_3080;
   wire n_1_737_3081;
   wire n_1_737_3082;
   wire n_1_737_3083;
   wire n_1_737_3084;
   wire n_1_737_3085;
   wire n_1_737_3086;
   wire n_1_737_3087;
   wire n_1_737_3088;
   wire n_1_737_3089;
   wire n_1_737_3090;
   wire n_1_737_3091;
   wire n_1_737_3092;
   wire n_1_737_3093;
   wire n_1_737_3094;
   wire n_1_737_3095;
   wire n_1_737_3096;
   wire n_1_737_3097;
   wire n_1_737_3098;
   wire n_1_737_3099;
   wire n_1_737_3100;
   wire n_1_737_3101;
   wire n_1_737_3102;
   wire n_1_737_3103;
   wire n_1_737_3104;
   wire n_1_737_3105;
   wire n_1_737_3106;
   wire n_1_737_3107;
   wire n_1_737_3108;
   wire n_1_737_3109;
   wire n_1_737_3111;
   wire n_1_737_3112;
   wire n_1_737_3113;
   wire n_1_737_3114;
   wire n_1_737_3115;
   wire n_1_737_3116;
   wire n_1_737_3117;
   wire n_1_737_3118;
   wire n_1_737_3119;
   wire n_1_737_3120;
   wire n_1_737_3121;
   wire n_1_737_3122;
   wire n_1_737_3123;
   wire n_1_737_3124;
   wire n_1_737_3125;
   wire n_1_737_3126;
   wire n_1_737_3127;
   wire n_1_737_3128;
   wire n_1_737_3129;
   wire n_1_737_3130;
   wire n_1_737_3131;
   wire n_1_737_3132;
   wire n_1_737_3133;
   wire n_1_737_3134;
   wire n_1_737_3135;
   wire n_1_737_3136;
   wire n_1_737_3137;
   wire n_1_737_3138;
   wire n_1_737_3139;
   wire n_1_737_3140;
   wire n_1_737_3141;
   wire n_1_737_3142;
   wire n_1_737_3143;
   wire n_1_737_3144;
   wire n_1_737_3145;
   wire n_1_737_3146;
   wire n_1_737_3147;
   wire n_1_737_3148;
   wire n_1_737_3149;
   wire n_1_737_3150;
   wire n_1_737_3151;
   wire n_1_737_3152;
   wire n_1_737_3153;
   wire n_1_737_3154;
   wire n_1_737_3155;
   wire n_1_737_3156;
   wire n_1_737_3157;
   wire n_1_737_3158;
   wire n_1_737_3159;
   wire n_1_737_3160;
   wire n_1_737_3161;
   wire n_1_737_3162;
   wire n_1_737_3163;
   wire n_1_737_3164;
   wire n_1_737_3165;
   wire n_1_737_3166;
   wire n_1_737_3167;
   wire n_1_737_3168;
   wire n_1_737_3169;
   wire n_1_737_3170;
   wire n_1_737_3171;
   wire n_1_737_3172;
   wire n_1_737_3173;
   wire n_1_737_3174;
   wire n_1_737_3175;
   wire n_1_737_3176;
   wire n_1_737_3177;
   wire n_1_737_3178;
   wire n_1_737_3179;
   wire n_1_737_3180;
   wire n_1_737_3181;
   wire n_1_737_3182;
   wire n_1_737_3183;
   wire n_1_737_3184;
   wire n_1_737_3185;
   wire n_1_737_3186;
   wire n_1_737_3187;
   wire n_1_737_3188;
   wire n_1_737_3189;
   wire n_1_737_3190;
   wire n_1_737_3191;
   wire n_1_737_3192;
   wire n_1_737_3193;
   wire n_1_737_3194;
   wire n_1_737_3195;
   wire n_1_737_3196;
   wire n_1_737_3197;
   wire n_1_737_3198;
   wire n_1_737_3199;
   wire n_1_737_3200;
   wire n_1_737_3201;
   wire n_1_737_3202;
   wire n_1_737_3203;
   wire n_1_737_3204;
   wire n_1_737_3205;
   wire n_1_737_3206;
   wire n_1_737_3207;
   wire n_1_737_3208;
   wire n_1_737_3209;
   wire n_1_737_3210;
   wire n_1_737_3211;
   wire n_1_737_3212;
   wire n_1_737_3213;
   wire n_1_737_3214;
   wire n_1_737_3215;
   wire n_1_737_3216;
   wire n_1_737_3217;
   wire n_1_737_3218;
   wire n_1_737_3219;
   wire n_1_737_3220;
   wire n_1_737_3221;
   wire n_1_737_3222;
   wire n_1_737_3223;
   wire n_1_737_3224;
   wire n_1_737_3225;
   wire n_1_737_3226;
   wire n_1_737_3227;
   wire n_1_737_3228;
   wire n_1_737_3229;
   wire n_1_737_3230;
   wire n_1_737_3231;
   wire n_1_737_3232;
   wire n_1_737_3233;
   wire n_1_737_3234;
   wire n_1_737_3235;
   wire n_1_737_3236;
   wire n_1_737_3237;
   wire n_1_737_3238;
   wire n_1_737_3239;
   wire n_1_737_3240;
   wire n_1_737_3241;
   wire n_1_737_3242;
   wire n_1_737_3243;
   wire n_1_737_3244;
   wire n_1_737_3245;
   wire n_1_737_3246;
   wire n_1_737_3247;
   wire n_1_737_3248;
   wire n_1_737_3249;
   wire n_1_737_3250;
   wire n_1_737_3251;
   wire n_1_737_3252;
   wire n_1_737_3253;
   wire n_1_737_3254;
   wire n_1_737_3255;
   wire n_1_737_3256;
   wire n_1_737_3257;
   wire n_1_737_3258;
   wire n_1_737_3259;
   wire n_1_737_3260;
   wire n_1_737_3261;
   wire n_1_737_3262;
   wire n_1_737_3263;
   wire n_1_737_3264;
   wire n_1_737_3265;
   wire n_1_737_3266;
   wire n_1_737_3267;
   wire n_1_737_3268;
   wire n_1_737_3269;
   wire n_1_737_3270;
   wire n_1_737_3271;
   wire n_1_737_3272;
   wire n_1_737_3273;
   wire n_1_737_3274;
   wire n_1_737_3275;
   wire n_1_737_3276;
   wire n_1_737_3277;
   wire n_1_737_3278;
   wire n_1_737_3279;
   wire n_1_737_3280;
   wire n_1_737_3281;
   wire n_1_737_3282;
   wire n_1_737_3283;
   wire n_1_737_3284;
   wire n_1_737_3285;
   wire n_1_737_3286;
   wire n_1_737_3287;
   wire n_1_737_3288;
   wire n_1_737_3289;
   wire n_1_737_3290;
   wire n_1_737_3291;
   wire n_1_737_3292;
   wire n_1_737_3293;
   wire n_1_737_3294;
   wire n_1_737_3295;
   wire n_1_737_3296;
   wire n_1_737_3297;
   wire n_1_737_3298;
   wire n_1_737_3299;
   wire n_1_737_3300;
   wire n_1_737_3301;
   wire n_1_737_3302;
   wire n_1_737_3303;
   wire n_1_737_3304;
   wire n_1_737_3305;
   wire n_1_737_3306;
   wire n_1_737_3307;
   wire n_1_737_3308;
   wire n_1_737_3309;
   wire n_1_737_3310;
   wire n_1_737_3311;
   wire n_1_737_3312;
   wire n_1_737_3313;
   wire n_1_737_3314;
   wire n_1_737_3315;
   wire n_1_737_3316;
   wire n_1_737_3317;
   wire n_1_737_3318;
   wire n_1_737_3319;
   wire n_1_737_3320;
   wire n_1_737_3321;
   wire n_1_737_3322;
   wire n_1_737_3323;
   wire n_1_737_3324;
   wire n_1_737_3325;
   wire n_1_737_3326;
   wire n_1_737_3327;
   wire n_1_737_3328;
   wire n_1_737_3329;
   wire n_1_737_3330;
   wire n_1_737_3331;
   wire n_1_737_3332;
   wire n_1_737_3333;
   wire n_1_737_3334;
   wire n_1_737_3335;
   wire n_1_737_3336;
   wire n_1_737_3337;
   wire n_1_737_3338;
   wire n_1_737_3339;
   wire n_1_737_3340;
   wire n_1_737_3341;
   wire n_1_737_3342;
   wire n_1_737_3343;
   wire n_1_737_3344;
   wire n_1_737_3345;
   wire n_1_737_3346;
   wire n_1_737_3347;
   wire n_1_737_3348;
   wire n_1_737_3349;
   wire n_1_737_3350;
   wire n_1_737_3351;
   wire n_1_737_3352;
   wire n_1_737_3353;
   wire n_1_737_3354;
   wire n_1_737_3355;
   wire n_1_737_3356;
   wire n_1_737_3357;
   wire n_1_737_3358;
   wire n_1_737_3359;
   wire n_1_737_3360;
   wire n_1_737_3361;
   wire n_1_737_3362;
   wire n_1_737_3363;
   wire n_1_737_3364;
   wire n_1_737_3365;
   wire n_1_737_3366;
   wire n_1_737_3367;
   wire n_1_737_3368;
   wire n_1_737_3369;
   wire n_1_737_3370;
   wire n_1_737_3371;
   wire n_1_737_3372;
   wire n_1_737_3373;
   wire n_1_737_3374;
   wire n_1_737_3375;
   wire n_1_737_3376;
   wire n_1_737_3377;
   wire n_1_737_3378;
   wire n_1_737_3379;
   wire n_1_737_3380;
   wire n_1_737_3381;
   wire n_1_737_3382;
   wire n_1_737_3383;
   wire n_1_737_3384;
   wire n_1_737_3385;
   wire n_1_737_3386;
   wire n_1_737_3387;
   wire n_1_737_3388;
   wire n_1_737_3389;
   wire n_1_737_3390;
   wire n_1_737_3391;
   wire n_1_737_3392;
   wire n_1_737_3393;
   wire n_1_737_3394;
   wire n_1_737_3395;
   wire n_1_737_3396;
   wire n_1_737_3397;
   wire n_1_737_3398;
   wire n_1_737_3399;
   wire n_1_737_3400;
   wire n_1_737_3401;
   wire n_1_737_3402;
   wire n_1_737_3403;
   wire n_1_737_3404;
   wire n_1_737_3405;
   wire n_1_737_3406;
   wire n_1_737_3407;
   wire n_1_737_3408;
   wire n_1_737_3409;
   wire n_1_737_3410;
   wire n_1_737_3411;
   wire n_1_737_3412;
   wire n_1_737_3413;
   wire n_1_737_3414;
   wire n_1_737_3415;
   wire n_1_737_3416;
   wire n_1_737_3417;
   wire n_1_737_3418;
   wire n_1_737_3419;
   wire n_1_737_3420;
   wire n_1_737_3421;
   wire n_1_737_3422;
   wire n_1_737_3423;
   wire n_1_737_3424;
   wire n_1_737_3425;
   wire n_1_737_3426;
   wire n_1_737_3427;
   wire n_1_737_3428;
   wire n_1_737_3429;
   wire n_1_737_3430;
   wire n_1_737_3431;
   wire n_1_737_3432;
   wire n_1_737_3433;
   wire n_1_737_3434;
   wire n_1_737_3435;
   wire n_1_737_3436;
   wire n_1_737_3437;
   wire n_1_737_3438;
   wire n_1_737_3439;
   wire n_1_737_3440;
   wire n_1_737_3441;
   wire n_1_737_3442;
   wire n_1_737_3443;
   wire n_1_737_3444;
   wire n_1_737_3445;
   wire n_1_737_3446;
   wire n_1_737_3447;
   wire n_1_737_3448;
   wire n_1_737_3449;
   wire n_1_737_3450;
   wire n_1_737_3451;
   wire n_1_737_3452;
   wire n_1_737_3453;
   wire n_1_737_3454;
   wire n_1_737_3455;
   wire n_1_737_3456;
   wire n_1_737_3457;
   wire n_1_737_3458;
   wire n_1_737_3459;
   wire n_1_737_3460;
   wire n_1_737_3461;
   wire n_1_737_3462;
   wire n_1_737_3463;
   wire n_1_737_3464;
   wire n_1_737_3465;
   wire n_1_737_3466;
   wire n_1_737_3467;
   wire n_1_737_3468;
   wire n_1_737_3469;
   wire n_1_737_3470;
   wire n_1_737_3471;
   wire n_1_737_3472;
   wire n_1_737_3473;
   wire n_1_737_3474;
   wire n_1_737_3475;
   wire n_1_737_3476;
   wire n_1_737_3477;
   wire n_1_737_3478;
   wire n_1_737_3479;
   wire n_1_737_3480;
   wire n_1_737_3481;
   wire n_1_737_3482;
   wire n_1_737_3483;
   wire n_1_737_3484;
   wire n_1_737_3485;
   wire n_1_737_3486;
   wire n_1_737_3487;
   wire n_1_737_3488;
   wire n_1_737_3489;
   wire n_1_737_3490;
   wire n_1_737_3491;
   wire n_1_737_3492;
   wire n_1_737_3493;
   wire n_1_737_3494;
   wire n_1_737_3495;
   wire n_1_737_3496;
   wire n_1_737_3497;
   wire n_1_737_3498;
   wire n_1_737_3499;
   wire n_1_737_3500;
   wire n_1_737_3501;
   wire n_1_737_3502;
   wire n_1_737_3503;
   wire n_1_737_3504;
   wire n_1_737_3505;
   wire n_1_737_3506;
   wire n_1_737_3507;
   wire n_1_737_3508;
   wire n_1_737_3509;
   wire n_1_737_3510;
   wire n_1_737_3511;
   wire n_1_737_3512;
   wire n_1_737_3513;
   wire n_1_737_3514;
   wire n_1_737_3515;
   wire n_1_737_3516;
   wire n_1_737_3517;
   wire n_1_737_3518;
   wire n_1_737_3519;
   wire n_1_737_3520;
   wire n_1_737_3521;
   wire n_1_737_3522;
   wire n_1_737_3523;
   wire n_1_737_3524;
   wire n_1_737_3525;
   wire n_1_737_3526;
   wire n_1_737_3527;
   wire n_1_737_3528;
   wire n_1_737_3529;
   wire n_1_737_3530;
   wire n_1_737_3531;
   wire n_1_737_3532;
   wire n_1_737_3533;
   wire n_1_737_3534;
   wire n_1_737_3535;
   wire n_1_737_3536;
   wire n_1_737_3537;
   wire n_1_737_3538;
   wire n_1_737_3539;
   wire n_1_737_3540;
   wire n_1_737_3541;
   wire n_1_737_3542;
   wire n_1_737_3543;
   wire n_1_737_3544;
   wire n_1_737_3545;
   wire n_1_737_3546;
   wire n_1_737_3547;
   wire n_1_737_3548;
   wire n_1_737_3549;
   wire n_1_737_3550;
   wire n_1_737_3551;
   wire n_1_737_3552;
   wire n_1_737_3553;
   wire n_1_737_3554;
   wire n_1_737_3555;
   wire n_1_737_3556;
   wire n_1_737_3557;
   wire n_1_737_3558;
   wire n_1_737_3559;
   wire n_1_737_3560;
   wire n_1_737_3561;
   wire n_1_737_3562;
   wire n_1_737_3563;
   wire n_1_737_3564;
   wire n_1_737_3565;
   wire n_1_737_3566;
   wire n_1_737_3567;
   wire n_1_737_3568;
   wire n_1_737_3569;
   wire n_1_737_3570;
   wire n_1_737_3571;
   wire n_1_737_3572;
   wire n_1_737_3573;
   wire n_1_737_3574;
   wire n_1_737_3575;
   wire n_1_737_3576;
   wire n_1_737_3577;
   wire n_1_737_3578;
   wire n_1_737_3579;
   wire n_1_737_3580;
   wire n_1_737_3581;
   wire n_1_737_3582;
   wire n_1_737_3583;
   wire n_1_737_3584;
   wire n_1_737_3585;
   wire n_1_737_3586;
   wire n_1_737_3587;
   wire n_1_737_3588;
   wire n_1_737_3589;
   wire n_1_737_3590;
   wire n_1_737_3591;
   wire n_1_737_3592;
   wire n_1_737_3593;
   wire n_1_737_3594;
   wire n_1_737_3595;
   wire n_1_737_3596;
   wire n_1_737_3597;
   wire n_1_737_3598;
   wire n_1_737_3599;
   wire n_1_737_3600;
   wire n_1_737_3601;
   wire n_1_737_3602;
   wire n_1_737_3603;
   wire n_1_737_3604;
   wire n_1_737_3605;
   wire n_1_737_3606;
   wire n_1_737_3607;
   wire n_1_737_3608;
   wire n_1_737_3609;
   wire n_1_737_3610;
   wire n_1_737_3611;
   wire n_1_737_3612;
   wire n_1_737_3613;
   wire n_1_737_3614;
   wire n_1_737_3615;
   wire n_1_737_3616;
   wire n_1_737_3617;
   wire n_1_737_3618;
   wire n_1_737_3619;
   wire n_1_737_3620;
   wire n_1_737_3621;
   wire n_1_737_3622;
   wire n_1_737_3623;
   wire n_1_737_3624;
   wire n_1_737_3625;
   wire n_1_737_3626;
   wire n_1_737_3627;
   wire n_1_737_3628;
   wire n_1_737_3629;
   wire n_1_737_3630;
   wire n_1_737_3631;
   wire n_1_737_3632;
   wire n_1_737_3633;
   wire n_1_737_3634;
   wire n_1_737_3635;
   wire n_1_737_3636;
   wire n_1_737_3637;
   wire n_1_737_3638;
   wire n_1_737_3639;
   wire n_1_737_3640;
   wire n_1_737_3641;
   wire n_1_737_3642;
   wire n_1_737_3643;
   wire n_1_737_3644;
   wire n_1_737_3645;
   wire n_1_737_3646;
   wire n_1_737_3647;
   wire n_1_737_3648;
   wire n_1_737_3649;
   wire n_1_737_3650;
   wire n_1_737_3651;
   wire n_1_737_3652;
   wire n_1_737_3653;
   wire n_1_737_3654;
   wire n_1_737_3655;
   wire n_1_737_3656;
   wire n_1_737_3657;
   wire n_1_737_3658;
   wire n_1_737_3659;
   wire n_1_737_3660;
   wire n_1_737_3661;
   wire n_1_737_3662;
   wire n_1_737_3663;
   wire n_1_737_3664;
   wire n_1_737_3665;
   wire n_1_737_3666;
   wire n_1_737_3667;
   wire n_1_737_3668;
   wire n_1_737_3669;
   wire n_1_737_3670;
   wire n_1_737_3671;
   wire n_1_737_3672;
   wire n_1_737_3673;
   wire n_1_737_3674;
   wire n_1_737_3675;
   wire n_1_737_3676;
   wire n_1_737_3677;
   wire n_1_737_3678;
   wire n_1_737_3679;
   wire n_1_737_3680;
   wire n_1_737_3681;
   wire n_1_737_3682;
   wire n_1_737_3683;
   wire n_1_737_3684;
   wire n_1_737_3685;
   wire n_1_737_3686;
   wire n_1_737_3687;
   wire n_1_737_3688;
   wire n_1_737_3689;
   wire n_1_737_3690;
   wire n_1_737_3691;
   wire n_1_737_3692;
   wire n_1_737_3693;
   wire n_1_737_3694;
   wire n_1_737_3695;
   wire n_1_737_3696;
   wire n_1_737_3697;
   wire n_1_737_3698;
   wire n_1_737_3699;
   wire n_1_737_3700;
   wire n_1_737_3701;
   wire n_1_737_3702;
   wire n_1_737_3703;
   wire n_1_737_3704;
   wire n_1_737_3705;
   wire n_1_737_3706;
   wire n_1_737_3707;
   wire n_1_737_3708;
   wire n_1_737_3709;
   wire n_1_737_3710;
   wire n_1_737_3711;
   wire n_1_737_3712;
   wire n_1_737_3713;
   wire n_1_737_3714;
   wire n_1_737_3715;
   wire n_1_737_3716;
   wire n_1_737_3717;
   wire n_1_737_3718;
   wire n_1_737_3719;
   wire n_1_737_3720;
   wire n_1_737_3721;
   wire n_1_737_3722;
   wire n_1_737_3723;
   wire n_1_737_3724;
   wire n_1_737_3725;
   wire n_1_737_3726;
   wire n_1_737_3727;
   wire n_1_737_3728;
   wire n_1_737_3729;
   wire n_1_737_3730;
   wire n_1_737_3731;
   wire n_1_737_3732;
   wire n_1_737_3733;
   wire n_1_737_3734;
   wire n_1_737_3735;
   wire n_1_737_3736;
   wire n_1_737_3737;
   wire n_1_737_3738;
   wire n_1_737_3739;
   wire n_1_737_3740;
   wire n_1_737_3741;
   wire n_1_737_3742;
   wire n_1_737_3743;
   wire n_1_737_3744;
   wire n_1_737_3745;
   wire n_1_737_3746;
   wire n_1_737_3747;
   wire n_1_737_3748;
   wire n_1_737_3749;
   wire n_1_737_3750;
   wire n_1_737_3751;
   wire n_1_737_3752;
   wire n_1_737_3753;
   wire n_1_737_3754;
   wire n_1_737_3755;
   wire n_1_737_3756;
   wire n_1_737_3757;
   wire n_1_737_3758;
   wire n_1_737_3759;
   wire n_1_737_3760;
   wire n_1_737_3761;
   wire n_1_737_3762;
   wire n_1_737_3763;
   wire n_1_737_3764;
   wire n_1_737_3765;
   wire n_1_737_3766;
   wire n_1_737_3767;
   wire n_1_737_3768;
   wire n_1_737_3769;
   wire n_1_737_3770;
   wire n_1_737_3771;
   wire n_1_737_3772;
   wire n_1_737_3773;
   wire n_1_737_3774;
   wire n_1_737_3775;
   wire n_1_737_3776;
   wire n_1_737_3777;
   wire n_1_737_3778;
   wire n_1_737_3779;
   wire n_1_737_3780;
   wire n_1_737_3781;
   wire n_1_737_3782;
   wire n_1_737_3783;
   wire n_1_737_3784;
   wire n_1_737_3785;
   wire n_1_737_3786;
   wire n_1_737_3787;
   wire n_1_737_3788;
   wire n_1_737_3789;
   wire n_1_737_3790;
   wire n_1_737_3791;
   wire n_1_737_3792;
   wire n_1_737_3793;
   wire n_1_737_3794;
   wire n_1_737_3795;
   wire n_1_737_3796;
   wire n_1_737_3797;
   wire n_1_737_3798;
   wire n_1_737_3799;
   wire n_1_737_3800;
   wire n_1_737_3801;
   wire n_1_737_3802;
   wire n_1_737_3803;
   wire n_1_737_3804;
   wire n_1_737_3805;
   wire n_1_737_3806;
   wire n_1_737_3807;
   wire n_1_737_3808;
   wire n_1_737_3809;
   wire n_1_737_3810;
   wire n_1_737_3811;
   wire n_1_737_3812;
   wire n_1_737_3813;
   wire n_1_737_3814;
   wire n_1_737_3815;
   wire n_1_737_3816;
   wire n_1_737_3817;
   wire n_1_737_3818;
   wire n_1_737_3819;
   wire n_1_737_3820;
   wire n_1_737_3821;
   wire n_1_737_3822;
   wire n_1_737_3823;
   wire n_1_737_3824;
   wire n_1_737_3825;
   wire n_1_737_3826;
   wire n_1_737_3827;
   wire n_1_737_3828;
   wire n_1_737_3829;
   wire n_1_737_3830;
   wire n_1_737_3831;
   wire n_1_737_3832;
   wire n_1_737_3833;
   wire n_1_737_3834;
   wire n_1_737_3835;
   wire n_1_737_3836;
   wire n_1_737_3837;
   wire n_1_737_3838;
   wire n_1_737_3839;
   wire n_1_737_3840;
   wire n_1_737_3841;
   wire n_1_737_3842;
   wire n_1_737_3843;
   wire n_1_737_3844;
   wire n_1_737_3845;
   wire n_1_737_3846;
   wire n_1_737_3847;
   wire n_1_737_3848;
   wire n_1_737_3849;
   wire n_1_737_3850;
   wire n_1_737_3851;
   wire n_1_737_3852;
   wire n_1_737_3853;
   wire n_1_737_3854;
   wire n_1_737_3855;
   wire n_1_737_3856;
   wire n_1_737_3857;
   wire n_1_737_3858;
   wire n_1_737_3859;
   wire n_1_737_3860;
   wire n_1_737_3861;
   wire n_1_737_3862;
   wire n_1_737_3863;
   wire n_1_737_3864;
   wire n_1_737_3865;
   wire n_1_737_3866;
   wire n_1_737_3867;
   wire n_1_737_3868;
   wire n_1_737_3869;
   wire n_1_737_3870;
   wire n_1_737_3871;
   wire n_1_737_3872;
   wire n_1_737_3873;
   wire n_1_737_3874;
   wire n_1_737_3875;
   wire n_1_737_3876;
   wire n_1_737_3877;
   wire n_1_737_3878;
   wire n_1_737_3879;
   wire n_1_737_3880;
   wire n_1_737_3881;
   wire n_1_737_3882;
   wire n_1_737_3883;
   wire n_1_737_3884;
   wire n_1_737_3885;
   wire n_1_737_3886;
   wire n_1_737_3887;
   wire n_1_737_3888;
   wire n_1_737_3889;
   wire n_1_737_3890;
   wire n_1_737_3891;
   wire n_1_737_3892;
   wire n_1_737_3893;
   wire n_1_737_3894;
   wire n_1_737_3895;
   wire n_1_737_3896;
   wire n_1_737_3897;
   wire n_1_737_3898;
   wire n_1_737_3899;
   wire n_1_737_3900;
   wire n_1_737_3901;
   wire n_1_737_3902;
   wire n_1_737_3903;
   wire n_1_737_3904;
   wire n_1_737_3905;
   wire n_1_737_3906;
   wire n_1_737_3907;
   wire n_1_737_3908;
   wire n_1_737_3909;
   wire n_1_737_3910;
   wire n_1_737_3911;
   wire n_1_737_3912;
   wire n_1_737_3913;
   wire n_1_737_3914;
   wire n_1_737_3915;
   wire n_1_737_3916;
   wire n_1_737_3917;
   wire n_1_737_3918;
   wire n_1_737_3919;
   wire n_1_737_3920;
   wire n_1_737_3921;
   wire n_1_737_3922;
   wire n_1_737_3923;
   wire n_1_737_3924;
   wire n_1_737_3925;
   wire n_1_737_3926;
   wire n_1_737_3927;
   wire n_1_737_3928;
   wire n_1_737_3929;
   wire n_1_737_3930;
   wire n_1_737_3931;
   wire n_1_737_3932;
   wire n_1_737_3933;
   wire n_1_737_3934;
   wire n_1_737_3935;
   wire n_1_737_3936;
   wire n_1_737_3937;
   wire n_1_737_3938;
   wire n_1_737_3939;
   wire n_1_737_3940;
   wire n_1_737_3941;
   wire n_1_737_3942;
   wire n_1_737_3943;
   wire n_1_737_3944;
   wire n_1_737_3945;
   wire n_1_737_3946;
   wire n_1_737_3947;
   wire n_1_737_3948;
   wire n_1_737_3949;
   wire n_1_737_3950;
   wire n_1_737_3951;
   wire n_1_737_3952;
   wire n_1_737_3953;
   wire n_1_737_3954;
   wire n_1_737_3955;
   wire n_1_737_3956;
   wire n_1_737_3957;
   wire n_1_737_3958;
   wire n_1_737_3959;
   wire n_1_737_3960;
   wire n_1_737_3961;
   wire n_1_737_3962;
   wire n_1_737_3963;
   wire n_1_737_3964;
   wire n_1_737_3965;
   wire n_1_737_3966;
   wire n_1_737_3967;
   wire n_1_737_3968;
   wire n_1_737_3969;
   wire n_1_737_3970;
   wire n_1_737_3971;
   wire n_1_737_3972;
   wire n_1_737_3973;
   wire n_1_737_3974;
   wire n_1_737_3975;
   wire n_1_737_3976;
   wire n_1_737_3977;
   wire n_1_737_3978;
   wire n_1_737_3979;
   wire n_1_737_3980;
   wire n_1_737_3981;
   wire n_1_737_3982;
   wire n_1_737_3983;
   wire n_1_737_3984;
   wire n_1_737_3985;
   wire n_1_737_3986;
   wire n_1_737_3987;
   wire n_1_737_3988;
   wire n_1_737_3989;
   wire n_1_737_3990;
   wire n_1_737_3991;
   wire n_1_737_3992;
   wire n_1_737_3993;
   wire n_1_737_3994;
   wire n_1_737_3995;
   wire n_1_737_3996;
   wire n_1_737_3997;
   wire n_1_737_3998;
   wire n_1_737_3999;
   wire n_1_737_4000;
   wire n_1_737_4001;
   wire n_1_737_4002;
   wire n_1_737_4003;
   wire n_1_737_4004;
   wire n_1_737_4005;
   wire n_1_737_4006;
   wire n_1_737_4007;
   wire n_1_737_4008;
   wire n_1_737_4009;
   wire n_1_737_4010;
   wire n_1_737_4011;
   wire n_1_737_4012;
   wire n_1_737_4013;
   wire n_1_737_4014;
   wire n_1_737_4015;
   wire n_1_737_4016;
   wire n_1_737_4017;
   wire n_1_737_4018;
   wire n_1_737_4019;
   wire n_1_737_4020;
   wire n_1_737_4021;
   wire n_1_737_4022;
   wire n_1_737_4023;
   wire n_1_737_4024;
   wire n_1_737_4025;
   wire n_1_737_4026;
   wire n_1_737_4027;
   wire n_1_737_4028;
   wire n_1_737_4029;
   wire n_1_737_4030;
   wire n_1_737_4031;
   wire n_1_737_4032;
   wire n_1_737_4033;
   wire n_1_737_4034;
   wire n_1_737_4035;
   wire n_1_737_4036;
   wire n_1_737_4037;
   wire n_1_737_4038;
   wire n_1_737_4039;
   wire n_1_737_4040;
   wire n_1_737_4041;
   wire n_1_737_4042;
   wire n_1_737_4043;
   wire n_1_737_4044;
   wire n_1_737_4045;
   wire n_1_737_4046;
   wire n_1_737_4047;
   wire n_1_737_4048;
   wire n_1_737_4049;
   wire n_1_737_4050;
   wire n_1_737_4051;
   wire n_1_737_4052;
   wire n_1_737_4053;
   wire n_1_737_4054;
   wire n_1_737_4055;
   wire n_1_737_4056;
   wire n_1_737_4057;
   wire n_1_737_4058;
   wire n_1_737_4059;
   wire n_1_737_4060;
   wire n_1_737_4061;
   wire n_1_737_4062;
   wire n_1_737_4063;
   wire n_1_737_4064;
   wire n_1_737_4065;
   wire n_1_737_4066;
   wire n_1_737_4067;
   wire n_1_737_4068;
   wire n_1_737_4069;
   wire n_1_737_4070;
   wire n_1_737_4071;
   wire n_1_737_4072;
   wire n_1_737_4073;
   wire n_1_737_4074;
   wire n_1_737_4075;
   wire n_1_737_4076;
   wire n_1_737_4077;
   wire n_1_737_4078;
   wire n_1_737_4079;
   wire n_1_737_4080;
   wire n_1_737_4081;
   wire n_1_737_4082;
   wire n_1_737_4083;
   wire n_1_737_4084;
   wire n_1_737_4085;
   wire n_1_737_4086;
   wire n_1_737_4087;
   wire n_1_737_4088;
   wire n_1_737_4089;
   wire n_1_737_4090;
   wire n_1_737_4091;
   wire n_1_737_4093;
   wire n_1_737_4094;
   wire n_1_737_4095;
   wire n_1_737_4096;
   wire n_1_737_4097;
   wire n_1_737_4098;
   wire n_1_737_4099;
   wire n_1_737_4100;
   wire n_1_737_4101;
   wire n_1_737_4102;
   wire n_1_737_4103;
   wire n_1_737_4104;
   wire n_1_737_4105;
   wire n_1_737_4106;
   wire n_1_737_4107;
   wire n_1_737_4108;
   wire n_1_737_4109;
   wire n_1_737_4110;
   wire n_1_737_4111;
   wire n_1_737_4112;
   wire n_1_737_4113;
   wire n_1_737_4114;
   wire n_1_737_4115;
   wire n_1_737_4116;
   wire n_1_737_4117;
   wire n_1_737_4118;
   wire n_1_737_4119;
   wire n_1_737_4120;
   wire n_1_737_4121;
   wire n_1_737_4122;
   wire n_1_737_4123;
   wire n_1_737_4124;
   wire n_1_737_4125;
   wire n_1_737_4126;
   wire n_1_737_4127;
   wire n_1_737_4128;
   wire n_1_737_4129;
   wire n_1_737_4130;
   wire n_1_737_4131;
   wire n_1_737_4132;
   wire n_1_737_4133;
   wire n_1_737_4134;
   wire n_1_737_4135;
   wire n_1_737_4136;
   wire n_1_737_4137;
   wire n_1_737_4138;
   wire n_1_737_4139;
   wire n_1_737_4140;
   wire n_1_737_4141;
   wire n_1_737_4142;
   wire n_1_737_4143;
   wire n_1_737_4144;
   wire n_1_737_4145;
   wire n_1_737_4146;
   wire n_1_737_4147;
   wire n_1_737_4148;
   wire n_1_737_4149;
   wire n_1_737_4150;
   wire n_1_737_4151;
   wire n_1_737_4152;
   wire n_1_737_4153;
   wire n_1_737_4154;
   wire n_1_737_4155;
   wire n_1_737_4156;
   wire n_1_737_4157;
   wire n_1_737_4158;
   wire n_1_737_4159;
   wire n_1_737_4160;
   wire n_1_737_4161;
   wire n_1_737_4162;
   wire n_1_737_4163;
   wire n_1_737_4164;
   wire n_1_737_4165;
   wire n_1_737_4166;
   wire n_1_737_4167;
   wire n_1_737_4168;
   wire n_1_737_4169;
   wire n_1_737_4170;
   wire n_1_737_4171;
   wire n_1_737_4172;
   wire n_1_737_4173;
   wire n_1_737_4174;
   wire n_1_737_4175;
   wire n_1_737_4176;
   wire n_1_737_4177;
   wire n_1_737_4178;
   wire n_1_737_4179;
   wire n_1_737_4180;
   wire n_1_737_4181;
   wire n_1_737_4182;
   wire n_1_737_4183;
   wire n_1_737_4184;
   wire n_1_737_4185;
   wire n_1_737_4186;
   wire n_1_737_4187;
   wire n_1_737_4188;
   wire n_1_737_4189;
   wire n_1_737_4190;
   wire n_1_737_4191;
   wire n_1_737_4192;
   wire n_1_737_4193;
   wire n_1_737_4194;
   wire n_1_737_4195;
   wire n_1_737_4196;
   wire n_1_737_4197;
   wire n_1_737_4198;
   wire n_1_737_4199;
   wire n_1_737_4200;
   wire n_1_737_4201;
   wire n_1_737_4202;
   wire n_1_737_4203;
   wire n_1_737_4204;
   wire n_1_737_4205;
   wire n_1_737_4206;
   wire n_1_737_4207;
   wire n_1_737_4208;
   wire n_1_737_4209;
   wire n_1_737_4210;
   wire n_1_737_4211;
   wire n_1_737_4212;
   wire n_1_737_4213;
   wire n_1_737_4214;
   wire n_1_737_4215;
   wire n_1_737_4216;
   wire n_1_737_4217;
   wire n_1_737_4218;
   wire n_1_737_4219;
   wire n_1_737_4220;
   wire n_1_737_4221;
   wire n_1_737_4222;
   wire n_1_737_4223;
   wire n_1_737_4224;
   wire n_1_737_4225;
   wire n_1_737_4226;
   wire n_1_737_4227;
   wire n_1_737_4228;
   wire n_1_737_4229;
   wire n_1_737_4230;
   wire n_1_737_4231;
   wire n_1_737_4232;
   wire n_1_737_4233;
   wire n_1_737_4234;
   wire n_1_737_4235;
   wire n_1_737_4236;
   wire n_1_737_4237;
   wire n_1_737_4238;
   wire n_1_737_4239;
   wire n_1_737_4240;
   wire n_1_737_4241;
   wire n_1_737_4242;
   wire n_1_737_4243;
   wire n_1_737_4244;
   wire n_1_737_4245;
   wire n_1_737_4246;
   wire n_1_737_4247;
   wire n_1_737_4248;
   wire n_1_737_4249;
   wire n_1_737_4250;
   wire n_1_737_4251;
   wire n_1_737_4252;
   wire n_1_737_4253;
   wire n_1_737_4254;
   wire n_1_737_4255;
   wire n_1_737_4256;
   wire n_1_737_4257;
   wire n_1_737_4258;
   wire n_1_737_4259;
   wire n_1_737_4260;
   wire n_1_737_4261;
   wire n_1_737_4262;
   wire n_1_737_4263;
   wire n_1_737_4264;
   wire n_1_737_4265;
   wire n_1_737_4266;
   wire n_1_737_4267;
   wire n_1_737_4268;
   wire n_1_737_4269;
   wire n_1_737_4270;
   wire n_1_737_4271;
   wire n_1_737_4272;
   wire n_1_737_4273;
   wire n_1_737_4274;
   wire n_1_737_4275;
   wire n_1_737_4276;
   wire n_1_737_4277;
   wire n_1_737_4278;
   wire n_1_737_4279;
   wire n_1_737_4280;
   wire n_1_737_4281;
   wire n_1_737_4282;
   wire n_1_737_4283;
   wire n_1_737_4284;
   wire n_1_737_4285;
   wire n_1_737_4286;
   wire n_1_737_4287;
   wire n_1_737_4288;
   wire n_1_737_4289;
   wire n_1_737_4290;
   wire n_1_737_4291;
   wire n_1_737_4292;
   wire n_1_737_4293;
   wire n_1_737_4294;
   wire n_1_737_4295;
   wire n_1_737_4296;
   wire n_1_737_4297;
   wire n_1_737_4298;
   wire n_1_737_4299;
   wire n_1_737_4300;
   wire n_1_737_4301;
   wire n_1_737_4302;
   wire n_1_737_4303;
   wire n_1_737_4304;
   wire n_1_737_4305;
   wire n_1_737_4306;
   wire n_1_737_4307;
   wire n_1_737_4308;
   wire n_1_737_4309;
   wire n_1_737_4310;
   wire n_1_737_4311;
   wire n_1_737_4312;
   wire n_1_737_4313;
   wire n_1_737_4314;
   wire n_1_737_4315;
   wire n_1_737_4316;
   wire n_1_737_4317;
   wire n_1_737_4318;
   wire n_1_737_4319;
   wire n_1_737_4320;
   wire n_1_737_4321;
   wire n_1_737_4322;
   wire n_1_737_4323;
   wire n_1_737_4324;
   wire n_1_737_4325;
   wire n_1_737_4326;
   wire n_1_737_4327;
   wire n_1_737_4328;
   wire n_1_737_4329;
   wire n_1_737_4330;
   wire n_1_737_4331;
   wire n_1_737_4332;
   wire n_1_737_4333;
   wire n_1_737_4334;
   wire n_1_737_4335;
   wire n_1_737_4336;
   wire n_1_737_4337;
   wire n_1_737_4338;
   wire n_1_737_4339;
   wire n_1_737_4340;
   wire n_1_737_4341;
   wire n_1_737_4342;
   wire n_1_737_4343;
   wire n_1_737_4344;
   wire n_1_737_4345;
   wire n_1_737_4346;
   wire n_1_737_4347;
   wire n_1_737_4348;
   wire n_1_737_4349;
   wire n_1_737_4350;
   wire n_1_737_4351;
   wire n_1_737_4352;
   wire n_1_737_4353;
   wire n_1_737_4354;
   wire n_1_737_4355;
   wire n_1_737_4356;
   wire n_1_737_4357;
   wire n_1_737_4358;
   wire n_1_737_4359;
   wire n_1_737_4360;
   wire n_1_737_4361;
   wire n_1_737_4362;
   wire n_1_737_4363;
   wire n_1_737_4364;
   wire n_1_737_4365;
   wire n_1_737_4366;
   wire n_1_737_4367;
   wire n_1_737_4368;
   wire n_1_737_4369;
   wire n_1_737_4370;
   wire n_1_737_4371;
   wire n_1_737_4372;
   wire n_1_737_4373;
   wire n_1_737_4374;
   wire n_1_737_4375;
   wire n_1_737_4376;
   wire n_1_737_4377;
   wire n_1_737_4378;
   wire n_1_737_4379;
   wire n_1_737_4380;
   wire n_1_737_4381;
   wire n_1_737_4382;
   wire n_1_737_4383;
   wire n_1_737_4384;
   wire n_1_737_4385;
   wire n_1_737_4386;
   wire n_1_737_4387;
   wire n_1_737_4388;
   wire n_1_737_4389;
   wire n_1_737_4390;
   wire n_1_737_4391;
   wire n_1_737_4392;
   wire n_1_737_4393;
   wire n_1_737_4394;
   wire n_1_737_4395;
   wire n_1_737_4396;
   wire n_1_737_4397;
   wire n_1_737_4398;
   wire n_1_737_4399;
   wire n_1_737_4403;
   wire n_1_737_4405;
   wire n_1_737_4406;
   wire n_1_737_4407;
   wire n_1_737_4408;
   wire n_1_737_4409;
   wire n_1_737_4410;
   wire n_1_737_4411;
   wire n_1_737_4412;
   wire n_1_737_4413;
   wire n_1_737_4414;
   wire n_1_737_4415;
   wire n_1_737_4416;
   wire n_1_737_4417;
   wire n_1_737_4418;
   wire n_1_737_4419;
   wire n_1_737_4420;
   wire n_1_737_4421;
   wire n_1_737_4422;
   wire n_1_737_4423;
   wire n_1_737_4424;
   wire n_1_737_4425;
   wire n_1_737_4426;
   wire n_1_737_4427;
   wire n_1_737_4428;
   wire n_1_737_4429;
   wire n_1_737_4430;
   wire n_1_737_4431;
   wire n_1_737_4432;
   wire n_1_737_4433;
   wire n_1_737_4434;
   wire n_1_737_4435;
   wire n_1_737_4436;
   wire n_1_737_4437;
   wire n_1_737_4438;
   wire n_1_737_4439;
   wire n_1_737_4440;
   wire n_1_737_4441;
   wire n_1_737_4442;
   wire n_1_737_4443;
   wire n_1_737_4444;
   wire n_1_737_4445;
   wire n_1_737_4446;
   wire n_1_737_4447;
   wire n_1_737_4448;
   wire n_1_737_4449;
   wire n_1_737_4450;
   wire n_1_737_4451;
   wire n_1_737_4452;
   wire n_1_737_4454;
   wire n_1_737_4455;
   wire n_1_737_4456;
   wire n_1_737_4457;
   wire n_1_737_4458;
   wire n_1_737_4459;
   wire n_1_737_4460;
   wire n_1_737_4461;
   wire n_1_737_4462;
   wire n_1_737_4463;
   wire n_1_737_4464;
   wire n_1_737_4465;
   wire n_1_737_4466;
   wire n_1_737_4467;
   wire n_1_737_4468;
   wire n_1_737_4469;
   wire n_1_737_4470;
   wire n_1_737_4471;
   wire n_1_737_4472;
   wire n_1_737_4473;
   wire n_1_737_4474;
   wire n_1_737_4475;
   wire n_1_737_4476;
   wire n_1_737_4477;
   wire n_1_737_4478;
   wire n_1_737_4479;
   wire n_1_737_4480;
   wire n_1_737_4481;
   wire n_1_737_4482;
   wire n_1_737_4483;
   wire n_1_737_4484;
   wire n_1_737_4485;
   wire n_1_737_4486;
   wire n_1_737_4487;
   wire n_1_737_4488;
   wire n_1_737_4489;
   wire n_1_737_4490;
   wire n_1_737_4491;
   wire n_1_737_4492;
   wire n_1_737_4493;
   wire n_1_737_4494;
   wire n_1_737_4495;
   wire n_1_737_4496;
   wire n_1_737_4497;
   wire n_1_737_4498;
   wire n_1_737_4499;
   wire n_1_737_4500;
   wire n_1_737_4501;
   wire n_1_737_4502;
   wire n_1_737_4503;
   wire n_1_737_4504;
   wire n_1_737_4505;
   wire n_1_737_4506;
   wire n_1_737_4507;
   wire n_1_737_4508;
   wire n_1_737_4509;
   wire n_1_737_4510;
   wire n_1_737_4511;
   wire n_1_737_4512;
   wire n_1_737_4513;
   wire n_1_737_4514;
   wire n_1_737_4515;
   wire n_1_737_4516;
   wire n_1_737_4517;
   wire n_1_737_4518;
   wire n_1_737_4519;
   wire n_1_737_4520;
   wire n_1_737_4521;
   wire n_1_737_4522;
   wire n_1_737_4523;
   wire n_1_737_4524;
   wire n_1_737_4525;
   wire n_1_737_4526;
   wire n_1_737_4527;
   wire n_1_737_4528;
   wire n_1_737_4529;
   wire n_1_737_4530;
   wire n_1_737_4531;
   wire n_1_737_4532;
   wire n_1_737_4533;
   wire n_1_737_4534;
   wire n_1_737_4535;
   wire n_1_737_4536;
   wire n_1_737_4537;
   wire n_1_737_4538;
   wire n_1_737_4539;
   wire n_1_737_4540;
   wire n_1_737_4541;
   wire n_1_737_4542;
   wire n_1_737_4543;
   wire n_1_737_4544;
   wire n_1_737_4545;
   wire n_1_737_4546;
   wire n_1_737_4547;
   wire n_1_737_4548;
   wire n_1_737_4549;
   wire n_1_737_4550;
   wire n_1_737_4551;
   wire n_1_737_4552;
   wire n_1_737_4553;
   wire n_1_737_4554;
   wire n_1_737_4555;
   wire n_1_737_4556;
   wire n_1_737_4557;
   wire n_1_737_4558;
   wire n_1_737_4559;
   wire n_1_737_4560;
   wire n_1_737_4561;
   wire n_1_737_4562;
   wire n_1_737_4563;
   wire n_1_737_4564;
   wire n_1_737_4565;
   wire n_1_737_4566;
   wire n_1_737_4567;
   wire n_1_737_4568;
   wire n_1_737_4569;
   wire n_1_737_4570;
   wire n_1_737_4571;
   wire n_1_737_4572;
   wire n_1_737_4573;
   wire n_1_737_4574;
   wire n_1_737_4575;
   wire n_1_737_4576;
   wire n_1_737_4577;
   wire n_1_737_4578;
   wire n_1_737_4579;
   wire n_1_737_4580;
   wire n_1_737_4581;
   wire n_1_737_4582;
   wire n_1_737_4583;
   wire n_1_737_4584;
   wire n_1_737_4585;
   wire n_1_737_4586;
   wire n_1_737_4587;
   wire n_1_737_4588;
   wire n_1_737_4589;
   wire n_1_737_4590;
   wire n_1_737_4591;
   wire n_1_737_4592;
   wire n_1_737_4593;
   wire n_1_737_4594;
   wire n_1_737_4595;
   wire n_1_737_4596;
   wire n_1_737_4597;
   wire n_1_737_4598;
   wire n_1_737_4599;
   wire n_1_737_4600;
   wire n_1_737_4601;
   wire n_1_737_4602;
   wire n_1_737_4603;
   wire n_1_737_4604;
   wire n_1_737_4605;
   wire n_1_737_4606;
   wire n_1_737_4607;
   wire n_1_737_4608;
   wire n_1_737_4609;
   wire n_1_737_4610;
   wire n_1_737_4611;
   wire n_1_737_4612;
   wire n_1_737_4613;
   wire n_1_737_4614;
   wire n_1_737_4615;
   wire n_1_737_4616;
   wire n_1_737_4617;
   wire n_1_737_4618;
   wire n_1_737_4619;
   wire n_1_737_4620;
   wire n_1_737_4621;
   wire n_1_737_4622;
   wire n_1_737_4623;
   wire n_1_737_4624;
   wire n_1_737_4625;
   wire n_1_737_4626;
   wire n_1_737_4627;
   wire n_1_737_4628;
   wire n_1_737_4629;
   wire n_1_737_4630;
   wire n_1_737_4631;
   wire n_1_737_4632;
   wire n_1_737_4633;
   wire n_1_737_4634;
   wire n_1_737_4635;
   wire n_1_737_4636;
   wire n_1_737_4637;
   wire n_1_737_4638;
   wire n_1_737_4639;
   wire n_1_737_4640;
   wire n_1_737_4641;
   wire n_1_737_4642;
   wire n_1_737_4643;
   wire n_1_737_4644;
   wire n_1_737_4645;
   wire n_1_737_4646;
   wire n_1_737_4647;
   wire n_1_737_4648;
   wire n_1_737_4649;
   wire n_1_737_4650;
   wire n_1_737_4651;
   wire n_1_737_4652;
   wire n_1_737_4653;
   wire n_1_737_4654;
   wire n_1_737_4655;
   wire n_1_737_4656;
   wire n_1_737_4657;
   wire n_1_737_4658;
   wire n_1_737_4659;
   wire n_1_737_4660;
   wire n_1_737_4661;
   wire n_1_737_4662;
   wire n_1_737_4663;
   wire n_1_737_4664;
   wire n_1_737_4665;
   wire n_1_737_4666;
   wire n_1_737_4667;
   wire n_1_737_4668;
   wire n_1_737_4669;
   wire n_1_737_4670;
   wire n_1_737_4671;
   wire n_1_737_4672;
   wire n_1_737_4673;
   wire n_1_737_4674;
   wire n_1_737_4675;
   wire n_1_737_4676;
   wire n_1_737_4677;
   wire n_1_737_4678;
   wire n_1_737_4679;
   wire n_1_737_4680;
   wire n_1_737_4681;
   wire n_1_737_4682;
   wire n_1_737_4683;
   wire n_1_737_4684;
   wire n_1_737_4685;
   wire n_1_737_4686;
   wire n_1_737_4687;
   wire n_1_737_4688;
   wire n_1_737_4689;
   wire n_1_737_4690;
   wire n_1_737_4691;
   wire n_1_737_4692;
   wire n_1_737_4693;
   wire n_1_737_4694;
   wire n_1_737_4695;
   wire n_1_737_4696;
   wire n_1_737_4697;
   wire n_1_737_4698;
   wire n_1_737_4699;
   wire n_1_737_4700;
   wire n_1_737_4701;
   wire n_1_737_4702;
   wire n_1_737_4703;
   wire n_1_737_4704;
   wire n_1_737_4705;
   wire n_1_737_4706;
   wire n_1_737_4707;
   wire n_1_737_4708;
   wire n_1_737_4709;
   wire n_1_737_4710;
   wire n_1_737_4711;
   wire n_1_737_4712;
   wire n_1_737_4713;
   wire n_1_737_4714;
   wire n_1_737_4715;
   wire n_1_737_4716;
   wire n_1_737_4717;
   wire n_1_737_4718;
   wire n_1_737_4719;
   wire n_1_737_4720;
   wire n_1_737_4721;
   wire n_1_737_4722;
   wire n_1_737_4723;
   wire n_1_737_4724;
   wire n_1_737_4725;
   wire n_1_737_4726;
   wire n_1_737_4727;
   wire n_1_737_4728;
   wire n_1_737_4729;
   wire n_1_737_4730;
   wire n_1_737_4731;
   wire n_1_737_4732;
   wire n_1_737_4733;
   wire n_1_737_4734;
   wire n_1_737_4735;
   wire n_1_737_4736;
   wire n_1_737_4737;
   wire n_1_737_4738;
   wire n_1_737_4739;
   wire n_1_737_4740;
   wire n_1_737_4741;
   wire n_1_737_4742;
   wire n_1_737_4743;
   wire n_1_737_4744;
   wire n_1_737_4745;
   wire n_1_737_4746;
   wire n_1_737_4747;
   wire n_1_737_4748;
   wire n_1_737_4749;
   wire n_1_737_4750;
   wire n_1_737_4751;
   wire n_1_737_4752;
   wire n_1_737_4753;
   wire n_1_737_4754;
   wire n_1_737_4755;
   wire n_1_737_4756;
   wire n_1_737_4757;
   wire n_1_737_4758;
   wire n_1_737_4759;
   wire n_1_737_4760;
   wire n_1_737_4761;
   wire n_1_737_4762;
   wire n_1_737_4763;
   wire n_1_737_4764;
   wire n_1_737_4765;
   wire n_1_737_4766;
   wire n_1_737_4767;
   wire n_1_737_4768;
   wire n_1_737_4769;
   wire n_1_737_4770;
   wire n_1_737_4771;
   wire n_1_737_4772;
   wire n_1_737_4773;
   wire n_1_737_4774;
   wire n_1_737_4775;
   wire n_1_737_4776;
   wire n_1_737_4777;
   wire n_1_737_4778;
   wire n_1_737_4779;
   wire n_1_737_4780;
   wire n_1_737_4781;
   wire n_1_737_4782;
   wire n_1_737_4783;
   wire n_1_737_4784;
   wire n_1_737_4785;
   wire n_1_737_4786;
   wire n_1_737_4787;
   wire n_1_737_4788;
   wire n_1_737_4789;
   wire n_1_737_4790;
   wire n_1_737_4791;
   wire n_1_737_4792;
   wire n_1_737_4793;
   wire n_1_737_4794;
   wire n_1_737_4795;
   wire n_1_737_4796;
   wire n_1_737_4797;
   wire n_1_737_4798;
   wire n_1_737_4799;
   wire n_1_737_4800;
   wire n_1_737_4801;
   wire n_1_737_4802;
   wire n_1_737_4803;
   wire n_1_737_4804;
   wire n_1_737_4805;
   wire n_1_737_4806;
   wire n_1_737_4807;
   wire n_1_737_4808;
   wire n_1_737_4809;
   wire n_1_737_4810;
   wire n_1_737_4811;
   wire n_1_737_4812;
   wire n_1_737_4813;
   wire n_1_737_4814;
   wire n_1_737_4815;
   wire n_1_737_4816;
   wire n_1_737_4817;
   wire n_1_737_4818;
   wire n_1_737_4819;
   wire n_1_737_4820;
   wire n_1_737_4821;
   wire n_1_737_4822;
   wire n_1_737_4823;
   wire n_1_737_4824;
   wire n_1_737_4825;
   wire n_1_737_4826;
   wire n_1_737_4827;
   wire n_1_737_4828;
   wire n_1_737_4829;
   wire n_1_737_4830;
   wire n_1_737_4831;
   wire n_1_737_4832;
   wire n_1_737_4833;
   wire n_1_737_4834;
   wire n_1_737_4835;
   wire n_1_737_4836;
   wire n_1_737_4837;
   wire n_1_737_4838;
   wire n_1_737_4839;
   wire n_1_737_4840;
   wire n_1_737_4841;
   wire n_1_737_4842;
   wire n_1_737_4843;
   wire n_1_737_4844;
   wire n_1_737_4845;
   wire n_1_737_4846;
   wire n_1_737_4847;
   wire n_1_737_4848;
   wire n_1_737_4849;
   wire n_1_737_4850;
   wire n_1_737_4851;
   wire n_1_737_4852;
   wire n_1_737_4853;
   wire n_1_737_4854;
   wire n_1_737_4855;
   wire n_1_737_4856;
   wire n_1_737_4857;
   wire n_1_737_4858;
   wire n_1_737_4859;
   wire n_1_737_4860;
   wire n_1_737_4861;
   wire n_1_737_4862;
   wire n_1_737_4863;
   wire n_1_737_4864;
   wire n_1_737_4865;
   wire n_1_737_4866;
   wire n_1_737_4867;
   wire n_1_737_4868;
   wire n_1_737_4869;
   wire n_1_737_4870;
   wire n_1_737_4871;
   wire n_1_737_4872;
   wire n_1_737_4873;
   wire n_1_737_4874;
   wire n_1_737_4875;
   wire n_1_737_4876;
   wire n_1_737_4877;
   wire n_1_737_4878;
   wire n_1_737_4879;
   wire n_1_737_4880;
   wire n_1_737_4881;
   wire n_1_737_4882;
   wire n_1_737_4883;
   wire n_1_737_4884;
   wire n_1_737_4885;
   wire n_1_737_4886;
   wire n_1_737_4887;
   wire n_1_737_4888;
   wire n_1_737_4889;
   wire n_1_737_4890;
   wire n_1_737_4891;
   wire n_1_737_4892;
   wire n_1_737_4893;
   wire n_1_737_4894;
   wire n_1_737_4895;
   wire n_1_737_4896;
   wire n_1_737_4897;
   wire n_1_737_4898;
   wire n_1_737_4899;
   wire n_1_737_4900;
   wire n_1_737_4901;
   wire n_1_737_4902;
   wire n_1_737_4903;
   wire n_1_737_4904;
   wire n_1_737_4905;
   wire n_1_737_4906;
   wire n_1_737_4907;
   wire n_1_737_4908;
   wire n_1_737_4909;
   wire n_1_737_4910;
   wire n_1_737_4911;
   wire n_1_737_4912;
   wire n_1_737_4913;
   wire n_1_737_4914;
   wire n_1_737_4915;
   wire n_1_737_4916;
   wire n_1_737_4917;
   wire n_1_737_4918;
   wire n_1_737_4919;
   wire n_1_737_4920;
   wire n_1_737_4921;
   wire n_1_737_4922;
   wire n_1_737_4923;
   wire n_1_737_4924;
   wire n_1_737_4925;
   wire n_1_737_4926;
   wire n_1_737_4927;
   wire n_1_737_4928;
   wire n_1_737_4929;
   wire n_1_737_4930;
   wire n_1_737_4931;
   wire n_1_737_4932;
   wire n_1_737_4933;
   wire n_1_737_4934;
   wire n_1_737_4935;
   wire n_1_737_4936;
   wire n_1_737_4937;
   wire n_1_737_4938;
   wire n_1_737_4939;
   wire n_1_737_4940;
   wire n_1_737_4941;
   wire n_1_737_4942;
   wire n_1_737_4943;
   wire n_1_737_4944;
   wire n_1_737_4945;
   wire n_1_737_4946;
   wire n_1_737_4947;
   wire n_1_737_4948;
   wire n_1_737_4949;
   wire n_1_737_4950;
   wire n_1_737_4951;
   wire n_1_737_4952;
   wire n_1_737_4953;
   wire n_1_737_4954;
   wire n_1_737_4955;
   wire n_1_737_4956;
   wire n_1_737_4957;
   wire n_1_737_4958;
   wire n_1_737_4959;
   wire n_1_737_4960;
   wire n_1_737_4961;
   wire n_1_737_4962;
   wire n_1_737_4963;
   wire n_1_737_4964;
   wire n_1_737_4966;
   wire n_1_737_4967;
   wire n_1_737_4968;
   wire n_1_737_4969;
   wire n_1_737_4970;
   wire n_1_737_4971;
   wire n_1_737_4972;
   wire n_1_737_4973;
   wire n_1_737_4974;
   wire n_1_737_4975;
   wire n_1_737_4976;
   wire n_1_737_4977;
   wire n_1_737_4978;
   wire n_1_737_4979;
   wire n_1_737_4980;
   wire n_1_737_4981;
   wire n_1_737_4982;
   wire n_1_737_4983;
   wire n_1_737_4984;
   wire n_1_737_4985;
   wire n_1_737_4986;
   wire n_1_737_4987;
   wire n_1_737_4988;
   wire n_1_737_4989;
   wire n_1_737_4990;
   wire n_1_737_4991;
   wire n_1_737_4992;
   wire n_1_737_4993;
   wire n_1_737_4994;
   wire n_1_737_4995;
   wire n_1_737_4996;
   wire n_1_737_4997;
   wire n_1_737_4998;
   wire n_1_737_4999;
   wire n_1_737_5000;
   wire n_1_737_5001;
   wire n_1_737_5002;
   wire n_1_737_5003;
   wire n_1_737_5004;
   wire n_1_737_5005;
   wire n_1_737_5006;
   wire n_1_737_5007;
   wire n_1_737_5008;
   wire n_1_737_5009;
   wire n_1_737_5010;
   wire n_1_737_5011;
   wire n_1_737_5012;
   wire n_1_737_5013;
   wire n_1_737_5014;
   wire n_1_737_5015;
   wire n_1_737_5016;
   wire n_1_737_5017;
   wire n_1_737_5018;
   wire n_1_737_5019;
   wire n_1_737_5020;
   wire n_1_737_5021;
   wire n_1_737_5022;
   wire n_1_737_5023;
   wire n_1_737_5024;
   wire n_1_737_5025;
   wire n_1_737_5026;
   wire n_1_737_5027;
   wire n_1_737_5028;
   wire n_1_737_5029;
   wire n_1_737_5030;
   wire n_1_737_5031;
   wire n_1_737_5032;
   wire n_1_737_5033;
   wire n_1_737_5034;
   wire n_1_737_5035;
   wire n_1_737_5036;
   wire n_1_737_5037;
   wire n_1_737_5038;
   wire n_1_737_5039;
   wire n_1_737_5040;
   wire n_1_737_5041;
   wire n_1_737_5042;
   wire n_1_737_5043;
   wire n_1_737_5044;
   wire n_1_737_5045;
   wire n_1_737_5046;
   wire n_1_737_5047;
   wire n_1_737_5048;
   wire n_1_737_5049;
   wire n_1_737_5050;
   wire n_1_737_5051;
   wire n_1_737_5052;
   wire n_1_737_5053;
   wire n_1_737_5054;
   wire n_1_737_5055;
   wire n_1_737_5056;
   wire n_1_737_5057;
   wire n_1_737_5058;
   wire n_1_737_5059;
   wire n_1_737_5060;
   wire n_1_737_5061;
   wire n_1_737_5062;
   wire n_1_737_5063;
   wire n_1_737_5064;
   wire n_1_737_5065;
   wire n_1_737_5066;
   wire n_1_737_5067;
   wire n_1_737_5068;
   wire n_1_737_5069;
   wire n_1_737_5070;
   wire n_1_737_5071;
   wire n_1_737_5072;
   wire n_1_737_5073;
   wire n_1_737_5074;
   wire n_1_737_5075;
   wire n_1_737_5076;
   wire n_1_737_5077;
   wire n_1_737_5078;
   wire n_1_737_5079;
   wire n_1_737_5080;
   wire n_1_737_5081;
   wire n_1_737_5082;
   wire n_1_737_5083;
   wire n_1_737_5084;
   wire n_1_737_5085;
   wire n_1_737_5086;
   wire n_1_737_5087;
   wire n_1_737_5088;
   wire n_1_737_5089;
   wire n_1_737_5090;
   wire n_1_737_5091;
   wire n_1_737_5092;
   wire n_1_737_5093;
   wire n_1_737_5094;
   wire n_1_737_5095;
   wire n_1_737_5096;
   wire n_1_737_5097;
   wire n_1_737_5098;
   wire n_1_737_5099;
   wire n_1_737_5100;
   wire n_1_737_5101;
   wire n_1_737_5102;
   wire n_1_737_5103;
   wire n_1_737_5104;
   wire n_1_737_5105;
   wire n_1_737_5106;
   wire n_1_737_5107;
   wire n_1_737_5108;
   wire n_1_737_5109;
   wire n_1_737_5110;
   wire n_1_737_5111;
   wire n_1_737_5112;
   wire n_1_737_5113;
   wire n_1_737_5114;
   wire n_1_737_5115;
   wire n_1_737_5116;
   wire n_1_737_5117;
   wire n_1_737_5118;
   wire n_1_737_5119;
   wire n_1_737_5120;
   wire n_1_737_5121;
   wire n_1_737_5122;
   wire n_1_737_5123;
   wire n_1_737_5124;
   wire n_1_737_5125;
   wire n_1_737_5126;
   wire n_1_737_5127;
   wire n_1_737_5128;
   wire n_1_737_5129;
   wire n_1_737_5130;
   wire n_1_737_5131;
   wire n_1_737_5132;
   wire n_1_737_5133;
   wire n_1_737_5134;
   wire n_1_737_5135;
   wire n_1_737_5136;
   wire n_1_737_5137;
   wire n_1_737_5138;
   wire n_1_737_5139;
   wire n_1_737_5140;
   wire n_1_737_5141;
   wire n_1_737_5142;
   wire n_1_737_5143;
   wire n_1_737_5144;
   wire n_1_737_5145;
   wire n_1_737_5146;
   wire n_1_737_5147;
   wire n_1_737_5148;
   wire n_1_737_5149;
   wire n_1_737_5150;
   wire n_1_737_5151;
   wire n_1_737_5152;
   wire n_1_737_5153;
   wire n_1_737_5154;
   wire n_1_737_5155;
   wire n_1_737_5156;
   wire n_1_737_5157;
   wire n_1_737_5158;
   wire n_1_737_5159;
   wire n_1_737_5160;
   wire n_1_737_5161;
   wire n_1_737_5162;
   wire n_1_737_5163;
   wire n_1_737_5164;
   wire n_1_737_5165;
   wire n_1_737_5166;
   wire n_1_737_5168;
   wire n_1_737_5169;
   wire n_1_737_5170;
   wire n_1_737_5171;
   wire n_1_737_5172;
   wire n_1_737_5173;
   wire n_1_737_5174;
   wire n_1_737_5175;
   wire n_1_737_5176;
   wire n_1_737_5177;
   wire n_1_737_5178;
   wire n_1_737_5179;
   wire n_1_737_5180;
   wire n_1_737_5183;
   wire n_1_737_5184;
   wire n_1_737_5185;
   wire n_1_737_5186;
   wire n_1_737_5187;
   wire n_1_737_5188;
   wire n_1_737_5189;
   wire n_1_737_5190;
   wire n_1_737_5191;
   wire n_1_737_5192;
   wire n_1_737_5193;
   wire n_1_737_5194;
   wire n_1_737_5195;
   wire n_1_737_5196;
   wire n_1_737_5197;
   wire n_1_737_5198;
   wire n_1_737_5199;
   wire n_1_737_5200;
   wire n_1_737_5201;
   wire n_1_737_5202;
   wire n_1_737_5203;
   wire n_1_737_5204;
   wire n_1_737_5205;
   wire n_1_737_5206;
   wire n_1_737_5207;
   wire n_1_737_5208;
   wire n_1_737_5209;
   wire n_1_737_5210;
   wire n_1_737_5211;
   wire n_1_737_5212;
   wire n_1_737_5213;
   wire n_1_737_5214;
   wire n_1_737_5215;
   wire n_1_737_5216;
   wire n_1_737_5217;
   wire n_1_737_5218;
   wire n_1_737_5219;
   wire n_1_737_5220;
   wire n_1_737_5221;
   wire n_1_737_5222;
   wire n_1_737_5223;
   wire n_1_737_5224;
   wire n_1_737_5225;
   wire n_1_737_5226;
   wire n_1_737_5227;
   wire n_1_737_5228;
   wire n_1_737_5229;
   wire n_1_737_5230;
   wire n_1_737_5231;
   wire n_1_737_5232;
   wire n_1_737_5233;
   wire n_1_737_5234;
   wire n_1_737_5235;
   wire n_1_737_5236;
   wire n_1_737_5237;
   wire n_1_737_5238;
   wire n_1_737_5239;
   wire n_1_737_5240;
   wire n_1_737_5241;
   wire n_1_737_5242;
   wire n_1_737_5243;
   wire n_1_737_5244;
   wire n_1_737_5245;
   wire n_1_737_5246;
   wire n_1_737_5247;
   wire n_1_737_5248;
   wire n_1_737_5249;
   wire n_1_737_5250;
   wire n_1_737_5251;
   wire n_1_737_5252;
   wire n_1_737_5253;
   wire n_1_737_5254;
   wire n_1_737_5255;
   wire n_1_737_5256;
   wire n_1_737_5257;
   wire n_1_737_5258;
   wire n_1_737_5259;
   wire n_1_737_5260;
   wire n_1_737_5261;
   wire n_1_737_5262;
   wire n_1_737_5263;
   wire n_1_737_5264;
   wire n_1_737_5265;
   wire n_1_737_5266;
   wire n_1_737_5267;
   wire n_1_737_5268;
   wire n_1_737_5269;
   wire n_1_737_5270;
   wire n_1_737_5271;
   wire n_1_737_5272;
   wire n_1_737_5273;
   wire n_1_737_5274;
   wire n_1_737_5275;
   wire n_1_737_5276;
   wire n_1_737_5277;
   wire n_1_737_5278;
   wire n_1_737_5279;
   wire n_1_737_5280;
   wire n_1_737_5281;
   wire n_1_737_5282;
   wire n_1_737_5283;
   wire n_1_737_5284;
   wire n_1_737_5285;
   wire n_1_737_5286;
   wire n_1_737_5287;
   wire n_1_737_5288;
   wire n_1_737_5289;
   wire n_1_737_5290;
   wire n_1_737_5291;
   wire n_1_737_5292;
   wire n_1_737_5293;
   wire n_1_737_5294;
   wire n_1_737_5295;
   wire n_1_737_5296;
   wire n_1_737_5297;
   wire n_1_737_5298;
   wire n_1_737_5299;
   wire n_1_737_5300;
   wire n_1_737_5301;
   wire n_1_737_5302;
   wire n_1_737_5303;
   wire n_1_737_5304;
   wire n_1_737_5305;
   wire n_1_737_5306;
   wire n_1_737_5307;
   wire n_1_737_5308;
   wire n_1_737_5309;
   wire n_1_737_5310;
   wire n_1_737_5311;
   wire n_1_737_5312;
   wire n_1_737_5313;
   wire n_1_737_5314;
   wire n_1_737_5315;
   wire n_1_737_5316;
   wire n_1_737_5317;
   wire n_1_737_5318;
   wire n_1_737_5319;
   wire n_1_737_5320;
   wire n_1_737_5321;
   wire n_1_737_5322;
   wire n_1_737_5323;
   wire n_1_737_5324;
   wire n_1_737_5325;
   wire n_1_737_5326;
   wire n_1_737_5327;
   wire n_1_737_5328;
   wire n_1_737_5329;
   wire n_1_737_5330;
   wire n_1_737_5331;
   wire n_1_737_5332;
   wire n_1_737_5333;
   wire n_1_737_5334;
   wire n_1_737_5335;
   wire n_1_737_5336;
   wire n_1_737_5338;
   wire n_1_737_5339;
   wire n_1_737_5340;
   wire n_1_737_5341;
   wire n_1_737_5342;
   wire n_1_737_5343;
   wire n_1_737_5344;
   wire n_1_737_5345;
   wire n_1_737_5346;
   wire n_1_737_5347;
   wire n_1_737_5348;
   wire n_1_737_5349;
   wire n_1_737_5350;
   wire n_1_737_5351;
   wire n_1_737_5352;
   wire n_1_737_5353;
   wire n_1_737_5354;
   wire n_1_737_5355;
   wire n_1_737_5356;
   wire n_1_737_5357;
   wire n_1_737_5358;
   wire n_1_737_5359;
   wire n_1_737_5360;
   wire n_1_737_5361;
   wire n_1_737_5362;
   wire n_1_737_5363;
   wire n_1_737_5364;
   wire n_1_737_5365;
   wire n_1_737_5366;
   wire n_1_737_5367;
   wire n_1_737_5368;
   wire n_1_737_5369;
   wire n_1_737_5370;
   wire n_1_737_5371;
   wire n_1_737_5372;
   wire n_1_737_5373;
   wire n_1_737_5374;
   wire n_1_737_5375;
   wire n_1_737_5376;
   wire n_1_737_5377;
   wire n_1_737_5378;
   wire n_1_737_5379;
   wire n_1_737_5380;
   wire n_1_737_5381;
   wire n_1_737_5382;
   wire n_1_737_5383;
   wire n_1_737_5384;
   wire n_1_737_5385;
   wire n_1_737_5386;
   wire n_1_737_5387;
   wire n_1_737_5388;
   wire n_1_737_5389;
   wire n_1_737_5390;
   wire n_1_737_5391;
   wire n_1_737_5392;
   wire n_1_737_5393;
   wire n_1_737_5394;
   wire n_1_737_5395;
   wire n_1_737_5396;
   wire n_1_737_5397;
   wire n_1_737_5398;
   wire n_1_737_5399;
   wire n_1_737_5400;
   wire n_1_737_5401;
   wire n_1_737_5402;
   wire n_1_737_5403;
   wire n_1_737_5404;
   wire n_1_737_5405;
   wire n_1_737_5406;
   wire n_1_737_5407;
   wire n_1_737_5408;
   wire n_1_737_5409;
   wire n_1_737_5410;
   wire n_1_737_5411;
   wire n_1_737_5412;
   wire n_1_737_5413;
   wire n_1_737_5414;
   wire n_1_737_5415;
   wire n_1_737_5416;
   wire n_1_737_5417;
   wire n_1_737_5418;
   wire n_1_737_5419;
   wire n_1_737_5420;
   wire n_1_737_5421;
   wire n_1_737_5422;
   wire n_1_737_5423;
   wire n_1_737_5424;
   wire n_1_737_5425;
   wire n_1_737_5426;
   wire n_1_737_5427;
   wire n_1_737_5428;
   wire n_1_737_5429;
   wire n_1_737_5430;
   wire n_1_737_5431;
   wire n_1_737_5432;
   wire n_1_737_5433;
   wire n_1_737_5434;
   wire n_1_737_5435;
   wire n_1_737_5436;
   wire n_1_737_5437;
   wire n_1_737_5438;
   wire n_1_737_5439;
   wire n_1_737_5440;
   wire n_1_737_5441;
   wire n_1_737_5442;
   wire n_1_737_5443;
   wire n_1_737_5444;
   wire n_1_737_5445;
   wire n_1_737_5446;
   wire n_1_737_5447;
   wire n_1_737_5448;
   wire n_1_737_5449;
   wire n_1_737_5450;
   wire n_1_737_5451;
   wire n_1_737_5452;
   wire n_1_737_5453;
   wire n_1_737_5454;
   wire n_1_737_5455;
   wire n_1_737_5456;
   wire n_1_737_5457;
   wire n_1_737_5458;
   wire n_1_737_5459;
   wire n_1_737_5460;
   wire n_1_737_5461;
   wire n_1_737_5462;
   wire n_1_737_5463;
   wire n_1_737_5464;
   wire n_1_737_5465;
   wire n_1_737_5466;
   wire n_1_737_5467;
   wire n_1_737_5468;
   wire n_1_737_5469;
   wire n_1_737_5470;
   wire n_1_737_5471;
   wire n_1_737_5472;
   wire n_1_737_5473;
   wire n_1_737_5474;
   wire n_1_737_5475;
   wire n_1_737_5476;
   wire n_1_737_5477;
   wire n_1_737_5478;
   wire n_1_737_5479;
   wire n_1_737_5480;
   wire n_1_737_5481;
   wire n_1_737_5482;
   wire n_1_737_5483;
   wire n_1_737_5484;
   wire n_1_737_5485;
   wire n_1_737_5486;
   wire n_1_737_5487;
   wire n_1_737_5488;
   wire n_1_737_5489;
   wire n_1_737_5490;
   wire n_1_737_5491;
   wire n_1_737_5492;
   wire n_1_737_5493;
   wire n_1_737_5494;
   wire n_1_737_5495;
   wire n_1_737_5496;
   wire n_1_737_5497;
   wire n_1_737_5498;
   wire n_1_737_5499;
   wire n_1_737_5500;
   wire n_1_737_5501;
   wire n_1_737_5502;
   wire n_1_737_5503;
   wire n_1_737_5504;
   wire n_1_737_5505;
   wire n_1_737_5506;
   wire n_1_737_5507;
   wire n_1_737_5508;
   wire n_1_737_5509;
   wire n_1_737_5510;
   wire n_1_737_5511;
   wire n_1_737_5512;
   wire n_1_737_5513;
   wire n_1_737_5514;
   wire n_1_737_5515;
   wire n_1_737_5516;
   wire n_1_737_5517;
   wire n_1_737_5518;
   wire n_1_737_5519;
   wire n_1_737_5520;
   wire n_1_737_5521;
   wire n_1_737_5522;
   wire n_1_737_5523;
   wire n_1_737_5524;
   wire n_1_737_5525;
   wire n_1_737_5526;
   wire n_1_737_5527;
   wire n_1_737_5528;
   wire n_1_737_5529;
   wire n_1_737_5530;
   wire n_1_737_5531;
   wire n_1_737_5532;
   wire n_1_737_5533;
   wire n_1_737_5534;
   wire n_1_737_5535;
   wire n_1_737_5536;
   wire n_1_737_5537;
   wire n_1_737_5538;
   wire n_1_737_5539;
   wire n_1_737_5540;
   wire n_1_737_5541;
   wire n_1_737_5542;
   wire n_1_737_5543;
   wire n_1_737_5544;
   wire n_1_737_5545;
   wire n_1_737_5546;
   wire n_1_737_5547;
   wire n_1_737_5548;
   wire n_1_737_5549;
   wire n_1_737_5550;
   wire n_1_737_5551;
   wire n_1_737_5552;
   wire n_1_737_5553;
   wire n_1_737_5554;
   wire n_1_737_5555;
   wire n_1_737_5556;
   wire n_1_737_5557;
   wire n_1_737_5558;
   wire n_1_737_5559;
   wire n_1_737_5560;
   wire n_1_737_5561;
   wire n_1_737_5562;
   wire n_1_737_5563;
   wire n_1_737_5564;
   wire n_1_737_5565;
   wire n_1_737_5566;
   wire n_1_737_5567;
   wire n_1_737_5568;
   wire n_1_737_5569;
   wire n_1_737_5570;
   wire n_1_737_5571;
   wire n_1_737_5572;
   wire n_1_737_5573;
   wire n_1_737_5574;
   wire n_1_737_5575;
   wire n_1_737_5576;
   wire n_1_737_5577;
   wire n_1_737_5578;
   wire n_1_737_5579;
   wire n_1_737_5580;
   wire n_1_737_5581;
   wire n_1_737_5582;
   wire n_1_737_5583;
   wire n_1_737_5584;
   wire n_1_737_5585;
   wire n_1_737_5586;
   wire n_1_737_5587;
   wire n_1_737_5588;
   wire n_1_737_5589;
   wire n_1_737_5590;
   wire n_1_737_5591;
   wire n_1_737_5592;
   wire n_1_737_5593;
   wire n_1_737_5594;
   wire n_1_737_5595;
   wire n_1_737_5597;
   wire n_1_737_5598;
   wire n_1_737_5599;
   wire n_1_737_5600;
   wire n_1_737_5601;
   wire n_1_737_5603;
   wire n_1_737_5604;
   wire n_1_737_5605;
   wire n_1_737_5606;
   wire n_1_737_5607;
   wire n_1_737_5608;
   wire n_1_737_5609;
   wire n_1_737_5610;
   wire n_1_737_5611;
   wire n_1_737_5612;
   wire n_1_737_5613;
   wire n_1_737_5614;
   wire n_1_737_5615;
   wire n_1_737_5616;
   wire n_1_737_5617;
   wire n_1_737_5618;
   wire n_1_737_5619;
   wire n_1_737_5620;
   wire n_1_737_5621;
   wire n_1_737_5622;
   wire n_1_737_5623;
   wire n_1_737_5624;
   wire n_1_737_5625;
   wire n_1_737_5626;
   wire n_1_737_5627;
   wire n_1_737_5628;
   wire n_1_737_5629;
   wire n_1_737_5630;
   wire n_1_737_5631;
   wire n_1_737_5632;
   wire n_1_737_5633;
   wire n_1_737_5634;
   wire n_1_737_5635;
   wire n_1_737_5636;
   wire n_1_737_5637;
   wire n_1_737_5638;
   wire n_1_737_5639;
   wire n_1_737_5640;
   wire n_1_737_5641;
   wire n_1_737_5642;
   wire n_1_737_5643;
   wire n_1_737_5644;
   wire n_1_737_5645;
   wire n_1_737_5646;
   wire n_1_737_5647;
   wire n_1_737_5648;
   wire n_1_737_5649;
   wire n_1_737_5650;
   wire n_1_737_5651;
   wire n_1_737_5652;
   wire n_1_737_5653;
   wire n_1_737_5654;
   wire n_1_737_5655;
   wire n_1_737_5656;
   wire n_1_737_5657;
   wire n_1_737_5658;
   wire n_1_737_5659;
   wire n_1_737_5660;
   wire n_1_737_5661;
   wire n_1_737_5662;
   wire n_1_737_5663;
   wire n_1_737_5664;
   wire n_1_737_5665;
   wire n_1_737_5666;
   wire n_1_737_5667;
   wire n_1_737_5668;
   wire n_1_737_5669;
   wire n_1_737_5670;
   wire n_1_737_5671;
   wire n_1_737_5672;
   wire n_1_737_5673;
   wire n_1_737_5674;
   wire n_1_737_5675;
   wire n_1_737_5676;
   wire n_1_737_5677;
   wire n_1_737_5678;
   wire n_1_737_5679;
   wire n_1_737_5680;
   wire n_1_737_1870;
   wire n_1_737_1871;
   wire n_1_737_1874;
   wire n_1_737_1875;
   wire n_1_737_4402;
   wire n_1_737_5181;
   wire n_1_737_5596;
   wire n_1_737_1973;
   wire n_1_737_1969;
   wire n_1_737_1979;
   wire n_1_737_4400;
   wire n_1_737_5681;
   wire n_1_737_1970;
   wire n_1_737_5682;
   wire n_1_737_5683;
   wire n_1_737_5684;
   wire n_1_737_5685;
   wire n_1_737_5686;
   wire n_1_737_5687;
   wire n_1_737_5688;
   wire n_1_737_5689;
   wire n_1_737_5690;
   wire n_1_737_5691;
   wire n_1_737_5692;
   wire n_1_737_5693;
   wire n_1_737_5694;
   wire n_1_737_5695;
   wire n_1_737_5696;
   wire n_1_737_5697;
   wire n_1_737_5698;
   wire n_1_737_5699;
   wire n_1_737_1971;
   wire n_1_737_5700;
   wire n_1_737_5701;
   wire n_1_737_5702;
   wire n_1_737_5703;
   wire n_1_737_5704;
   wire n_1_737_5705;
   wire n_1_737_5706;
   wire n_1_737_5182;
   wire n_1_737_4401;
   wire n_1_737_4404;
   wire n_1_737_3110;
   wire n_1_737_4092;
   wire n_1_737_5602;
   wire n_1_737_4965;
   wire n_1_737_5167;
   wire n_1_737_4453;
   wire n_1_737_1978;
   wire n_1_737_1976;
   wire n_1_737_5337;
   wire n_4_1_0;
   wire n_4_1_1;
   wire n_4_513_0;
   wire n_4_513_1;
   wire n_4_513_2;
   wire n_4_513_3;
   wire n_4_0;
   wire n_4_54_0;
   wire n_4_54_1;
   wire n_4_1;
   wire n_4_2;
   wire n_4_3;
   wire n_0_2;
   wire n_0_129;
   wire n_0_390;
   wire n_0_5;
   wire n_0_0;
   wire n_0_711;
   wire n_0_701;
   wire n_0_688;
   wire n_0_683;
   wire n_0_677;
   wire n_0_672;
   wire n_0_667;
   wire n_0_657;
   wire n_0_651;
   wire n_0_645;
   wire n_0_639;
   wire n_0_633;
   wire n_0_627;
   wire n_0_621;
   wire n_0_615;
   wire n_0_609;
   wire n_0_603;
   wire n_0_597;
   wire n_0_592;
   wire n_0_586;
   wire n_0_580;
   wire n_0_574;
   wire n_0_568;
   wire n_0_562;
   wire n_0_556;
   wire n_0_550;
   wire n_0_545;
   wire n_0_541;
   wire n_0_535;
   wire n_0_529;
   wire n_0_523;
   wire n_0_517;
   wire n_0_511;
   wire n_0_505;
   wire n_0_499;
   wire n_0_493;
   wire n_0_487;
   wire n_0_481;
   wire n_0_475;
   wire n_0_469;
   wire n_0_463;
   wire n_0_457;
   wire n_0_452;
   wire n_0_449;
   wire n_0_443;
   wire n_0_437;
   wire n_0_432;
   wire n_0_426;
   wire n_0_420;
   wire n_0_414;
   wire n_0_408;
   wire n_0_403;
   wire n_0_708;
   wire n_0_680;
   wire n_0_648;
   wire n_0_636;
   wire n_0_624;
   wire n_0_612;
   wire n_0_600;
   wire n_0_589;
   wire n_0_577;
   wire n_0_565;
   wire n_0_553;
   wire n_0_544;
   wire n_0_532;
   wire n_0_520;
   wire n_0_508;
   wire n_0_496;
   wire n_0_484;
   wire n_0_472;
   wire n_0_460;
   wire n_0_440;
   wire n_0_429;
   wire n_0_417;
   wire n_0_411;
   wire n_0_405;
   wire n_0_400;
   wire n_0_392;
   wire n_0_654;
   wire n_0_630;
   wire n_0_606;
   wire n_0_583;
   wire n_0_559;
   wire n_0_538;
   wire n_0_514;
   wire n_0_490;
   wire n_0_466;
   wire n_0_446;
   wire n_0_423;
   wire n_0_397;
   wire n_0_664;
   wire n_0_618;
   wire n_0_571;
   wire n_0_526;
   wire n_0_478;
   wire n_0_404;
   wire n_0_502;
   wire n_0_642;
   wire n_0_1;
   wire n_0_128;
   wire n_0_106_0;
   wire n_0_106_1;
   wire n_0_106_2;
   wire n_0_131;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_145;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_157;
   wire n_0_162;
   wire n_0_168;
   wire n_0_169;
   wire n_0_171;
   wire n_0_172;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_177;
   wire n_0_178;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_190;
   wire n_0_192;
   wire n_0_193;
   wire n_0_194;
   wire n_0_199;
   wire n_0_203;
   wire n_0_206;
   wire n_0_209;
   wire n_0_210;
   wire n_0_211;
   wire n_0_212;
   wire n_0_213;
   wire n_0_214;
   wire n_0_215;
   wire n_0_216;
   wire n_0_218;
   wire n_0_219;
   wire n_0_220;
   wire n_0_227;
   wire n_0_230;
   wire n_0_233;
   wire n_0_234;
   wire n_0_236;
   wire n_0_239;
   wire n_0_243;
   wire n_0_244;
   wire n_0_245;
   wire n_0_246;
   wire n_0_247;
   wire n_0_249;
   wire n_0_255;
   wire n_0_143;
   wire n_0_107_0;
   wire n_0_107_1;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_144;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_152;
   wire n_0_156;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_166;
   wire n_0_167;
   wire n_0_170;
   wire n_0_179;
   wire n_0_180;
   wire n_0_181;
   wire n_0_191;
   wire n_0_195;
   wire n_0_196;
   wire n_0_197;
   wire n_0_198;
   wire n_0_200;
   wire n_0_201;
   wire n_0_202;
   wire n_0_204;
   wire n_0_205;
   wire n_0_207;
   wire n_0_208;
   wire n_0_217;
   wire n_0_221;
   wire n_0_222;
   wire n_0_223;
   wire n_0_224;
   wire n_0_225;
   wire n_0_226;
   wire n_0_228;
   wire n_0_229;
   wire n_0_231;
   wire n_0_232;
   wire n_0_235;
   wire n_0_237;
   wire n_0_238;
   wire n_0_240;
   wire n_0_241;
   wire n_0_242;
   wire n_0_248;
   wire n_0_250;
   wire n_0_251;
   wire n_0_252;
   wire n_0_253;
   wire n_0_254;
   wire n_0_256;
   wire n_0_257;
   wire n_0_258;
   wire n_0_259;
   wire n_0_108_0;
   wire n_0_108_1;
   wire n_0_108_2;
   wire n_0_260;
   wire n_0_130;
   wire n_0_395;
   wire n_0_112_0;
   wire n_0_112_1;
   wire n_0_261;
   wire n_0_3;
   wire n_0_712;
   wire n_0_4;
   wire n_0_702;
   wire n_0_6;
   wire n_0_689;
   wire n_0_7;
   wire n_0_684;
   wire n_0_8;
   wire n_0_678;
   wire n_0_9;
   wire n_0_673;
   wire n_0_10;
   wire n_0_668;
   wire n_0_11;
   wire n_0_658;
   wire n_0_12;
   wire n_0_652;
   wire n_0_13;
   wire n_0_646;
   wire n_0_14;
   wire n_0_640;
   wire n_0_15;
   wire n_0_634;
   wire n_0_16;
   wire n_0_628;
   wire n_0_17;
   wire n_0_622;
   wire n_0_18;
   wire n_0_616;
   wire n_0_19;
   wire n_0_610;
   wire n_0_20;
   wire n_0_604;
   wire n_0_21;
   wire n_0_598;
   wire n_0_22;
   wire n_0_593;
   wire n_0_23;
   wire n_0_587;
   wire n_0_24;
   wire n_0_581;
   wire n_0_25;
   wire n_0_575;
   wire n_0_26;
   wire n_0_569;
   wire n_0_27;
   wire n_0_563;
   wire n_0_28;
   wire n_0_557;
   wire n_0_29;
   wire n_0_551;
   wire n_0_30;
   wire n_0_546;
   wire n_0_31;
   wire n_0_542;
   wire n_0_32;
   wire n_0_536;
   wire n_0_33;
   wire n_0_530;
   wire n_0_34;
   wire n_0_524;
   wire n_0_35;
   wire n_0_518;
   wire n_0_36;
   wire n_0_512;
   wire n_0_37;
   wire n_0_506;
   wire n_0_38;
   wire n_0_500;
   wire n_0_39;
   wire n_0_494;
   wire n_0_40;
   wire n_0_488;
   wire n_0_41;
   wire n_0_482;
   wire n_0_42;
   wire n_0_476;
   wire n_0_43;
   wire n_0_470;
   wire n_0_44;
   wire n_0_464;
   wire n_0_194_0;
   wire n_0_194_1;
   wire n_0_45;
   wire n_0_458;
   wire n_0_196_0;
   wire n_0_196_1;
   wire n_0_46;
   wire n_0_453;
   wire n_0_47;
   wire n_0_450;
   wire n_0_48;
   wire n_0_444;
   wire n_0_49;
   wire n_0_438;
   wire n_0_50;
   wire n_0_433;
   wire n_0_51;
   wire n_0_427;
   wire n_0_52;
   wire n_0_421;
   wire n_0_53;
   wire n_0_415;
   wire n_0_54;
   wire n_0_409;
   wire n_0_214_0;
   wire n_0_214_1;
   wire n_0_55;
   wire n_0_709;
   wire n_0_56;
   wire n_0_681;
   wire n_0_57;
   wire n_0_649;
   wire n_0_58;
   wire n_0_637;
   wire n_0_59;
   wire n_0_625;
   wire n_0_60;
   wire n_0_613;
   wire n_0_61;
   wire n_0_601;
   wire n_0_62;
   wire n_0_590;
   wire n_0_63;
   wire n_0_578;
   wire n_0_64;
   wire n_0_566;
   wire n_0_65;
   wire n_0_554;
   wire n_0_66;
   wire n_0_533;
   wire n_0_67;
   wire n_0_521;
   wire n_0_68;
   wire n_0_509;
   wire n_0_69;
   wire n_0_497;
   wire n_0_70;
   wire n_0_485;
   wire n_0_71;
   wire n_0_473;
   wire n_0_72;
   wire n_0_461;
   wire n_0_252_0;
   wire n_0_252_1;
   wire n_0_73;
   wire n_0_441;
   wire n_0_74;
   wire n_0_430;
   wire n_0_75;
   wire n_0_418;
   wire n_0_76;
   wire n_0_412;
   wire n_0_77;
   wire n_0_406;
   wire n_0_262_0;
   wire n_0_262_1;
   wire n_0_78;
   wire n_0_401;
   wire n_0_79;
   wire n_0_393;
   wire n_0_80;
   wire n_0_655;
   wire n_0_81;
   wire n_0_631;
   wire n_0_82;
   wire n_0_607;
   wire n_0_83;
   wire n_0_584;
   wire n_0_84;
   wire n_0_560;
   wire n_0_85;
   wire n_0_539;
   wire n_0_278_0;
   wire n_0_278_1;
   wire n_0_86;
   wire n_0_515;
   wire n_0_87;
   wire n_0_491;
   wire n_0_88;
   wire n_0_467;
   wire n_0_284_0;
   wire n_0_284_1;
   wire n_0_89;
   wire n_0_447;
   wire n_0_90;
   wire n_0_424;
   wire n_0_91;
   wire n_0_92;
   wire n_0_398;
   wire n_0_93;
   wire n_0_665;
   wire n_0_94;
   wire n_0_619;
   wire n_0_95;
   wire n_0_572;
   wire n_0_96;
   wire n_0_527;
   wire n_0_97;
   wire n_0_479;
   wire n_0_435;
   wire n_0_98;
   wire n_0_503;
   wire n_0_305_0;
   wire n_0_305_1;
   wire n_0_99;
   wire n_0_643;
   wire n_0_308_0;
   wire n_0_308_1;
   wire n_0_262;
   wire n_0_263;
   wire n_0_309_0;
   wire n_0_309_1;
   wire n_0_264;
   wire n_0_310_0;
   wire n_0_310_1;
   wire n_0_310_2;
   wire n_0_265;
   wire n_0_311_0;
   wire n_0_311_1;
   wire n_0_311_2;
   wire n_0_266;
   wire n_0_312_0;
   wire n_0_312_1;
   wire n_0_312_2;
   wire n_0_267;
   wire n_0_313_0;
   wire n_0_313_1;
   wire n_0_313_2;
   wire n_0_268;
   wire n_0_314_0;
   wire n_0_314_1;
   wire n_0_314_2;
   wire n_0_269;
   wire n_0_315_0;
   wire n_0_315_1;
   wire n_0_270;
   wire n_0_316_0;
   wire n_0_316_1;
   wire n_0_271;
   wire n_0_317_0;
   wire n_0_317_1;
   wire n_0_317_2;
   wire n_0_272;
   wire n_0_318_0;
   wire n_0_318_1;
   wire n_0_318_2;
   wire n_0_273;
   wire n_0_319_0;
   wire n_0_319_1;
   wire n_0_319_2;
   wire n_0_274;
   wire n_0_320_0;
   wire n_0_320_1;
   wire n_0_320_2;
   wire n_0_275;
   wire n_0_321_0;
   wire n_0_321_1;
   wire n_0_321_2;
   wire n_0_276;
   wire n_0_322_0;
   wire n_0_322_1;
   wire n_0_322_2;
   wire n_0_277;
   wire n_0_323_0;
   wire n_0_323_1;
   wire n_0_323_2;
   wire n_0_278;
   wire n_0_324_0;
   wire n_0_324_1;
   wire n_0_324_2;
   wire n_0_279;
   wire n_0_325_0;
   wire n_0_325_1;
   wire n_0_325_2;
   wire n_0_280;
   wire n_0_326_0;
   wire n_0_326_1;
   wire n_0_281;
   wire n_0_327_0;
   wire n_0_327_1;
   wire n_0_327_2;
   wire n_0_282;
   wire n_0_328_0;
   wire n_0_328_1;
   wire n_0_328_2;
   wire n_0_283;
   wire n_0_329_0;
   wire n_0_329_1;
   wire n_0_284;
   wire n_0_330_0;
   wire n_0_330_1;
   wire n_0_330_2;
   wire n_0_285;
   wire n_0_331_0;
   wire n_0_331_1;
   wire n_0_331_2;
   wire n_0_286;
   wire n_0_332_0;
   wire n_0_332_1;
   wire n_0_332_2;
   wire n_0_287;
   wire n_0_333_0;
   wire n_0_333_1;
   wire n_0_288;
   wire n_0_334_0;
   wire n_0_334_1;
   wire n_0_289;
   wire n_0_335_0;
   wire n_0_335_1;
   wire n_0_290;
   wire n_0_336_0;
   wire n_0_336_1;
   wire n_0_291;
   wire n_0_337_0;
   wire n_0_337_1;
   wire n_0_337_2;
   wire n_0_292;
   wire n_0_338_0;
   wire n_0_338_1;
   wire n_0_338_2;
   wire n_0_293;
   wire n_0_339_0;
   wire n_0_339_1;
   wire n_0_340_0;
   wire n_0_340_1;
   wire n_0_294;
   wire n_0_341_0;
   wire n_0_341_1;
   wire n_0_295;
   wire n_0_342_0;
   wire n_0_342_1;
   wire n_0_296;
   wire n_0_343_0;
   wire n_0_343_1;
   wire n_0_297;
   wire n_0_298;
   wire n_0_344_0;
   wire n_0_344_1;
   wire n_0_344_2;
   wire n_0_345_0;
   wire n_0_345_1;
   wire n_0_299;
   wire n_0_346_0;
   wire n_0_346_1;
   wire n_0_300;
   wire n_0_347_0;
   wire n_0_347_1;
   wire n_0_301;
   wire n_0_302;
   wire n_0_348_0;
   wire n_0_348_1;
   wire n_0_303;
   wire n_0_349_0;
   wire n_0_349_1;
   wire n_0_349_2;
   wire n_0_304;
   wire n_0_350_0;
   wire n_0_350_1;
   wire n_0_350_2;
   wire n_0_305;
   wire n_0_351_0;
   wire n_0_351_1;
   wire n_0_351_2;
   wire n_0_352_0;
   wire n_0_352_1;
   wire n_0_306;
   wire n_0_353_0;
   wire n_0_353_1;
   wire n_0_307;
   wire n_0_308;
   wire n_0_354_0;
   wire n_0_354_1;
   wire n_0_354_2;
   wire n_0_355_0;
   wire n_0_355_1;
   wire n_0_309;
   wire n_0_356_0;
   wire n_0_356_1;
   wire n_0_310;
   wire n_0_311;
   wire n_0_357_0;
   wire n_0_357_1;
   wire n_0_357_2;
   wire n_0_358_0;
   wire n_0_358_1;
   wire n_0_312;
   wire n_0_313;
   wire n_0_359_0;
   wire n_0_359_1;
   wire n_0_359_2;
   wire n_0_314;
   wire n_0_360_0;
   wire n_0_360_1;
   wire n_0_315;
   wire n_0_361_0;
   wire n_0_361_1;
   wire n_0_361_2;
   wire n_0_316;
   wire n_0_362_0;
   wire n_0_362_1;
   wire n_0_362_2;
   wire n_0_317;
   wire n_0_363_0;
   wire n_0_363_1;
   wire n_0_363_2;
   wire n_0_318;
   wire n_0_364_0;
   wire n_0_364_1;
   wire n_0_364_2;
   wire n_0_365_0;
   wire n_0_365_1;
   wire n_0_319;
   wire n_0_320;
   wire n_0_366_0;
   wire n_0_366_1;
   wire n_0_366_2;
   wire n_0_367_0;
   wire n_0_367_1;
   wire n_0_321;
   wire n_0_322;
   wire n_0_368_0;
   wire n_0_368_1;
   wire n_0_368_2;
   wire n_0_369_0;
   wire n_0_369_1;
   wire n_0_323;
   wire n_0_370_0;
   wire n_0_370_1;
   wire n_0_324;
   wire n_0_371_0;
   wire n_0_371_1;
   wire n_0_325;
   wire n_0_372_0;
   wire n_0_372_1;
   wire n_0_326;
   wire n_0_373_0;
   wire n_0_373_1;
   wire n_0_327;
   wire n_0_374_0;
   wire n_0_374_1;
   wire n_0_328;
   wire n_0_375_0;
   wire n_0_375_1;
   wire n_0_329;
   wire n_0_330;
   wire n_0_376_0;
   wire n_0_376_1;
   wire n_0_376_2;
   wire n_0_377_0;
   wire n_0_377_1;
   wire n_0_331;
   wire n_0_332;
   wire n_0_378_0;
   wire n_0_378_1;
   wire n_0_378_2;
   wire n_0_333;
   wire n_0_379_0;
   wire n_0_379_1;
   wire n_0_379_2;
   wire n_0_334;
   wire n_0_380_0;
   wire n_0_380_1;
   wire n_0_335;
   wire n_0_381_0;
   wire n_0_381_1;
   wire n_0_381_2;
   wire n_0_382_0;
   wire n_0_382_1;
   wire n_0_336;
   wire n_0_337;
   wire n_0_383_0;
   wire n_0_383_1;
   wire n_0_383_2;
   wire n_0_338;
   wire n_0_384_0;
   wire n_0_384_1;
   wire n_0_384_2;
   wire n_0_339;
   wire n_0_385_0;
   wire n_0_385_1;
   wire n_0_385_2;
   wire n_0_386_0;
   wire n_0_386_1;
   wire n_0_340;
   wire n_0_341;
   wire n_0_387_0;
   wire n_0_387_1;
   wire n_0_387_2;
   wire n_0_388_0;
   wire n_0_388_1;
   wire n_0_342;
   wire n_0_343;
   wire n_0_389_0;
   wire n_0_389_1;
   wire n_0_389_2;
   wire n_0_344;
   wire n_0_390_0;
   wire n_0_390_1;
   wire n_0_390_2;
   wire n_0_345;
   wire n_0_391_0;
   wire n_0_391_1;
   wire n_0_346;
   wire n_0_392_0;
   wire n_0_392_1;
   wire n_0_392_2;
   wire n_0_347;
   wire n_0_393_0;
   wire n_0_393_1;
   wire n_0_393_2;
   wire n_0_348;
   wire n_0_394_0;
   wire n_0_394_1;
   wire n_0_394_2;
   wire n_0_349;
   wire n_0_395_0;
   wire n_0_395_1;
   wire n_0_395_2;
   wire n_0_396_0;
   wire n_0_396_1;
   wire n_0_350;
   wire n_0_351;
   wire n_0_397_0;
   wire n_0_397_1;
   wire n_0_397_2;
   wire n_0_352;
   wire n_0_398_0;
   wire n_0_398_1;
   wire n_0_398_2;
   wire n_0_353;
   wire n_0_399_0;
   wire n_0_399_1;
   wire n_0_399_2;
   wire n_0_354;
   wire n_0_400_0;
   wire n_0_400_1;
   wire n_0_400_2;
   wire n_0_401_0;
   wire n_0_401_1;
   wire n_0_355;
   wire n_0_356;
   wire n_0_402_0;
   wire n_0_402_1;
   wire n_0_402_2;
   wire n_0_357;
   wire n_0_403_0;
   wire n_0_403_1;
   wire n_0_403_2;
   wire n_0_358;
   wire n_0_404_0;
   wire n_0_404_1;
   wire n_0_404_2;
   wire n_0_359;
   wire n_0_405_0;
   wire n_0_405_1;
   wire n_0_405_2;
   wire n_0_360;
   wire n_0_406_0;
   wire n_0_406_1;
   wire n_0_406_2;
   wire n_0_361;
   wire n_0_407_0;
   wire n_0_407_1;
   wire n_0_407_2;
   wire n_0_362;
   wire n_0_408_0;
   wire n_0_408_1;
   wire n_0_408_2;
   wire n_0_363;
   wire n_0_409_0;
   wire n_0_409_1;
   wire n_0_409_2;
   wire n_0_364;
   wire n_0_410_0;
   wire n_0_410_1;
   wire n_0_410_2;
   wire n_0_365;
   wire n_0_411_0;
   wire n_0_411_1;
   wire n_0_411_2;
   wire n_0_366;
   wire n_0_412_0;
   wire n_0_412_1;
   wire n_0_412_2;
   wire n_0_367;
   wire n_0_413_0;
   wire n_0_413_1;
   wire n_0_413_2;
   wire n_0_368;
   wire n_0_414_0;
   wire n_0_414_1;
   wire n_0_414_2;
   wire n_0_369;
   wire n_0_415_0;
   wire n_0_415_1;
   wire n_0_415_2;
   wire n_0_370;
   wire n_0_416_0;
   wire n_0_416_1;
   wire n_0_416_2;
   wire n_0_371;
   wire n_0_417_0;
   wire n_0_417_1;
   wire n_0_372;
   wire n_0_418_0;
   wire n_0_418_1;
   wire n_0_418_2;
   wire n_0_373;
   wire n_0_419_0;
   wire n_0_419_1;
   wire n_0_419_2;
   wire n_0_420_0;
   wire n_0_420_1;
   wire n_0_374;
   wire n_0_421_0;
   wire n_0_421_1;
   wire n_0_375;
   wire n_0_376;
   wire n_0_422_0;
   wire n_0_422_1;
   wire n_0_422_2;
   wire n_0_377;
   wire n_0_423_0;
   wire n_0_423_1;
   wire n_0_423_2;
   wire n_0_378;
   wire n_0_424_0;
   wire n_0_424_1;
   wire n_0_424_2;
   wire n_0_379;
   wire n_0_425_0;
   wire n_0_425_1;
   wire n_0_425_2;
   wire n_0_380;
   wire n_0_426_0;
   wire n_0_426_1;
   wire n_0_426_2;
   wire n_0_381;
   wire n_0_427_0;
   wire n_0_427_1;
   wire n_0_427_2;
   wire n_0_382;
   wire n_0_428_0;
   wire n_0_428_1;
   wire n_0_428_2;
   wire n_0_429_0;
   wire n_0_429_1;
   wire n_0_383;
   wire n_0_384;
   wire n_0_430_0;
   wire n_0_430_1;
   wire n_0_430_2;
   wire n_0_385;
   wire n_0_431_0;
   wire n_0_431_1;
   wire n_0_386;
   wire n_0_432_0;
   wire n_0_432_1;
   wire n_0_432_2;
   wire n_0_387;
   wire n_0_433_0;
   wire n_0_433_1;
   wire n_0_433_2;
   wire n_0_388;
   wire n_0_434_0;
   wire n_0_434_1;
   wire n_0_434_2;
   wire n_0_435_0;
   wire n_0_435_1;
   wire n_0_389;
   wire n_0_436_0;
   wire n_0_436_1;
   wire n_0_391;
   wire n_0_394;
   wire n_0_437_0;
   wire n_0_437_1;
   wire n_0_437_2;
   wire n_0_438_0;
   wire n_0_438_1;
   wire n_0_396;
   wire n_0_399;
   wire n_0_439_0;
   wire n_0_439_1;
   wire n_0_439_2;
   wire n_0_440_0;
   wire n_0_440_1;
   wire n_0_402;
   wire n_0_407;
   wire n_0_441_0;
   wire n_0_441_1;
   wire n_0_441_2;
   wire n_0_442_0;
   wire n_0_442_1;
   wire n_0_410;
   wire n_0_413;
   wire n_0_443_0;
   wire n_0_443_1;
   wire n_0_416;
   wire n_0_444_0;
   wire n_0_444_1;
   wire n_0_419;
   wire n_0_445_0;
   wire n_0_445_1;
   wire n_0_422;
   wire n_0_446_0;
   wire n_0_446_1;
   wire n_0_447_0;
   wire n_0_447_1;
   wire n_0_425;
   wire n_0_428;
   wire n_0_448_0;
   wire n_0_448_1;
   wire n_0_448_2;
   wire n_0_449_0;
   wire n_0_449_1;
   wire n_0_431;
   wire n_0_450_0;
   wire n_0_450_1;
   wire n_0_434;
   wire n_0_451_0;
   wire n_0_451_1;
   wire n_0_436;
   wire n_0_452_0;
   wire n_0_452_1;
   wire n_0_439;
   wire n_0_453_0;
   wire n_0_453_1;
   wire n_0_442;
   wire n_0_454_0;
   wire n_0_454_1;
   wire n_0_445;
   wire n_0_455_0;
   wire n_0_455_1;
   wire n_0_448;
   wire n_0_456_0;
   wire n_0_456_1;
   wire n_0_451;
   wire n_0_457_0;
   wire n_0_457_1;
   wire n_0_454;
   wire n_0_458_0;
   wire n_0_458_1;
   wire n_0_455;
   wire n_0_459_0;
   wire n_0_459_1;
   wire n_0_456;
   wire n_0_460_0;
   wire n_0_460_1;
   wire n_0_459;
   wire n_0_461_0;
   wire n_0_461_1;
   wire n_0_462;
   wire n_0_462_0;
   wire n_0_462_1;
   wire n_0_465;
   wire n_0_468;
   wire n_0_463_0;
   wire n_0_463_1;
   wire n_0_464_0;
   wire n_0_464_1;
   wire n_0_471;
   wire n_0_474;
   wire n_0_465_0;
   wire n_0_465_1;
   wire n_0_465_2;
   wire n_0_477;
   wire n_0_466_0;
   wire n_0_466_1;
   wire n_0_466_2;
   wire n_0_480;
   wire n_0_467_0;
   wire n_0_467_1;
   wire n_0_467_2;
   wire n_0_483;
   wire n_0_468_0;
   wire n_0_468_1;
   wire n_0_468_2;
   wire n_0_486;
   wire n_0_469_0;
   wire n_0_469_1;
   wire n_0_469_2;
   wire n_0_489;
   wire n_0_470_0;
   wire n_0_470_1;
   wire n_0_470_2;
   wire n_0_471_0;
   wire n_0_471_1;
   wire n_0_492;
   wire n_0_472_0;
   wire n_0_472_1;
   wire n_0_495;
   wire n_0_473_0;
   wire n_0_473_1;
   wire n_0_498;
   wire n_0_474_0;
   wire n_0_474_1;
   wire n_0_501;
   wire n_0_504;
   wire n_0_475_0;
   wire n_0_475_1;
   wire n_0_475_2;
   wire n_0_476_0;
   wire n_0_476_1;
   wire n_0_507;
   wire n_0_477_0;
   wire n_0_477_1;
   wire n_0_510;
   wire n_0_513;
   wire n_0_478_0;
   wire n_0_478_1;
   wire n_0_478_2;
   wire n_0_479_0;
   wire n_0_479_1;
   wire n_0_516;
   wire n_0_480_0;
   wire n_0_480_1;
   wire n_0_519;
   wire n_0_481_0;
   wire n_0_481_1;
   wire n_0_522;
   wire n_0_525;
   wire n_0_482_0;
   wire n_0_482_1;
   wire n_0_482_2;
   wire n_0_483_0;
   wire n_0_483_1;
   wire n_0_528;
   wire n_0_484_0;
   wire n_0_484_1;
   wire n_0_531;
   wire n_0_534;
   wire n_0_485_0;
   wire n_0_485_1;
   wire n_0_485_2;
   wire n_0_486_0;
   wire n_0_486_1;
   wire n_0_537;
   wire n_0_540;
   wire n_0_487_0;
   wire n_0_487_1;
   wire n_0_487_2;
   wire n_0_488_0;
   wire n_0_488_1;
   wire n_0_543;
   wire n_0_489_0;
   wire n_0_489_1;
   wire n_0_547;
   wire n_0_548;
   wire n_0_490_0;
   wire n_0_490_1;
   wire n_0_490_2;
   wire n_0_491_0;
   wire n_0_491_1;
   wire n_0_549;
   wire n_0_552;
   wire n_0_492_0;
   wire n_0_492_1;
   wire n_0_492_2;
   wire n_0_555;
   wire n_0_493_0;
   wire n_0_493_1;
   wire n_0_493_2;
   wire n_0_558;
   wire n_0_494_0;
   wire n_0_494_1;
   wire n_0_494_2;
   wire n_0_495_0;
   wire n_0_495_1;
   wire n_0_561;
   wire n_0_564;
   wire n_0_496_0;
   wire n_0_496_1;
   wire n_0_496_2;
   wire n_0_567;
   wire n_0_497_0;
   wire n_0_497_1;
   wire n_0_497_2;
   wire n_0_570;
   wire n_0_498_0;
   wire n_0_498_1;
   wire n_0_498_2;
   wire n_0_573;
   wire n_0_499_0;
   wire n_0_499_1;
   wire n_0_499_2;
   wire n_0_576;
   wire n_0_500_0;
   wire n_0_500_1;
   wire n_0_500_2;
   wire n_0_579;
   wire n_0_501_0;
   wire n_0_501_1;
   wire n_0_501_2;
   wire n_0_582;
   wire n_0_502_0;
   wire n_0_502_1;
   wire n_0_502_2;
   wire n_0_585;
   wire n_0_503_0;
   wire n_0_503_1;
   wire n_0_503_2;
   wire n_0_588;
   wire n_0_504_0;
   wire n_0_504_1;
   wire n_0_504_2;
   wire n_0_505_0;
   wire n_0_505_1;
   wire n_0_591;
   wire n_0_506_0;
   wire n_0_506_1;
   wire n_0_594;
   wire n_0_507_0;
   wire n_0_507_1;
   wire n_0_595;
   wire n_0_596;
   wire n_0_508_0;
   wire n_0_508_1;
   wire n_0_508_2;
   wire n_0_599;
   wire n_0_509_0;
   wire n_0_509_1;
   wire n_0_509_2;
   wire n_0_602;
   wire n_0_511_0;
   wire n_0_511_1;
   wire n_0_605;
   wire n_0_512_0;
   wire n_0_512_1;
   wire n_0_512_2;
   wire n_0_608;
   wire n_0_513_0;
   wire n_0_513_1;
   wire n_0_513_2;
   wire n_0_611;
   wire n_0_514_0;
   wire n_0_514_1;
   wire n_0_514_2;
   wire n_0_614;
   wire n_0_515_0;
   wire n_0_515_1;
   wire n_0_515_2;
   wire n_0_617;
   wire n_0_516_0;
   wire n_0_516_1;
   wire n_0_516_2;
   wire n_0_620;
   wire n_0_517_0;
   wire n_0_517_1;
   wire n_0_517_2;
   wire n_0_623;
   wire n_0_518_0;
   wire n_0_518_1;
   wire n_0_518_2;
   wire n_0_519_0;
   wire n_0_519_1;
   wire n_0_626;
   wire n_0_520_0;
   wire n_0_520_1;
   wire n_0_629;
   wire n_0_521_0;
   wire n_0_521_1;
   wire n_0_632;
   wire n_0_635;
   wire n_0_522_0;
   wire n_0_522_1;
   wire n_0_522_2;
   wire n_0_523_0;
   wire n_0_523_1;
   wire n_0_638;
   wire n_0_641;
   wire n_0_524_0;
   wire n_0_524_1;
   wire n_0_524_2;
   wire n_0_525_0;
   wire n_0_525_1;
   wire n_0_644;
   wire n_0_526_0;
   wire n_0_526_1;
   wire n_0_647;
   wire n_0_650;
   wire n_0_527_0;
   wire n_0_527_1;
   wire n_0_527_2;
   wire n_0_528_0;
   wire n_0_528_1;
   wire n_0_653;
   wire n_0_656;
   wire n_0_529_0;
   wire n_0_529_1;
   wire n_0_530_0;
   wire n_0_530_1;
   wire n_0_659;
   wire n_0_531_0;
   wire n_0_531_1;
   wire n_0_660;
   wire n_0_532_0;
   wire n_0_532_1;
   wire n_0_661;
   wire n_0_533_0;
   wire n_0_533_1;
   wire n_0_662;
   wire n_0_534_0;
   wire n_0_534_1;
   wire n_0_663;
   wire n_0_535_0;
   wire n_0_535_1;
   wire n_0_666;
   wire n_0_536_0;
   wire n_0_536_1;
   wire n_0_669;
   wire n_0_670;
   wire n_0_537_0;
   wire n_0_537_1;
   wire n_0_537_2;
   wire n_0_671;
   wire n_0_538_0;
   wire n_0_538_1;
   wire n_0_538_2;
   wire n_0_539_0;
   wire n_0_539_1;
   wire n_0_674;
   wire n_0_675;
   wire n_0_540_0;
   wire n_0_540_1;
   wire n_0_540_2;
   wire n_0_541_0;
   wire n_0_541_1;
   wire n_0_676;
   wire n_0_679;
   wire n_0_682;
   wire n_0_543_0;
   wire n_0_543_1;
   wire n_0_685;
   wire n_0_686;
   wire n_0_687;
   wire n_0_546_0;
   wire n_0_546_1;
   wire n_0_690;
   wire n_0_547_0;
   wire n_0_547_1;
   wire n_0_691;
   wire n_0_692;
   wire n_0_693;
   wire n_0_694;
   wire n_0_695;
   wire n_0_696;
   wire n_0_697;
   wire n_0_698;
   wire n_0_699;
   wire n_0_700;
   wire n_0_703;
   wire n_0_704;
   wire n_0_705;
   wire n_0_560_0;
   wire n_0_560_1;
   wire n_0_706;
   wire n_0_707;
   wire n_0_710;
   wire n_0_713;
   wire n_0_564_0;
   wire n_0_564_1;
   wire n_0_714;
   wire n_0_565_0;
   wire n_0_565_1;
   wire n_0_715;
   wire n_0_566_0;
   wire n_0_566_1;
   wire n_0_716;
   wire n_0_567_0;
   wire n_0_567_1;
   wire n_0_717;
   wire n_0_718;
   wire n_0_719;
   wire n_0_570_0;
   wire n_0_570_1;
   wire n_0_720;
   wire n_0_721;
   wire n_0_722;
   wire n_0_723;
   wire n_0_724;
   wire n_0_725;
   wire n_0_726;
   wire n_0_727;
   wire n_0_728;
   wire n_0_579_0;
   wire n_0_579_1;
   wire n_0_729;
   wire n_0_730;
   wire n_0_731;
   wire n_0_732;
   wire n_0_733;
   wire n_0_734;
   wire n_0_735;
   wire n_0_736;
   wire n_0_737;
   wire n_0_738;
   wire n_0_739;
   wire n_0_740;
   wire n_0_591_0;
   wire n_0_591_1;
   wire n_0_741;
   wire n_0_742;
   wire n_0_743;
   wire n_0_744;
   wire n_0_745;
   wire n_0_746;
   wire n_0_747;
   wire n_0_748;
   wire n_0_749;
   wire n_0_750;
   wire n_0_751;
   wire n_0_752;
   wire n_0_753;
   wire n_0_754;
   wire n_0_755;
   wire n_0_756;
   wire n_0_757;
   wire n_0_758;
   wire n_0_759;
   wire n_0_760;
   wire n_0_761;
   wire n_0_762;
   wire n_0_763;
   wire n_0_764;
   wire n_0_765;
   wire n_0_766;
   wire n_0_767;
   wire n_0_768;
   wire n_0_769;
   wire n_0_770;
   wire n_0_621_0;
   wire n_0_621_1;
   wire n_0_771;
   wire n_0_772;
   wire n_0_773;
   wire n_0_774;
   wire n_0_775;
   wire n_0_776;
   wire n_0_777;
   wire n_0_778;
   wire n_0_779;
   wire n_0_780;
   wire n_0_781;
   wire n_0_782;
   wire n_0_783;
   wire n_0_784;
   wire n_0_785;
   wire n_0_786;
   wire n_0_787;
   wire n_0_788;
   wire n_0_789;
   wire n_0_790;
   wire n_0_791;
   wire n_0_792;
   wire n_0_793;
   wire n_0_794;
   wire n_0_795;
   wire n_0_796;
   wire n_0_797;
   wire n_0_798;
   wire n_0_799;
   wire n_0_800;
   wire n_0_801;
   wire n_0_802;
   wire n_0_803;
   wire n_0_804;
   wire n_0_805;
   wire n_0_901;
   wire n_0_658_0;
   wire n_0_658_1;
   wire n_0_658_2;
   wire n_0_658_3;
   wire [6:0]\out_bs[7] ;
   wire [6:0]\out_as[7] ;
   wire n_0_806;
   wire n_0_100;
   wire n_0_680_0;
   wire n_0_680_1;
   wire n_0_680_2;
   wire n_0_680_3;
   wire n_0_101;
   wire n_0_681_0;
   wire n_0_681_1;
   wire n_0_681_2;
   wire n_0_681_3;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_697_0;
   wire n_0_118;
   wire n_0_807;
   wire n_0_699_0;
   wire n_0_699_1;
   wire n_0_808;
   wire n_0_700_0;
   wire n_0_700_1;
   wire n_0_700_2;
   wire n_0_809;
   wire n_0_701_0;
   wire n_0_701_1;
   wire n_0_810;
   wire n_0_702_0;
   wire n_0_702_1;
   wire n_0_811;
   wire n_0_703_0;
   wire n_0_703_1;
   wire n_0_812;
   wire n_0_704_0;
   wire n_0_704_1;
   wire n_0_813;
   wire n_0_705_0;
   wire n_0_705_1;
   wire n_0_705_2;
   wire n_0_814;
   wire n_0_706_0;
   wire n_0_706_1;
   wire n_0_706_2;
   wire n_0_815;
   wire n_0_707_0;
   wire n_0_707_1;
   wire n_0_119;
   wire n_0_708_0;
   wire n_0_708_1;
   wire n_0_708_2;
   wire n_0_708_3;
   wire n_0_709_0;
   wire n_0_709_1;
   wire n_0_709_2;
   wire n_0_709_3;
   wire n_0_710_0;
   wire n_0_710_1;
   wire n_0_710_2;
   wire n_0_710_3;
   wire n_0_711_0;
   wire n_0_711_1;
   wire n_0_711_2;
   wire n_0_711_3;
   wire n_0_712_0;
   wire n_0_712_1;
   wire n_0_712_2;
   wire n_0_712_3;
   wire n_0_713_0;
   wire n_0_713_1;
   wire n_0_713_2;
   wire n_0_713_3;
   wire n_0_714_0;
   wire n_0_714_1;
   wire n_0_714_2;
   wire n_0_714_3;
   wire n_0_900;
   wire n_0_715_0;
   wire n_0_715_1;
   wire n_0_715_2;
   wire n_0_715_3;
   wire n_0_899;
   wire n_0_716_0;
   wire n_0_716_1;
   wire n_0_716_2;
   wire n_0_716_3;
   wire n_0_898;
   wire n_0_717_0;
   wire n_0_717_1;
   wire n_0_717_2;
   wire n_0_717_3;
   wire n_0_897;
   wire n_0_718_0;
   wire n_0_718_1;
   wire n_0_718_2;
   wire n_0_718_3;
   wire n_0_896;
   wire n_0_719_0;
   wire n_0_719_1;
   wire n_0_719_2;
   wire n_0_719_3;
   wire n_0_720_0;
   wire n_0_720_1;
   wire n_0_720_2;
   wire n_0_720_3;
   wire n_0_895;
   wire n_0_721_0;
   wire n_0_721_1;
   wire n_0_721_2;
   wire n_0_721_3;
   wire n_0_120;
   wire n_0_722_0;
   wire n_0_722_1;
   wire n_0_722_2;
   wire n_0_722_3;
   wire n_0_121;
   wire n_0_723_0;
   wire n_0_723_1;
   wire n_0_723_2;
   wire n_0_723_3;
   wire n_0_122;
   wire n_0_724_0;
   wire n_0_724_1;
   wire n_0_724_2;
   wire n_0_724_3;
   wire n_0_123;
   wire n_0_725_0;
   wire n_0_725_1;
   wire n_0_725_2;
   wire n_0_725_3;
   wire n_0_124;
   wire n_0_726_0;
   wire n_0_726_1;
   wire n_0_726_2;
   wire n_0_726_3;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_657_0;
   wire n_0_657_1;
   wire n_0_657_2;
   wire n_0_657_3;
   wire n_0_848;
   wire n_0_657_4;
   wire n_0_657_5;
   wire n_0_657_6;
   wire n_0_657_7;
   wire n_0_657_8;
   wire n_0_657_9;
   wire n_0_657_10;
   wire n_0_657_11;
   wire n_0_657_12;
   wire n_0_657_13;
   wire n_0_657_14;
   wire n_0_657_15;
   wire n_0_657_16;
   wire n_0_657_17;
   wire n_0_657_18;
   wire n_0_657_19;
   wire n_0_657_20;
   wire n_0_657_21;
   wire n_0_879;
   wire n_0_657_22;
   wire n_0_657_23;
   wire n_0_657_24;
   wire n_0_657_25;
   wire n_0_657_26;
   wire n_0_657_27;
   wire n_0_911;
   wire n_0_657_28;
   wire n_0_657_29;
   wire n_0_657_30;
   wire n_0_657_31;
   wire n_0_657_32;
   wire n_0_657_33;
   wire n_0_920;
   wire n_0_657_34;
   wire n_0_657_35;
   wire n_0_657_36;
   wire n_0_657_37;
   wire n_0_657_38;
   wire n_0_657_39;
   wire n_0_922;
   wire n_0_657_40;
   wire n_0_657_41;
   wire n_0_657_42;
   wire n_0_657_43;
   wire n_0_657_44;
   wire n_0_657_45;
   wire n_0_934;
   wire n_0_657_46;
   wire n_0_657_47;
   wire n_0_657_48;
   wire n_0_657_49;
   wire n_0_657_50;
   wire n_0_657_51;
   wire n_0_657_52;
   wire n_0_657_53;
   wire n_0_657_54;
   wire n_0_657_55;
   wire n_0_939;
   wire n_0_657_56;
   wire n_0_657_57;
   wire n_0_657_58;
   wire n_0_657_59;
   wire n_0_657_60;
   wire n_0_657_61;
   wire n_0_941;
   wire n_0_657_62;
   wire n_0_657_63;
   wire n_0_657_64;
   wire n_0_657_65;
   wire n_0_657_66;
   wire n_0_657_67;
   wire n_0_945;
   wire n_0_657_68;
   wire n_0_657_69;
   wire n_0_657_70;
   wire n_0_657_71;
   wire n_0_657_72;
   wire n_0_657_73;
   wire n_0_657_74;
   wire n_0_657_75;
   wire n_0_950;
   wire n_0_657_76;
   wire n_0_657_77;
   wire n_0_657_78;
   wire n_0_657_79;
   wire n_0_657_80;
   wire n_0_816;
   wire n_0_657_81;
   wire n_0_657_82;
   wire n_0_657_83;
   wire n_0_657_84;
   wire n_0_657_85;
   wire n_0_657_86;
   wire n_0_657_87;
   wire n_0_817;
   wire n_0_657_88;
   wire n_0_657_89;
   wire n_0_657_90;
   wire n_0_657_91;
   wire n_0_657_92;
   wire n_0_657_93;
   wire n_0_657_94;
   wire n_0_818;
   wire n_0_657_95;
   wire n_0_657_96;
   wire n_0_657_97;
   wire n_0_657_98;
   wire n_0_657_99;
   wire n_0_657_100;
   wire n_0_657_101;
   wire n_0_819;
   wire n_0_657_102;
   wire n_0_657_103;
   wire n_0_657_104;
   wire n_0_657_105;
   wire n_0_657_106;
   wire n_0_657_107;
   wire n_0_657_108;
   wire n_0_820;
   wire n_0_657_109;
   wire n_0_657_110;
   wire n_0_657_111;
   wire n_0_657_112;
   wire n_0_657_113;
   wire n_0_657_114;
   wire n_0_657_115;
   wire n_0_821;
   wire n_0_657_116;
   wire n_0_657_117;
   wire n_0_657_118;
   wire n_0_657_119;
   wire n_0_657_120;
   wire n_0_657_121;
   wire n_0_822;
   wire n_0_657_122;
   wire n_0_657_123;
   wire n_0_657_124;
   wire n_0_657_125;
   wire n_0_657_126;
   wire n_0_657_127;
   wire n_0_657_128;
   wire n_0_823;
   wire n_0_657_129;
   wire n_0_657_130;
   wire n_0_657_131;
   wire n_0_657_132;
   wire n_0_657_133;
   wire n_0_657_134;
   wire n_0_657_135;
   wire n_0_824;
   wire n_0_657_136;
   wire n_0_657_137;
   wire n_0_657_138;
   wire n_0_657_139;
   wire n_0_657_140;
   wire n_0_657_141;
   wire n_0_657_142;
   wire n_0_825;
   wire n_0_657_143;
   wire n_0_657_144;
   wire n_0_657_145;
   wire n_0_657_146;
   wire n_0_657_147;
   wire n_0_657_148;
   wire n_0_657_149;
   wire n_0_657_150;
   wire n_0_826;
   wire n_0_657_151;
   wire n_0_657_152;
   wire n_0_657_153;
   wire n_0_657_154;
   wire n_0_657_155;
   wire n_0_657_156;
   wire n_0_657_157;
   wire n_0_827;
   wire n_0_657_158;
   wire n_0_657_159;
   wire n_0_657_160;
   wire n_0_657_161;
   wire n_0_657_162;
   wire n_0_657_163;
   wire n_0_657_164;
   wire n_0_828;
   wire n_0_657_165;
   wire n_0_657_166;
   wire n_0_657_167;
   wire n_0_657_168;
   wire n_0_657_169;
   wire n_0_657_170;
   wire n_0_657_171;
   wire n_0_657_172;
   wire n_0_829;
   wire n_0_657_173;
   wire n_0_657_174;
   wire n_0_657_175;
   wire n_0_657_176;
   wire n_0_657_177;
   wire n_0_657_178;
   wire n_0_657_179;
   wire n_0_830;
   wire n_0_657_180;
   wire n_0_657_181;
   wire n_0_657_182;
   wire n_0_657_183;
   wire n_0_657_184;
   wire n_0_657_185;
   wire n_0_657_186;
   wire n_0_831;
   wire n_0_657_187;
   wire n_0_657_188;
   wire n_0_657_189;
   wire n_0_657_190;
   wire n_0_657_191;
   wire n_0_657_192;
   wire n_0_657_193;
   wire n_0_832;
   wire n_0_657_194;
   wire n_0_657_195;
   wire n_0_657_196;
   wire n_0_657_197;
   wire n_0_657_198;
   wire n_0_657_199;
   wire n_0_657_200;
   wire n_0_833;
   wire n_0_657_201;
   wire n_0_657_202;
   wire n_0_657_203;
   wire n_0_657_204;
   wire n_0_657_205;
   wire n_0_657_206;
   wire n_0_657_207;
   wire n_0_834;
   wire n_0_657_208;
   wire n_0_657_209;
   wire n_0_657_210;
   wire n_0_657_211;
   wire n_0_657_212;
   wire n_0_657_213;
   wire n_0_657_214;
   wire n_0_835;
   wire n_0_657_215;
   wire n_0_657_216;
   wire n_0_657_217;
   wire n_0_657_218;
   wire n_0_657_219;
   wire n_0_657_220;
   wire n_0_657_221;
   wire n_0_836;
   wire n_0_657_222;
   wire n_0_657_223;
   wire n_0_657_224;
   wire n_0_657_225;
   wire n_0_657_226;
   wire n_0_657_227;
   wire n_0_657_228;
   wire n_0_837;
   wire n_0_657_229;
   wire n_0_657_230;
   wire n_0_657_231;
   wire n_0_657_232;
   wire n_0_657_233;
   wire n_0_657_234;
   wire n_0_657_235;
   wire n_0_838;
   wire n_0_657_236;
   wire n_0_657_237;
   wire n_0_657_238;
   wire n_0_657_239;
   wire n_0_657_240;
   wire n_0_657_241;
   wire n_0_657_242;
   wire n_0_839;
   wire n_0_657_243;
   wire n_0_657_244;
   wire n_0_657_245;
   wire n_0_657_246;
   wire n_0_657_247;
   wire n_0_657_248;
   wire n_0_657_249;
   wire n_0_840;
   wire n_0_657_250;
   wire n_0_657_251;
   wire n_0_657_252;
   wire n_0_657_253;
   wire n_0_657_254;
   wire n_0_657_255;
   wire n_0_657_256;
   wire n_0_841;
   wire n_0_657_257;
   wire n_0_657_258;
   wire n_0_657_259;
   wire n_0_657_260;
   wire n_0_657_261;
   wire n_0_657_262;
   wire n_0_657_263;
   wire n_0_657_264;
   wire n_0_842;
   wire n_0_657_265;
   wire n_0_657_266;
   wire n_0_657_267;
   wire n_0_657_268;
   wire n_0_657_269;
   wire n_0_657_270;
   wire n_0_843;
   wire n_0_657_271;
   wire n_0_657_272;
   wire n_0_657_273;
   wire n_0_657_274;
   wire n_0_657_275;
   wire n_0_657_276;
   wire n_0_657_277;
   wire n_0_844;
   wire n_0_657_278;
   wire n_0_657_279;
   wire n_0_657_280;
   wire n_0_657_281;
   wire n_0_657_282;
   wire n_0_657_283;
   wire n_0_657_284;
   wire n_0_845;
   wire n_0_657_285;
   wire n_0_657_286;
   wire n_0_657_287;
   wire n_0_657_288;
   wire n_0_657_289;
   wire n_0_657_290;
   wire n_0_657_291;
   wire n_0_657_292;
   wire n_0_846;
   wire n_0_657_293;
   wire n_0_657_294;
   wire n_0_657_295;
   wire n_0_657_296;
   wire n_0_657_297;
   wire n_0_657_298;
   wire n_0_657_299;
   wire n_0_847;
   wire n_0_657_300;
   wire n_0_657_301;
   wire n_0_657_302;
   wire n_0_657_303;
   wire n_0_657_304;
   wire n_0_657_305;
   wire n_0_657_306;
   wire n_0_657_307;
   wire n_0_849;
   wire n_0_657_308;
   wire n_0_657_309;
   wire n_0_657_310;
   wire n_0_657_311;
   wire n_0_657_312;
   wire n_0_657_313;
   wire n_0_657_314;
   wire n_0_850;
   wire n_0_657_315;
   wire n_0_657_316;
   wire n_0_657_317;
   wire n_0_657_318;
   wire n_0_657_319;
   wire n_0_657_320;
   wire n_0_657_321;
   wire n_0_851;
   wire n_0_657_322;
   wire n_0_657_323;
   wire n_0_657_324;
   wire n_0_657_325;
   wire n_0_657_326;
   wire n_0_657_327;
   wire n_0_657_328;
   wire n_0_852;
   wire n_0_657_329;
   wire n_0_657_330;
   wire n_0_657_331;
   wire n_0_657_332;
   wire n_0_657_333;
   wire n_0_657_334;
   wire n_0_657_335;
   wire n_0_853;
   wire n_0_657_336;
   wire n_0_657_337;
   wire n_0_657_338;
   wire n_0_657_339;
   wire n_0_657_340;
   wire n_0_657_341;
   wire n_0_657_342;
   wire n_0_854;
   wire n_0_657_343;
   wire n_0_657_344;
   wire n_0_657_345;
   wire n_0_657_346;
   wire n_0_657_347;
   wire n_0_657_348;
   wire n_0_657_349;
   wire n_0_657_350;
   wire n_0_657_351;
   wire n_0_855;
   wire n_0_657_352;
   wire n_0_657_353;
   wire n_0_657_354;
   wire n_0_657_355;
   wire n_0_657_356;
   wire n_0_657_357;
   wire n_0_657_358;
   wire n_0_657_359;
   wire n_0_856;
   wire n_0_657_360;
   wire n_0_657_361;
   wire n_0_657_362;
   wire n_0_657_363;
   wire n_0_657_364;
   wire n_0_657_365;
   wire n_0_657_366;
   wire n_0_657_367;
   wire n_0_657_368;
   wire n_0_857;
   wire n_0_657_369;
   wire n_0_657_370;
   wire n_0_657_371;
   wire n_0_657_372;
   wire n_0_657_373;
   wire n_0_657_374;
   wire n_0_657_375;
   wire n_0_657_376;
   wire n_0_858;
   wire n_0_657_377;
   wire n_0_657_378;
   wire n_0_657_379;
   wire n_0_657_380;
   wire n_0_657_381;
   wire n_0_657_382;
   wire n_0_657_383;
   wire n_0_859;
   wire n_0_657_384;
   wire n_0_657_385;
   wire n_0_657_386;
   wire n_0_657_387;
   wire n_0_657_388;
   wire n_0_657_389;
   wire n_0_657_390;
   wire n_0_860;
   wire n_0_657_391;
   wire n_0_657_392;
   wire n_0_657_393;
   wire n_0_657_394;
   wire n_0_657_395;
   wire n_0_657_396;
   wire n_0_657_397;
   wire n_0_861;
   wire n_0_657_398;
   wire n_0_657_399;
   wire n_0_657_400;
   wire n_0_657_401;
   wire n_0_657_402;
   wire n_0_657_403;
   wire n_0_657_404;
   wire n_0_657_405;
   wire n_0_862;
   wire n_0_657_406;
   wire n_0_657_407;
   wire n_0_657_408;
   wire n_0_657_409;
   wire n_0_657_410;
   wire n_0_657_411;
   wire n_0_657_412;
   wire n_0_863;
   wire n_0_657_413;
   wire n_0_657_414;
   wire n_0_657_415;
   wire n_0_657_416;
   wire n_0_657_417;
   wire n_0_657_418;
   wire n_0_657_419;
   wire n_0_657_420;
   wire n_0_657_421;
   wire n_0_657_422;
   wire n_0_864;
   wire n_0_657_423;
   wire n_0_657_424;
   wire n_0_657_425;
   wire n_0_657_426;
   wire n_0_657_427;
   wire n_0_657_428;
   wire n_0_657_429;
   wire n_0_865;
   wire n_0_657_430;
   wire n_0_657_431;
   wire n_0_657_432;
   wire n_0_657_433;
   wire n_0_657_434;
   wire n_0_657_435;
   wire n_0_657_436;
   wire n_0_866;
   wire n_0_657_437;
   wire n_0_657_438;
   wire n_0_657_439;
   wire n_0_657_440;
   wire n_0_657_441;
   wire n_0_657_442;
   wire n_0_867;
   wire n_0_657_443;
   wire n_0_657_444;
   wire n_0_657_445;
   wire n_0_657_446;
   wire n_0_657_447;
   wire n_0_657_448;
   wire n_0_657_449;
   wire n_0_868;
   wire n_0_657_450;
   wire n_0_657_451;
   wire n_0_657_452;
   wire n_0_657_453;
   wire n_0_657_454;
   wire n_0_657_455;
   wire n_0_657_456;
   wire n_0_657_457;
   wire n_0_869;
   wire n_0_657_458;
   wire n_0_657_459;
   wire n_0_657_460;
   wire n_0_657_461;
   wire n_0_657_462;
   wire n_0_657_463;
   wire n_0_657_464;
   wire n_0_657_465;
   wire n_0_870;
   wire n_0_657_466;
   wire n_0_657_467;
   wire n_0_657_468;
   wire n_0_657_469;
   wire n_0_657_470;
   wire n_0_657_471;
   wire n_0_657_472;
   wire n_0_657_473;
   wire n_0_871;
   wire n_0_657_474;
   wire n_0_657_475;
   wire n_0_657_476;
   wire n_0_657_477;
   wire n_0_657_478;
   wire n_0_657_479;
   wire n_0_657_480;
   wire n_0_657_481;
   wire n_0_872;
   wire n_0_657_482;
   wire n_0_657_483;
   wire n_0_657_484;
   wire n_0_657_485;
   wire n_0_657_486;
   wire n_0_657_487;
   wire n_0_873;
   wire n_0_657_488;
   wire n_0_657_489;
   wire n_0_657_490;
   wire n_0_657_491;
   wire n_0_657_492;
   wire n_0_657_493;
   wire n_0_874;
   wire n_0_657_494;
   wire n_0_657_495;
   wire n_0_657_496;
   wire n_0_657_497;
   wire n_0_657_498;
   wire n_0_657_499;
   wire n_0_875;
   wire n_0_657_500;
   wire n_0_657_501;
   wire n_0_657_502;
   wire n_0_657_503;
   wire n_0_657_504;
   wire n_0_657_505;
   wire n_0_657_506;
   wire n_0_657_507;
   wire n_0_657_508;
   wire n_0_876;
   wire n_0_657_509;
   wire n_0_657_510;
   wire n_0_657_511;
   wire n_0_657_512;
   wire n_0_657_513;
   wire n_0_657_514;
   wire n_0_877;
   wire n_0_657_515;
   wire n_0_657_516;
   wire n_0_657_517;
   wire n_0_657_518;
   wire n_0_657_519;
   wire n_0_657_520;
   wire n_0_657_521;
   wire n_0_878;
   wire n_0_657_522;
   wire n_0_657_523;
   wire n_0_657_524;
   wire n_0_657_525;
   wire n_0_657_526;
   wire n_0_657_527;
   wire n_0_880;
   wire n_0_657_528;
   wire n_0_657_529;
   wire n_0_657_530;
   wire n_0_657_531;
   wire n_0_657_532;
   wire n_0_657_533;
   wire n_0_657_534;
   wire n_0_881;
   wire n_0_657_535;
   wire n_0_657_536;
   wire n_0_657_537;
   wire n_0_657_538;
   wire n_0_657_539;
   wire n_0_657_540;
   wire n_0_657_541;
   wire n_0_882;
   wire n_0_657_542;
   wire n_0_657_543;
   wire n_0_657_544;
   wire n_0_657_545;
   wire n_0_657_546;
   wire n_0_657_547;
   wire n_0_657_548;
   wire n_0_883;
   wire n_0_657_549;
   wire n_0_657_550;
   wire n_0_657_551;
   wire n_0_657_552;
   wire n_0_657_553;
   wire n_0_657_554;
   wire n_0_657_555;
   wire n_0_657_556;
   wire n_0_657_557;
   wire n_0_657_558;
   wire n_0_657_559;
   wire n_0_884;
   wire n_0_657_560;
   wire n_0_657_561;
   wire n_0_657_562;
   wire n_0_657_563;
   wire n_0_657_564;
   wire n_0_657_565;
   wire n_0_657_566;
   wire n_0_885;
   wire n_0_657_567;
   wire n_0_657_568;
   wire n_0_657_569;
   wire n_0_657_570;
   wire n_0_657_571;
   wire n_0_657_572;
   wire n_0_657_573;
   wire n_0_657_574;
   wire n_0_886;
   wire n_0_657_575;
   wire n_0_657_576;
   wire n_0_657_577;
   wire n_0_657_578;
   wire n_0_657_579;
   wire n_0_657_580;
   wire n_0_657_581;
   wire n_0_887;
   wire n_0_657_582;
   wire n_0_657_583;
   wire n_0_657_584;
   wire n_0_657_585;
   wire n_0_657_586;
   wire n_0_657_587;
   wire n_0_657_588;
   wire n_0_657_589;
   wire n_0_888;
   wire n_0_657_590;
   wire n_0_657_591;
   wire n_0_657_592;
   wire n_0_657_593;
   wire n_0_657_594;
   wire n_0_657_595;
   wire n_0_657_596;
   wire n_0_657_597;
   wire n_0_889;
   wire n_0_657_598;
   wire n_0_657_599;
   wire n_0_657_600;
   wire n_0_657_601;
   wire n_0_657_602;
   wire n_0_657_603;
   wire n_0_657_604;
   wire n_0_890;
   wire n_0_657_605;
   wire n_0_657_606;
   wire n_0_657_607;
   wire n_0_657_608;
   wire n_0_657_609;
   wire n_0_657_610;
   wire n_0_657_611;
   wire n_0_657_612;
   wire n_0_891;
   wire n_0_657_613;
   wire n_0_657_614;
   wire n_0_657_615;
   wire n_0_657_616;
   wire n_0_657_617;
   wire n_0_657_618;
   wire n_0_657_619;
   wire n_0_657_620;
   wire n_0_892;
   wire n_0_657_621;
   wire n_0_657_622;
   wire n_0_657_623;
   wire n_0_657_624;
   wire n_0_657_625;
   wire n_0_657_626;
   wire n_0_657_627;
   wire n_0_893;
   wire n_0_657_628;
   wire n_0_657_629;
   wire n_0_657_630;
   wire n_0_657_631;
   wire n_0_657_632;
   wire n_0_657_633;
   wire n_0_657_634;
   wire n_0_894;
   wire n_0_657_635;
   wire n_0_657_636;
   wire n_0_657_637;
   wire n_0_657_638;
   wire n_0_657_639;
   wire n_0_657_640;
   wire n_0_657_641;
   wire n_0_902;
   wire n_0_657_642;
   wire n_0_657_643;
   wire n_0_657_644;
   wire n_0_657_645;
   wire n_0_657_646;
   wire n_0_657_647;
   wire n_0_657_648;
   wire n_0_657_649;
   wire n_0_657_650;
   wire n_0_657_651;
   wire n_0_657_652;
   wire n_0_903;
   wire n_0_657_653;
   wire n_0_657_654;
   wire n_0_657_655;
   wire n_0_657_656;
   wire n_0_657_657;
   wire n_0_657_658;
   wire n_0_657_659;
   wire n_0_657_660;
   wire n_0_904;
   wire n_0_657_661;
   wire n_0_657_662;
   wire n_0_657_663;
   wire n_0_657_664;
   wire n_0_657_665;
   wire n_0_657_666;
   wire n_0_657_667;
   wire n_0_657_668;
   wire n_0_905;
   wire n_0_657_669;
   wire n_0_657_670;
   wire n_0_657_671;
   wire n_0_657_672;
   wire n_0_657_673;
   wire n_0_657_674;
   wire n_0_657_675;
   wire n_0_657_676;
   wire n_0_906;
   wire n_0_657_677;
   wire n_0_657_678;
   wire n_0_657_679;
   wire n_0_657_680;
   wire n_0_657_681;
   wire n_0_657_682;
   wire n_0_657_683;
   wire n_0_907;
   wire n_0_657_684;
   wire n_0_657_685;
   wire n_0_657_686;
   wire n_0_657_687;
   wire n_0_657_688;
   wire n_0_657_689;
   wire n_0_657_690;
   wire n_0_657_691;
   wire n_0_908;
   wire n_0_657_692;
   wire n_0_657_693;
   wire n_0_657_694;
   wire n_0_657_695;
   wire n_0_657_696;
   wire n_0_657_697;
   wire n_0_657_698;
   wire n_0_657_699;
   wire n_0_909;
   wire n_0_657_700;
   wire n_0_657_701;
   wire n_0_657_702;
   wire n_0_657_703;
   wire n_0_657_704;
   wire n_0_657_705;
   wire n_0_657_706;
   wire n_0_657_707;
   wire n_0_910;
   wire n_0_657_708;
   wire n_0_657_709;
   wire n_0_657_710;
   wire n_0_657_711;
   wire n_0_657_712;
   wire n_0_657_713;
   wire n_0_657_714;
   wire n_0_657_715;
   wire n_0_912;
   wire n_0_657_716;
   wire n_0_657_717;
   wire n_0_657_718;
   wire n_0_657_719;
   wire n_0_657_720;
   wire n_0_657_721;
   wire n_0_657_722;
   wire n_0_913;
   wire n_0_657_723;
   wire n_0_657_724;
   wire n_0_657_725;
   wire n_0_657_726;
   wire n_0_657_727;
   wire n_0_657_728;
   wire n_0_657_729;
   wire n_0_914;
   wire n_0_657_730;
   wire n_0_657_731;
   wire n_0_657_732;
   wire n_0_657_733;
   wire n_0_657_734;
   wire n_0_657_735;
   wire n_0_657_736;
   wire n_0_657_737;
   wire n_0_657_738;
   wire n_0_657_739;
   wire n_0_657_740;
   wire n_0_915;
   wire n_0_657_741;
   wire n_0_657_742;
   wire n_0_657_743;
   wire n_0_657_744;
   wire n_0_657_745;
   wire n_0_657_746;
   wire n_0_657_747;
   wire n_0_657_748;
   wire n_0_657_749;
   wire n_0_657_750;
   wire n_0_657_751;
   wire n_0_916;
   wire n_0_657_752;
   wire n_0_657_753;
   wire n_0_657_754;
   wire n_0_657_755;
   wire n_0_657_756;
   wire n_0_657_757;
   wire n_0_657_758;
   wire n_0_657_759;
   wire n_0_657_760;
   wire n_0_657_761;
   wire n_0_657_762;
   wire n_0_917;
   wire n_0_657_763;
   wire n_0_657_764;
   wire n_0_657_765;
   wire n_0_657_766;
   wire n_0_657_767;
   wire n_0_657_768;
   wire n_0_657_769;
   wire n_0_657_770;
   wire n_0_657_771;
   wire n_0_657_772;
   wire n_0_657_773;
   wire n_0_918;
   wire n_0_657_774;
   wire n_0_657_775;
   wire n_0_657_776;
   wire n_0_657_777;
   wire n_0_657_778;
   wire n_0_657_779;
   wire n_0_657_780;
   wire n_0_919;
   wire n_0_657_781;
   wire n_0_657_782;
   wire n_0_657_783;
   wire n_0_657_784;
   wire n_0_657_785;
   wire n_0_657_786;
   wire n_0_657_787;
   wire n_0_921;
   wire n_0_657_788;
   wire n_0_657_789;
   wire n_0_657_790;
   wire n_0_657_791;
   wire n_0_657_792;
   wire n_0_657_793;
   wire n_0_657_794;
   wire n_0_923;
   wire n_0_657_795;
   wire n_0_657_796;
   wire n_0_657_797;
   wire n_0_657_798;
   wire n_0_657_799;
   wire n_0_657_800;
   wire n_0_657_801;
   wire n_0_924;
   wire n_0_657_802;
   wire n_0_657_803;
   wire n_0_657_804;
   wire n_0_657_805;
   wire n_0_657_806;
   wire n_0_657_807;
   wire n_0_657_808;
   wire n_0_657_809;
   wire n_0_657_810;
   wire n_0_925;
   wire n_0_657_811;
   wire n_0_657_812;
   wire n_0_657_813;
   wire n_0_657_814;
   wire n_0_657_815;
   wire n_0_657_816;
   wire n_0_657_817;
   wire n_0_657_818;
   wire n_0_657_819;
   wire n_0_657_820;
   wire n_0_926;
   wire n_0_657_821;
   wire n_0_657_822;
   wire n_0_657_823;
   wire n_0_657_824;
   wire n_0_657_825;
   wire n_0_657_826;
   wire n_0_657_827;
   wire n_0_927;
   wire n_0_657_828;
   wire n_0_657_829;
   wire n_0_657_830;
   wire n_0_657_831;
   wire n_0_657_832;
   wire n_0_657_833;
   wire n_0_657_834;
   wire n_0_928;
   wire n_0_657_835;
   wire n_0_657_836;
   wire n_0_657_837;
   wire n_0_657_838;
   wire n_0_657_839;
   wire n_0_657_840;
   wire n_0_657_841;
   wire n_0_929;
   wire n_0_657_842;
   wire n_0_657_843;
   wire n_0_657_844;
   wire n_0_657_845;
   wire n_0_657_846;
   wire n_0_657_847;
   wire n_0_657_848;
   wire n_0_930;
   wire n_0_657_849;
   wire n_0_657_850;
   wire n_0_657_851;
   wire n_0_657_852;
   wire n_0_657_853;
   wire n_0_657_854;
   wire n_0_657_855;
   wire n_0_931;
   wire n_0_657_856;
   wire n_0_657_857;
   wire n_0_657_858;
   wire n_0_657_859;
   wire n_0_657_860;
   wire n_0_657_861;
   wire n_0_657_862;
   wire n_0_932;
   wire n_0_657_863;
   wire n_0_657_864;
   wire n_0_657_865;
   wire n_0_657_866;
   wire n_0_657_867;
   wire n_0_657_868;
   wire n_0_657_869;
   wire n_0_933;
   wire n_0_657_870;
   wire n_0_657_871;
   wire n_0_657_872;
   wire n_0_657_873;
   wire n_0_657_874;
   wire n_0_657_875;
   wire n_0_657_876;
   wire n_0_935;
   wire n_0_657_877;
   wire n_0_657_878;
   wire n_0_657_879;
   wire n_0_657_880;
   wire n_0_657_881;
   wire n_0_936;
   wire n_0_657_882;
   wire n_0_657_883;
   wire n_0_657_884;
   wire n_0_657_885;
   wire n_0_657_886;
   wire n_0_657_887;
   wire n_0_657_888;
   wire n_0_937;
   wire n_0_657_889;
   wire n_0_657_890;
   wire n_0_657_891;
   wire n_0_657_892;
   wire n_0_657_893;
   wire n_0_657_894;
   wire n_0_657_895;
   wire n_0_657_896;
   wire n_0_657_897;
   wire n_0_657_898;
   wire n_0_938;
   wire n_0_657_899;
   wire n_0_657_900;
   wire n_0_657_901;
   wire n_0_657_902;
   wire n_0_657_903;
   wire n_0_940;
   wire n_0_657_904;
   wire n_0_657_905;
   wire n_0_657_906;
   wire n_0_657_907;
   wire n_0_657_908;
   wire n_0_657_909;
   wire n_0_657_910;
   wire n_0_657_911;
   wire n_0_657_912;
   wire n_0_657_913;
   wire n_0_942;
   wire n_0_657_914;
   wire n_0_657_915;
   wire n_0_657_916;
   wire n_0_657_917;
   wire n_0_657_918;
   wire n_0_657_919;
   wire n_0_657_920;
   wire n_0_943;
   wire n_0_657_921;
   wire n_0_657_922;
   wire n_0_657_923;
   wire n_0_657_924;
   wire n_0_657_925;
   wire n_0_657_926;
   wire n_0_657_927;
   wire n_0_944;
   wire n_0_657_928;
   wire n_0_657_929;
   wire n_0_657_930;
   wire n_0_657_931;
   wire n_0_657_932;
   wire n_0_657_933;
   wire n_0_657_934;
   wire n_0_946;
   wire n_0_657_935;
   wire n_0_657_936;
   wire n_0_657_937;
   wire n_0_657_938;
   wire n_0_657_939;
   wire n_0_657_940;
   wire n_0_657_941;
   wire n_0_947;
   wire n_0_657_942;
   wire n_0_657_943;
   wire n_0_657_944;
   wire n_0_657_945;
   wire n_0_657_946;
   wire n_0_948;
   wire n_0_657_947;
   wire n_0_657_948;
   wire n_0_657_949;
   wire n_0_657_950;
   wire n_0_657_951;
   wire n_0_657_952;
   wire n_0_657_953;
   wire n_0_657_954;
   wire n_0_657_955;
   wire n_0_949;
   wire n_0_657_956;
   wire n_0_657_957;
   wire n_0_657_958;
   wire n_0_657_959;
   wire n_0_657_960;
   wire n_0_657_961;
   wire n_0_657_962;
   wire n_0_657_963;
   wire n_0_657_964;
   wire n_2_0_0;
   wire n_2_0_1;
   wire n_2_1_0;
   wire n_2_1_1;
   wire n_2_2_0;
   wire n_2_2_1;
   wire n_2_3_0;
   wire n_2_3_1;
   wire n_2_4_0;
   wire n_2_4_1;
   wire n_2_5_0;
   wire n_2_5_1;
   wire n_2_6_0;
   wire n_2_6_1;
   wire n_2_7_0;
   wire n_2_7_1;
   wire n_2_8_0;
   wire n_2_8_1;
   wire n_2_9_0;
   wire n_2_9_1;
   wire n_2_10_0;
   wire n_2_10_1;
   wire n_2_11_0;
   wire n_2_11_1;
   wire n_2_12_0;
   wire n_2_12_1;
   wire n_2_13_0;
   wire n_2_13_1;
   wire n_2_14_0;
   wire n_2_14_1;
   wire n_2_15_0;
   wire n_2_15_1;
   wire n_2_16_0;
   wire n_2_16_1;
   wire n_2_17_0;
   wire n_2_17_1;
   wire n_2_18_0;
   wire n_2_18_1;
   wire n_2_19_0;
   wire n_2_19_1;
   wire n_2_20_0;
   wire n_2_20_1;
   wire n_2_21_0;
   wire n_2_21_1;
   wire n_2_22_0;
   wire n_2_22_1;
   wire n_2_23_0;
   wire n_2_23_1;
   wire n_2_24_0;
   wire n_2_24_1;
   wire n_2_25_0;
   wire n_2_25_1;
   wire n_2_26_0;
   wire n_2_26_1;
   wire n_2_27_0;
   wire n_2_27_1;
   wire n_2_28_0;
   wire n_2_28_1;
   wire n_2_29_0;
   wire n_2_29_1;
   wire n_2_30_0;
   wire n_2_30_1;
   wire n_2_31_0;
   wire n_2_31_1;
   wire n_2_32_0;
   wire n_2_32_1;
   wire n_2_33_0;
   wire n_2_33_1;
   wire n_2_34_0;
   wire n_2_34_1;
   wire n_2_35_0;
   wire n_2_35_1;
   wire n_2_36_0;
   wire n_2_36_1;
   wire n_2_37_0;
   wire n_2_37_1;
   wire n_2_38_0;
   wire n_2_38_1;
   wire n_2_39_0;
   wire n_2_39_1;
   wire n_2_40_0;
   wire n_2_40_1;
   wire n_2_41_0;
   wire n_2_41_1;
   wire n_2_42_0;
   wire n_2_42_1;
   wire n_2_43_0;
   wire n_2_43_1;
   wire n_2_44_0;
   wire n_2_44_1;
   wire n_2_45_0;
   wire n_2_45_1;
   wire n_2_46_0;
   wire n_2_46_1;
   wire n_2_47_0;
   wire n_2_47_1;
   wire n_2_48_0;
   wire n_2_48_1;
   wire n_2_49_0;
   wire n_2_49_1;
   wire n_2_50_0;
   wire n_2_50_1;
   wire n_2_51_0;
   wire n_2_51_1;
   wire n_2_52_0;
   wire n_2_52_1;
   wire n_2_53_0;
   wire n_2_53_1;
   wire n_2_54_0;
   wire n_2_54_1;
   wire n_2_55_0;
   wire n_2_55_1;
   wire n_2_56_0;
   wire n_2_56_1;
   wire n_2_57_0;
   wire n_2_57_1;
   wire n_2_58_0;
   wire n_2_58_1;
   wire n_2_59_0;
   wire n_2_59_1;
   wire n_2_60_0;
   wire n_2_60_1;
   wire n_2_61_0;
   wire n_2_61_1;
   wire n_2_62_0;
   wire n_2_62_1;
   wire n_2_63_0;
   wire n_2_63_1;
   wire n_2_64_0;
   wire n_2_64_1;
   wire n_2_65_0;
   wire n_2_65_1;
   wire n_2_66_0;
   wire n_2_66_1;
   wire n_2_67_0;
   wire n_2_67_1;
   wire n_2_68_0;
   wire n_2_68_1;
   wire n_2_69_0;
   wire n_2_69_1;
   wire n_2_70_0;
   wire n_2_70_1;
   wire n_2_71_0;
   wire n_2_71_1;
   wire n_2_72_0;
   wire n_2_72_1;
   wire n_2_72_2;
   wire n_2_72_3;
   wire n_2_73_0;
   wire n_2_73_1;
   wire n_2_73_2;
   wire n_2_73_3;
   wire n_2_74_0;
   wire n_2_74_1;
   wire n_2_74_2;
   wire n_2_74_3;
   wire n_2_75_0;
   wire n_2_75_1;
   wire n_2_75_2;
   wire n_2_75_3;
   wire n_2_1;
   wire n_2_76_0;
   wire n_2_76_1;
   wire n_2_4;
   wire n_2_77_0;
   wire n_2_77_1;
   wire n_2_5;
   wire n_2_78_0;
   wire n_2_78_1;
   wire n_2_17;
   wire n_2_79_0;
   wire n_2_79_1;
   wire n_2_21;
   wire n_2_81_0;
   wire n_2_81_1;
   wire n_2_22;
   wire n_2_82_0;
   wire n_2_82_1;
   wire n_2_28;
   wire n_2_83_0;
   wire n_2_83_1;
   wire n_2_38;
   wire n_2_84_0;
   wire n_2_84_1;
   wire n_2_50;
   wire n_2_85_0;
   wire n_2_85_1;
   wire n_2_53;
   wire n_2_86_0;
   wire n_2_86_1;
   wire n_2_56;
   wire n_2_87_0;
   wire n_2_87_1;
   wire n_2_60;
   wire n_2_88_0;
   wire n_2_88_1;
   wire n_2_67;
   wire n_2_89_0;
   wire n_2_89_1;
   wire n_2_68;
   wire n_2_90_0;
   wire n_2_90_1;
   wire n_2_69;
   wire n_2_91_0;
   wire n_2_91_1;
   wire n_2_70;
   wire n_2_92_0;
   wire n_2_92_1;
   wire n_2_71;
   wire n_2_93_0;
   wire n_2_93_1;
   wire n_2_75;
   wire n_2_94_0;
   wire n_2_94_1;
   wire n_2_76;
   wire n_2_95_0;
   wire n_2_95_1;
   wire n_2_77;
   wire n_2_96_0;
   wire n_2_96_1;
   wire n_2_78;
   wire n_2_97_0;
   wire n_2_97_1;
   wire n_2_80;
   wire n_2_98_0;
   wire n_2_98_1;
   wire n_2_83;
   wire n_2_99_0;
   wire n_2_99_1;
   wire n_2_86;
   wire n_2_100_0;
   wire n_2_100_1;
   wire n_2_89;
   wire n_2_101_0;
   wire n_2_101_1;
   wire n_2_90;
   wire n_2_102_0;
   wire n_2_102_1;
   wire n_2_91;
   wire n_2_103_0;
   wire n_2_103_1;
   wire n_2_93;
   wire n_2_104_0;
   wire n_2_104_1;
   wire n_2_94;
   wire n_2_105_0;
   wire n_2_105_1;
   wire n_2_97;
   wire n_2_106_0;
   wire n_2_106_1;
   wire n_2_100;
   wire n_2_107_0;
   wire n_2_107_1;
   wire n_2_102;
   wire n_2_108_0;
   wire n_2_108_1;
   wire n_2_104;
   wire n_2_109_0;
   wire n_2_109_1;
   wire n_2_112;
   wire n_2_110_0;
   wire n_2_110_1;
   wire n_2_113;
   wire n_2_111_0;
   wire n_2_111_1;
   wire n_2_116;
   wire n_2_112_0;
   wire n_2_112_1;
   wire n_2_119;
   wire n_2_113_0;
   wire n_2_113_1;
   wire n_2_120;
   wire n_2_114_0;
   wire n_2_114_1;
   wire n_2_121;
   wire n_2_115_0;
   wire n_2_115_1;
   wire n_2_122;
   wire n_2_116_0;
   wire n_2_116_1;
   wire n_2_123;
   wire n_2_117_0;
   wire n_2_117_1;
   wire n_2_126;
   wire n_2_118_0;
   wire n_2_118_1;
   wire n_2_127;
   wire n_2_119_0;
   wire n_2_119_1;
   wire n_2_128;
   wire n_2_120_0;
   wire n_2_120_1;
   wire n_2_129;
   wire n_2_121_0;
   wire n_2_121_1;
   wire n_2_138;
   wire n_2_122_0;
   wire n_2_122_1;
   wire n_2_142;
   wire n_2_123_0;
   wire n_2_123_1;
   wire n_2_150;
   wire n_2_124_0;
   wire n_2_124_1;
   wire n_2_153;
   wire n_2_125_0;
   wire n_2_125_1;
   wire n_2_156;
   wire n_2_126_0;
   wire n_2_126_1;
   wire n_2_157;
   wire n_2_127_0;
   wire n_2_127_1;
   wire n_2_160;
   wire n_2_128_0;
   wire n_2_128_1;
   wire n_2_161;
   wire n_2_129_0;
   wire n_2_129_1;
   wire n_2_162;
   wire n_2_130_0;
   wire n_2_130_1;
   wire n_2_163;
   wire n_2_131_0;
   wire n_2_131_1;
   wire n_2_167;
   wire n_2_132_0;
   wire n_2_132_1;
   wire n_2_168;
   wire n_2_133_0;
   wire n_2_133_1;
   wire n_2_172;
   wire n_2_134_0;
   wire n_2_134_1;
   wire n_2_173;
   wire n_2_135_0;
   wire n_2_135_1;
   wire n_2_174;
   wire n_2_136_0;
   wire n_2_136_1;
   wire n_2_180;
   wire n_2_137_0;
   wire n_2_137_1;
   wire n_2_184;
   wire n_2_138_0;
   wire n_2_138_1;
   wire n_2_185;
   wire n_2_139_0;
   wire n_2_139_1;
   wire n_2_188;
   wire n_2_140_0;
   wire n_2_140_1;
   wire n_2_194;
   wire n_2_141_0;
   wire n_2_141_1;
   wire n_2_196;
   wire n_2_142_0;
   wire n_2_142_1;
   wire n_2_197;
   wire n_2_143_0;
   wire n_2_143_1;
   wire n_2_198;
   wire n_2_144_0;
   wire n_2_144_1;
   wire n_2_201;
   wire n_2_145_0;
   wire n_2_145_1;
   wire n_2_202;
   wire n_2_146_0;
   wire n_2_146_1;
   wire n_2_203;
   wire n_2_147_0;
   wire n_2_147_1;
   wire n_2_205;
   wire n_2_148_0;
   wire n_2_148_1;
   wire n_2_225;
   wire n_2_149_0;
   wire n_2_149_1;
   wire n_2_149_2;
   wire n_2_149_3;
   wire n_2_226;
   wire n_2_150_0;
   wire n_2_150_1;
   wire n_2_150_2;
   wire n_2_150_3;
   wire n_2_227;
   wire n_2_151_0;
   wire n_2_151_1;
   wire n_2_151_2;
   wire n_2_151_3;
   wire n_2_228;
   wire n_2_152_0;
   wire n_2_152_1;
   wire n_2_152_2;
   wire n_2_152_3;
   wire n_2_154_0;
   wire n_2_154_1;
   wire n_2_154_2;
   wire n_2_154_3;
   wire n_2_241;
   wire n_2_339;
   wire n_2_156_0;
   wire n_2_156_1;
   wire n_2_156_2;
   wire n_2_156_3;
   wire n_2_157_0;
   wire n_2_157_1;
   wire n_2_157_2;
   wire n_2_157_3;
   wire n_2_158_0;
   wire n_2_158_1;
   wire n_2_158_2;
   wire n_2_158_3;
   wire n_2_159_0;
   wire n_2_159_1;
   wire n_2_159_2;
   wire n_2_159_3;
   wire n_2_160_0;
   wire n_2_160_1;
   wire n_2_160_2;
   wire n_2_160_3;
   wire n_2_161_0;
   wire n_2_161_1;
   wire n_2_161_2;
   wire n_2_161_3;
   wire n_2_162_0;
   wire n_2_162_1;
   wire n_2_162_2;
   wire n_2_162_3;
   wire n_2_163_0;
   wire n_2_163_1;
   wire n_2_163_2;
   wire n_2_163_3;
   wire n_2_164_0;
   wire n_2_164_1;
   wire n_2_164_2;
   wire n_2_164_3;
   wire n_2_165_0;
   wire n_2_165_1;
   wire n_2_165_2;
   wire n_2_165_3;
   wire n_2_166_0;
   wire n_2_166_1;
   wire n_2_166_2;
   wire n_2_166_3;
   wire n_2_167_0;
   wire n_2_167_1;
   wire n_2_167_2;
   wire n_2_167_3;
   wire n_2_168_0;
   wire n_2_168_1;
   wire n_2_168_2;
   wire n_2_168_3;
   wire n_2_169_0;
   wire n_2_169_1;
   wire n_2_169_2;
   wire n_2_169_3;
   wire n_2_170_0;
   wire n_2_170_1;
   wire n_2_170_2;
   wire n_2_170_3;
   wire n_2_171_0;
   wire n_2_171_1;
   wire n_2_171_2;
   wire n_2_171_3;
   wire n_2_172_0;
   wire n_2_172_1;
   wire n_2_172_2;
   wire n_2_172_3;
   wire n_2_173_0;
   wire n_2_173_1;
   wire n_2_173_2;
   wire n_2_173_3;
   wire n_2_174_0;
   wire n_2_174_1;
   wire n_2_174_2;
   wire n_2_174_3;
   wire n_2_175_0;
   wire n_2_175_1;
   wire n_2_175_2;
   wire n_2_175_3;
   wire n_2_176_0;
   wire n_2_176_1;
   wire n_2_176_2;
   wire n_2_176_3;
   wire n_2_177_0;
   wire n_2_177_1;
   wire n_2_177_2;
   wire n_2_177_3;
   wire n_2_178_0;
   wire n_2_178_1;
   wire n_2_178_2;
   wire n_2_178_3;
   wire n_2_179_0;
   wire n_2_179_1;
   wire n_2_179_2;
   wire n_2_179_3;
   wire n_2_180_0;
   wire n_2_180_1;
   wire n_2_180_2;
   wire n_2_180_3;
   wire n_2_181_0;
   wire n_2_181_1;
   wire n_2_181_2;
   wire n_2_181_3;
   wire n_2_182_0;
   wire n_2_182_1;
   wire n_2_182_2;
   wire n_2_182_3;
   wire n_2_183_0;
   wire n_2_183_1;
   wire n_2_183_2;
   wire n_2_183_3;
   wire n_2_184_0;
   wire n_2_184_1;
   wire n_2_184_2;
   wire n_2_184_3;
   wire n_2_185_0;
   wire n_2_185_1;
   wire n_2_185_2;
   wire n_2_185_3;
   wire n_2_186_0;
   wire n_2_186_1;
   wire n_2_186_2;
   wire n_2_186_3;
   wire n_2_187_0;
   wire n_2_187_1;
   wire n_2_187_2;
   wire n_2_187_3;
   wire n_2_188_0;
   wire n_2_188_1;
   wire n_2_188_2;
   wire n_2_188_3;
   wire n_2_189_0;
   wire n_2_189_1;
   wire n_2_189_2;
   wire n_2_189_3;
   wire n_2_190_0;
   wire n_2_190_1;
   wire n_2_190_2;
   wire n_2_190_3;
   wire n_2_191_0;
   wire n_2_191_1;
   wire n_2_191_2;
   wire n_2_191_3;
   wire n_2_192_0;
   wire n_2_192_1;
   wire n_2_192_2;
   wire n_2_192_3;
   wire n_2_193_0;
   wire n_2_193_1;
   wire n_2_193_2;
   wire n_2_193_3;
   wire n_2_194_0;
   wire n_2_194_1;
   wire n_2_194_2;
   wire n_2_194_3;
   wire n_2_195_0;
   wire n_2_195_1;
   wire n_2_195_2;
   wire n_2_195_3;
   wire n_2_196_0;
   wire n_2_196_1;
   wire n_2_196_2;
   wire n_2_196_3;
   wire n_2_197_0;
   wire n_2_197_1;
   wire n_2_197_2;
   wire n_2_197_3;
   wire n_2_198_0;
   wire n_2_198_1;
   wire n_2_198_2;
   wire n_2_198_3;
   wire n_2_199_0;
   wire n_2_199_1;
   wire n_2_199_2;
   wire n_2_199_3;
   wire n_2_200_0;
   wire n_2_200_1;
   wire n_2_200_2;
   wire n_2_200_3;
   wire n_2_201_0;
   wire n_2_201_1;
   wire n_2_201_2;
   wire n_2_201_3;
   wire n_2_202_0;
   wire n_2_202_1;
   wire n_2_202_2;
   wire n_2_202_3;
   wire n_2_203_0;
   wire n_2_203_1;
   wire n_2_203_2;
   wire n_2_203_3;
   wire n_2_204_0;
   wire n_2_204_1;
   wire n_2_204_2;
   wire n_2_204_3;
   wire n_2_205_0;
   wire n_2_205_1;
   wire n_2_205_2;
   wire n_2_205_3;
   wire n_2_206_0;
   wire n_2_206_1;
   wire n_2_206_2;
   wire n_2_206_3;
   wire n_2_207_0;
   wire n_2_207_1;
   wire n_2_207_2;
   wire n_2_207_3;
   wire n_2_208_0;
   wire n_2_208_1;
   wire n_2_208_2;
   wire n_2_208_3;
   wire n_2_209_0;
   wire n_2_209_1;
   wire n_2_209_2;
   wire n_2_209_3;
   wire n_2_210_0;
   wire n_2_210_1;
   wire n_2_210_2;
   wire n_2_210_3;
   wire n_2_211_0;
   wire n_2_211_1;
   wire n_2_211_2;
   wire n_2_211_3;
   wire n_2_212_0;
   wire n_2_212_1;
   wire n_2_212_2;
   wire n_2_212_3;
   wire n_2_213_0;
   wire n_2_213_1;
   wire n_2_213_2;
   wire n_2_213_3;
   wire n_2_214_0;
   wire n_2_214_1;
   wire n_2_214_2;
   wire n_2_214_3;
   wire n_2_215_0;
   wire n_2_215_1;
   wire n_2_215_2;
   wire n_2_215_3;
   wire n_2_216_0;
   wire n_2_216_1;
   wire n_2_216_2;
   wire n_2_216_3;
   wire n_2_217_0;
   wire n_2_217_1;
   wire n_2_217_2;
   wire n_2_217_3;
   wire n_2_218_0;
   wire n_2_218_1;
   wire n_2_218_2;
   wire n_2_218_3;
   wire n_2_219_0;
   wire n_2_219_1;
   wire n_2_219_2;
   wire n_2_219_3;
   wire n_2_220_0;
   wire n_2_220_1;
   wire n_2_220_2;
   wire n_2_220_3;
   wire n_2_221_0;
   wire n_2_221_1;
   wire n_2_221_2;
   wire n_2_221_3;
   wire n_2_222_0;
   wire n_2_222_1;
   wire n_2_222_2;
   wire n_2_222_3;
   wire n_2_223_0;
   wire n_2_223_1;
   wire n_2_223_2;
   wire n_2_223_3;
   wire n_2_224_0;
   wire n_2_224_1;
   wire n_2_224_2;
   wire n_2_224_3;
   wire n_2_225_0;
   wire n_2_225_1;
   wire n_2_225_2;
   wire n_2_225_3;
   wire n_2_226_0;
   wire n_2_226_1;
   wire n_2_226_2;
   wire n_2_226_3;
   wire n_2_227_0;
   wire n_2_227_1;
   wire n_2_227_2;
   wire n_2_227_3;
   wire n_2_228_0;
   wire n_2_228_1;
   wire n_2_228_2;
   wire n_2_228_3;
   wire n_2_229_0;
   wire n_2_229_1;
   wire n_2_229_2;
   wire n_2_229_3;
   wire n_2_230_0;
   wire n_2_230_1;
   wire n_2_230_2;
   wire n_2_230_3;
   wire n_2_231_0;
   wire n_2_231_1;
   wire n_2_231_2;
   wire n_2_231_3;
   wire n_2_232_0;
   wire n_2_232_1;
   wire n_2_232_2;
   wire n_2_232_3;
   wire n_2_233_0;
   wire n_2_233_1;
   wire n_2_233_2;
   wire n_2_233_3;
   wire n_2_234_0;
   wire n_2_234_1;
   wire n_2_234_2;
   wire n_2_234_3;
   wire n_2_235_0;
   wire n_2_235_1;
   wire n_2_235_2;
   wire n_2_235_3;
   wire n_2_0;
   wire n_2_236_0;
   wire n_2_236_1;
   wire n_2_236_2;
   wire n_2_236_3;
   wire n_2_237_0;
   wire n_2_237_1;
   wire n_2_237_2;
   wire n_2_237_3;
   wire n_2_238_0;
   wire n_2_238_1;
   wire n_2_238_2;
   wire n_2_238_3;
   wire n_2_239_0;
   wire n_2_239_1;
   wire n_2_239_2;
   wire n_2_239_3;
   wire n_2_240_0;
   wire n_2_240_1;
   wire n_2_240_2;
   wire n_2_240_3;
   wire n_2_241_0;
   wire n_2_241_1;
   wire n_2_241_2;
   wire n_2_241_3;
   wire n_2_242_0;
   wire n_2_242_1;
   wire n_2_242_2;
   wire n_2_242_3;
   wire n_2_243_0;
   wire n_2_243_1;
   wire n_2_243_2;
   wire n_2_243_3;
   wire n_2_244_0;
   wire n_2_244_1;
   wire n_2_244_2;
   wire n_2_244_3;
   wire n_2_245_0;
   wire n_2_245_1;
   wire n_2_245_2;
   wire n_2_245_3;
   wire n_2_246_0;
   wire n_2_246_1;
   wire n_2_246_2;
   wire n_2_246_3;
   wire n_2_247_0;
   wire n_2_247_1;
   wire n_2_247_2;
   wire n_2_247_3;
   wire n_2_248_0;
   wire n_2_248_1;
   wire n_2_248_2;
   wire n_2_248_3;
   wire n_2_249_0;
   wire n_2_249_1;
   wire n_2_249_2;
   wire n_2_249_3;
   wire n_2_250_0;
   wire n_2_250_1;
   wire n_2_250_2;
   wire n_2_250_3;
   wire n_2_251_0;
   wire n_2_251_1;
   wire n_2_251_2;
   wire n_2_251_3;
   wire n_2_252_0;
   wire n_2_252_1;
   wire n_2_252_2;
   wire n_2_252_3;
   wire n_2_253_0;
   wire n_2_253_1;
   wire n_2_253_2;
   wire n_2_253_3;
   wire n_2_254_0;
   wire n_2_254_1;
   wire n_2_254_2;
   wire n_2_254_3;
   wire n_2_255_0;
   wire n_2_255_1;
   wire n_2_255_2;
   wire n_2_255_3;
   wire n_2_256_0;
   wire n_2_256_1;
   wire n_2_256_2;
   wire n_2_256_3;
   wire n_2_257_0;
   wire n_2_257_1;
   wire n_2_257_2;
   wire n_2_257_3;
   wire n_2_208;
   wire n_2_258_0;
   wire n_2_258_1;
   wire n_2_258_2;
   wire n_2_258_3;
   wire n_2_209;
   wire n_2_259_0;
   wire n_2_259_1;
   wire n_2_259_2;
   wire n_2_259_3;
   wire n_2_210;
   wire n_2_260_0;
   wire n_2_260_1;
   wire n_2_260_2;
   wire n_2_260_3;
   wire n_2_261_0;
   wire n_2_261_1;
   wire n_2_261_2;
   wire n_2_261_3;
   wire n_2_211;
   wire n_2_262_0;
   wire n_2_262_1;
   wire n_2_262_2;
   wire n_2_262_3;
   wire n_2_212;
   wire n_2_263_0;
   wire n_2_263_1;
   wire n_2_263_2;
   wire n_2_263_3;
   wire n_2_213;
   wire n_2_264_0;
   wire n_2_264_1;
   wire n_2_264_2;
   wire n_2_264_3;
   wire n_2_214;
   wire n_2_265_0;
   wire n_2_265_1;
   wire n_2_265_2;
   wire n_2_265_3;
   wire n_2_215;
   wire n_2_266_0;
   wire n_2_266_1;
   wire n_2_266_2;
   wire n_2_266_3;
   wire n_2_216;
   wire n_2_267_0;
   wire n_2_267_1;
   wire n_2_267_2;
   wire n_2_267_3;
   wire n_2_217;
   wire n_2_268_0;
   wire n_2_268_1;
   wire n_2_268_2;
   wire n_2_268_3;
   wire n_2_269_0;
   wire n_2_269_1;
   wire n_2_269_2;
   wire n_2_269_3;
   wire n_2_218;
   wire n_2_270_0;
   wire n_2_270_1;
   wire n_2_270_2;
   wire n_2_270_3;
   wire n_2_271_0;
   wire n_2_271_1;
   wire n_2_271_2;
   wire n_2_271_3;
   wire n_2_219;
   wire n_2_272_0;
   wire n_2_272_1;
   wire n_2_272_2;
   wire n_2_272_3;
   wire n_2_220;
   wire n_2_273_0;
   wire n_2_273_1;
   wire n_2_273_2;
   wire n_2_273_3;
   wire n_2_221;
   wire n_2_274_0;
   wire n_2_274_1;
   wire n_2_274_2;
   wire n_2_274_3;
   wire n_2_275_0;
   wire n_2_275_1;
   wire n_2_275_2;
   wire n_2_275_3;
   wire n_2_222;
   wire n_2_276_0;
   wire n_2_276_1;
   wire n_2_276_2;
   wire n_2_276_3;
   wire n_2_277_0;
   wire n_2_277_1;
   wire n_2_277_2;
   wire n_2_277_3;
   wire n_2_223;
   wire n_2_278_0;
   wire n_2_278_1;
   wire n_2_278_2;
   wire n_2_278_3;
   wire n_2_224;
   wire n_2_279_0;
   wire n_2_279_1;
   wire n_2_279_2;
   wire n_2_279_3;
   wire n_2_280_0;
   wire n_2_280_1;
   wire n_2_280_2;
   wire n_2_280_3;
   wire n_2_281_0;
   wire n_2_281_1;
   wire n_2_281_2;
   wire n_2_281_3;
   wire n_2_2;
   wire n_2_3;
   wire n_2_6;
   wire n_2_7;
   wire n_2_18;
   wire n_2_19;
   wire n_2_23;
   wire n_2_24;
   wire n_2_29;
   wire n_2_30;
   wire n_2_39;
   wire n_2_40;
   wire n_2_51;
   wire n_2_52;
   wire n_2_54;
   wire n_2_55;
   wire n_2_57;
   wire n_2_58;
   wire n_2_61;
   wire n_2_62;
   wire n_2_81;
   wire n_2_82;
   wire n_2_84;
   wire n_2_85;
   wire n_2_87;
   wire n_2_88;
   wire n_2_95;
   wire n_2_98;
   wire n_2_99;
   wire n_2_114;
   wire n_2_115;
   wire n_2_117;
   wire n_2_118;
   wire n_2_124;
   wire n_2_125;
   wire n_2_130;
   wire n_2_131;
   wire n_2_151;
   wire n_2_152;
   wire n_2_154;
   wire n_2_155;
   wire n_2_158;
   wire n_2_159;
   wire n_2_169;
   wire n_2_170;
   wire n_2_181;
   wire n_2_182;
   wire n_2_186;
   wire n_2_187;
   wire n_2_189;
   wire n_2_190;
   wire n_2_199;
   wire n_2_200;
   wire n_2_206;
   wire n_2_8;
   wire n_2_349_0;
   wire n_2_349_1;
   wire n_2_16;
   wire n_2_350_0;
   wire n_2_350_1;
   wire n_2_20;
   wire n_2_351_0;
   wire n_2_351_1;
   wire n_2_26;
   wire n_2_352_0;
   wire n_2_352_1;
   wire n_2_27;
   wire n_2_353_0;
   wire n_2_353_1;
   wire n_2_59;
   wire n_2_354_0;
   wire n_2_354_1;
   wire n_2_63;
   wire n_2_355_0;
   wire n_2_355_1;
   wire n_2_74;
   wire n_2_356_0;
   wire n_2_356_1;
   wire n_2_108;
   wire n_2_357_0;
   wire n_2_357_1;
   wire n_2_109;
   wire n_2_358_0;
   wire n_2_358_1;
   wire n_2_164;
   wire n_2_359_0;
   wire n_2_359_1;
   wire n_2_360_0;
   wire n_2_360_1;
   wire n_2_204;
   wire n_2_361_0;
   wire n_2_361_1;
   wire n_2_195;
   wire n_2_362_0;
   wire n_2_362_1;
   wire n_2_193;
   wire n_2_363_0;
   wire n_2_363_1;
   wire n_2_178;
   wire n_2_364_0;
   wire n_2_364_1;
   wire n_2_175;
   wire n_2_365_0;
   wire n_2_365_1;
   wire n_2_171;
   wire n_2_366_0;
   wire n_2_366_1;
   wire n_2_147;
   wire n_2_367_0;
   wire n_2_367_1;
   wire n_2_143;
   wire n_2_368_0;
   wire n_2_368_1;
   wire n_2_139;
   wire n_2_369_0;
   wire n_2_369_1;
   wire n_2_135;
   wire n_2_370_0;
   wire n_2_370_1;
   wire n_2_132;
   wire n_2_371_0;
   wire n_2_371_1;
   wire n_2_107;
   wire n_2_372_0;
   wire n_2_372_1;
   wire n_2_105;
   wire n_2_373_0;
   wire n_2_373_1;
   wire n_2_103;
   wire n_2_374_0;
   wire n_2_374_1;
   wire n_2_101;
   wire n_2_375_0;
   wire n_2_375_1;
   wire n_2_96;
   wire n_2_376_0;
   wire n_2_376_1;
   wire n_2_92;
   wire n_2_377_0;
   wire n_2_377_1;
   wire n_2_79;
   wire n_2_378_0;
   wire n_2_378_1;
   wire n_2_73;
   wire n_2_379_0;
   wire n_2_379_1;
   wire n_2_72;
   wire n_2_380_0;
   wire n_2_380_1;
   wire n_2_44;
   wire n_2_381_0;
   wire n_2_381_1;
   wire n_2_35;
   wire n_2_382_0;
   wire n_2_382_1;
   wire n_2_9;
   wire n_2_383_0;
   wire n_2_383_1;
   wire n_2_146;
   wire n_2_384_0;
   wire n_2_384_1;
   wire n_2_64;
   wire n_2_385_0;
   wire n_2_385_1;
   wire n_2_47;
   wire n_2_386_0;
   wire n_2_386_1;
   wire n_2_41;
   wire n_2_387_0;
   wire n_2_387_1;
   wire n_2_32;
   wire n_2_388_0;
   wire n_2_388_1;
   wire n_2_31;
   wire n_2_389_0;
   wire n_2_389_1;
   wire n_2_25;
   wire n_2_390_0;
   wire n_2_390_1;
   wire n_2_192;
   wire n_2_391_0;
   wire n_2_391_1;
   wire n_2_191;
   wire n_2_392_0;
   wire n_2_392_1;
   wire n_2_183;
   wire n_2_393_0;
   wire n_2_393_1;
   wire n_2_106;
   wire n_2_394_0;
   wire n_2_394_1;
   wire n_2_13;
   wire n_2_395_0;
   wire n_2_395_1;
   wire n_2_10;
   wire n_2_396_0;
   wire n_2_396_1;
   wire n_2_207;
   wire n_2_397_0;
   wire n_2_397_1;
   wire n_2_179;
   wire n_2_398_0;
   wire n_2_398_1;
   wire n_2_298;
   wire n_2_360;
   wire n_2_340;
   wire n_2_341;
   wire n_2_342;
   wire n_2_343;
   wire n_2_344;
   wire n_2_345;
   wire [6:0]\out_as[0] ;
   wire n_2_361;
   wire n_2_346;
   wire n_2_347;
   wire n_2_370;
   wire n_2_372;
   wire n_2_362;
   wire n_2_348;
   wire [6:0]\out_as[1] ;
   wire [6:0]\out_bs[2] ;
   wire n_2_349;
   wire n_2_350;
   wire n_2_351;
   wire n_2_352;
   wire n_2_353;
   wire n_2_354;
   wire [6:0]\out_as[2] ;
   wire [6:0]\out_bs[3] ;
   wire n_2_363;
   wire n_2_355;
   wire n_2_364;
   wire n_2_356;
   wire n_2_357;
   wire n_2_358;
   wire [6:0]\out_as[3] ;
   wire [6:0]\out_bs[4] ;
   wire n_2_299;
   wire n_2_365;
   wire n_2_366;
   wire n_2_367;
   wire n_2_359;
   wire [6:0]\out_as[4] ;
   wire [6:0]\out_bs[5] ;
   wire [6:0]\out_as[5] ;
   wire n_2_399_0;
   wire n_2_400_0;
   wire n_2_400_1;
   wire n_2_400_2;
   wire n_2_400_3;
   wire n_2_401_0;
   wire n_2_401_1;
   wire n_2_402_0;
   wire n_2_402_1;
   wire n_2_403_0;
   wire n_2_403_1;
   wire n_2_404_0;
   wire n_2_404_1;
   wire n_2_405_0;
   wire n_2_405_1;
   wire n_2_406_0;
   wire n_2_406_1;
   wire n_2_407_0;
   wire n_2_407_1;
   wire n_2_408_0;
   wire n_2_408_1;
   wire n_2_409_0;
   wire n_2_409_1;
   wire n_2_410_0;
   wire n_2_410_1;
   wire n_2_411_0;
   wire n_2_411_1;
   wire n_2_412_0;
   wire n_2_412_1;
   wire n_2_413_0;
   wire n_2_413_1;
   wire n_2_414_0;
   wire n_2_414_1;
   wire n_2_415_0;
   wire n_2_415_1;
   wire n_2_416_0;
   wire n_2_416_1;
   wire n_2_417_0;
   wire n_2_417_1;
   wire n_2_418_0;
   wire n_2_418_1;
   wire n_2_419_0;
   wire n_2_419_1;
   wire n_2_420_0;
   wire n_2_420_1;
   wire n_2_421_0;
   wire n_2_421_1;
   wire n_2_422_0;
   wire n_2_422_1;
   wire n_2_423_0;
   wire n_2_423_1;
   wire n_2_424_0;
   wire n_2_424_1;
   wire n_2_425_0;
   wire n_2_425_1;
   wire n_2_426_0;
   wire n_2_426_1;
   wire n_2_427_0;
   wire n_2_427_1;
   wire n_2_428_0;
   wire n_2_428_1;
   wire n_2_429_0;
   wire n_2_429_1;
   wire n_2_430_0;
   wire n_2_430_1;
   wire n_2_431_0;
   wire n_2_431_1;
   wire n_2_432_0;
   wire n_2_432_1;
   wire n_2_433_0;
   wire n_2_433_1;
   wire n_2_434_0;
   wire n_2_434_1;
   wire n_2_435_0;
   wire n_2_435_1;
   wire n_2_436_0;
   wire n_2_436_1;
   wire n_2_437_0;
   wire n_2_437_1;
   wire n_2_438_0;
   wire n_2_438_1;
   wire n_2_439_0;
   wire n_2_439_1;
   wire n_2_440_0;
   wire n_2_440_1;
   wire n_2_441_0;
   wire n_2_441_1;
   wire n_2_442_0;
   wire n_2_442_1;
   wire n_2_443_0;
   wire n_2_443_1;
   wire n_2_444_0;
   wire n_2_444_1;
   wire n_2_445_0;
   wire n_2_445_1;
   wire n_2_446_0;
   wire n_2_446_1;
   wire n_2_447_0;
   wire n_2_447_1;
   wire n_2_448_0;
   wire n_2_448_1;
   wire n_2_449_0;
   wire n_2_449_1;
   wire n_2_450_0;
   wire n_2_450_1;
   wire n_2_451_0;
   wire n_2_451_1;
   wire n_2_452_0;
   wire n_2_452_1;
   wire n_2_453_0;
   wire n_2_453_1;
   wire n_2_11;
   wire n_2_12;
   wire n_2_14;
   wire n_2_15;
   wire n_2_33;
   wire n_2_34;
   wire n_2_36;
   wire n_2_37;
   wire n_2_42;
   wire n_2_43;
   wire n_2_45;
   wire n_2_46;
   wire n_2_65;
   wire n_2_66;
   wire n_2_110;
   wire n_2_111;
   wire n_2_133;
   wire n_2_134;
   wire n_2_136;
   wire n_2_137;
   wire n_2_140;
   wire n_2_141;
   wire n_2_144;
   wire n_2_145;
   wire n_2_148;
   wire n_2_149;
   wire n_2_480_0;
   wire n_2_480_1;
   wire n_2_176;
   wire n_2_177;
   wire n_2_165;
   wire n_2_166;
   wire n_2_485_0;
   wire n_2_485_1;
   wire n_2_485_2;
   wire n_2_48;
   wire n_2_49;
   wire n_2_229;
   wire n_2_230;
   wire n_2_231;
   wire n_2_238;
   wire n_2_242;
   wire n_2_243;
   wire n_2_249;
   wire n_2_252;
   wire n_2_256;
   wire n_2_257;
   wire n_2_258;
   wire n_2_260;
   wire n_2_264;
   wire n_2_265;
   wire n_2_266;
   wire n_2_267;
   wire n_2_269;
   wire n_2_270;
   wire n_2_271;
   wire n_2_272;
   wire n_2_278;
   wire n_2_279;
   wire n_2_280;
   wire n_2_281;
   wire n_2_283;
   wire n_2_285;
   wire n_2_286;
   wire n_2_287;
   wire n_2_288;
   wire n_2_289;
   wire n_2_290;
   wire n_2_291;
   wire n_2_523_0;
   wire n_2_523_1;
   wire n_2_232;
   wire n_2_525_0;
   wire n_2_525_1;
   wire n_2_292;
   wire n_2_528_0;
   wire n_2_528_1;
   wire n_2_236;
   wire n_2_530_0;
   wire n_2_530_1;
   wire n_2_293;
   wire n_2_533_0;
   wire n_2_533_1;
   wire n_2_239;
   wire n_2_535_0;
   wire n_2_535_1;
   wire n_2_294;
   wire n_2_538_0;
   wire n_2_538_1;
   wire n_2_539_0;
   wire n_2_539_1;
   wire n_2_247;
   wire n_2_541_0;
   wire n_2_541_1;
   wire n_2_544_0;
   wire n_2_544_1;
   wire n_2_261;
   wire n_2_546_0;
   wire n_2_546_1;
   wire n_2_297;
   wire buf_is_empty;
   wire n_2_300;
   wire n_2_301;
   wire n_2_549_0;
   wire n_2_549_1;
   wire n_2_302;
   wire n_2_549_2;
   wire n_2_549_3;
   wire n_2_303;
   wire n_2_549_4;
   wire n_2_549_5;
   wire n_2_304;
   wire n_2_549_6;
   wire n_2_549_7;
   wire n_2_305;
   wire n_2_549_8;
   wire n_2_549_9;
   wire n_2_306;
   wire n_2_549_10;
   wire n_2_549_11;
   wire n_2_307;
   wire n_2_549_12;
   wire n_2_549_13;
   wire n_2_308;
   wire n_2_549_14;
   wire n_2_549_15;
   wire n_2_309;
   wire n_2_549_16;
   wire n_2_549_17;
   wire n_2_310;
   wire n_2_549_18;
   wire n_2_549_19;
   wire n_2_311;
   wire n_2_549_20;
   wire n_2_549_21;
   wire n_2_312;
   wire n_2_549_22;
   wire n_2_549_23;
   wire n_2_313;
   wire n_2_549_24;
   wire n_2_549_25;
   wire n_2_314;
   wire n_2_549_26;
   wire n_2_549_27;
   wire n_2_315;
   wire n_2_549_28;
   wire n_2_549_29;
   wire n_2_316;
   wire n_2_549_30;
   wire n_2_549_31;
   wire n_2_317;
   wire n_2_549_32;
   wire n_2_549_33;
   wire n_2_318;
   wire n_2_549_34;
   wire n_2_549_35;
   wire n_2_319;
   wire n_2_549_36;
   wire n_2_549_37;
   wire n_2_320;
   wire n_2_549_38;
   wire n_2_549_39;
   wire n_2_321;
   wire n_2_549_40;
   wire n_2_549_41;
   wire n_2_322;
   wire n_2_549_42;
   wire n_2_549_43;
   wire n_2_323;
   wire n_2_549_44;
   wire n_2_549_45;
   wire n_2_324;
   wire n_2_549_46;
   wire n_2_549_47;
   wire n_2_325;
   wire n_2_549_48;
   wire n_2_549_49;
   wire n_2_326;
   wire n_2_549_50;
   wire n_2_549_51;
   wire n_2_327;
   wire n_2_549_52;
   wire n_2_549_53;
   wire n_2_328;
   wire n_2_549_54;
   wire n_2_549_55;
   wire n_2_329;
   wire n_2_549_56;
   wire n_2_549_57;
   wire n_2_330;
   wire n_2_549_58;
   wire n_2_549_59;
   wire n_2_331;
   wire n_2_549_60;
   wire n_2_549_61;
   wire n_2_332;
   wire n_2_549_62;
   wire n_2_549_63;
   wire n_2_549_64;
   wire n_2_549_65;
   wire n_2_549_66;
   wire n_2_333;
   wire n_2_549_67;
   wire n_2_334;
   wire n_2_549_68;
   wire n_2_549_69;
   wire n_2_549_70;
   wire n_2_549_71;
   wire n_2_549_72;
   wire n_2_549_73;
   wire n_2_549_74;
   wire n_2_549_75;
   wire n_2_549_76;
   wire n_2_549_77;
   wire n_2_373;
   wire n_2_549_78;
   wire n_2_549_79;
   wire [6:0]buf_fill_flush_diff;
   wire n_2_245;
   wire n_2_295;
   wire n_2_234;
   wire n_2_235;
   wire n_2_250;
   wire n_2_251;
   wire n_2_253;
   wire n_2_254;
   wire n_2_263;
   wire n_2_268;
   wire n_2_273;
   wire n_2_274;
   wire n_2_275;
   wire n_2_276;
   wire n_2_277;
   wire n_2_284;
   wire n_2_282;
   wire n_2_255;
   wire n_2_262;
   wire n_2_246;
   wire n_2_244;
   wire n_2_240;
   wire n_2_237;
   wire n_2_233;
   wire n_2_259;
   wire n_2_248;
   wire error_success_reg_enable_mux_n_0;
   wire n_2_335;
   wire [6:0]buf_flush_i_inc;
   wire [6:0]buf_flush_i_inv;
   wire [6:0]buf_fill_i;
   wire n_2_336;
   wire [6:0]buf_flush_i;
   wire n_2_337;
   wire n_2_338;
   wire [6:0]\out_bs[0] ;
   wire [6:0]\out_bs[1] ;
   wire n_2_368;
   wire n_2_369;
   wire n_2_371;
   wire n_2_542_0;
   wire n_2_542_1;
   wire n_2_296;
   wire n_2_542_2;
   wire n_2_542_3;
   wire n_2_542_4;

   datapath__1_13515 i_58_58 (.to_int6128({1'b0, \out_as[7] [6], \out_as[7] [5], 
      \out_as[7] [4], \out_as[7] [3], \out_as[7] [2], \out_as[7] [1], 1'b0}), 
      .p_0(n_0));
   datapath__1_13522 i_58_64 (.to_int6128({1'b0, \out_as[7] [6], \out_as[7] [5], 
      \out_as[7] [4], \out_as[7] [3], \out_as[7] [2], 1'b0, 1'b0}), .p_0(n_1));
   range_extractor__3_461 ranges_6_range_extr_i (.in_a(\out_bs[5] ), .in_size({
      in_data[7], in_data[6], in_data[5]}), .out_a(\out_as[6] ), .out_b(
      \out_bs[6] ));
   HA_X1 i_1_737_0 (.A(\out_as[7] [6]), .B(n_1_737_1301), .CO(n_1_737_0), .S());
   HA_X1 i_1_737_1 (.A(\out_as[7] [6]), .B(n_1_737_1300), .CO(n_1_737_1), .S());
   HA_X1 i_1_737_2 (.A(\out_as[7] [6]), .B(n_1_737_5141), .CO(n_1_737_2), .S());
   HA_X1 i_1_737_3 (.A(\out_as[7] [6]), .B(n_1_737_1299), .CO(n_1_737_3), .S());
   HA_X1 i_1_737_4 (.A(\out_as[7] [6]), .B(n_1_737_1298), .CO(n_1_737_4), .S());
   HA_X1 i_1_737_5 (.A(\out_as[7] [6]), .B(n_1_737_1297), .CO(n_1_737_5), .S());
   HA_X1 i_1_737_6 (.A(\out_as[7] [6]), .B(n_1_737_5138), .CO(n_1_737_6), .S());
   HA_X1 i_1_737_7 (.A(\out_as[7] [6]), .B(n_1_737_1296), .CO(n_1_737_7), .S());
   HA_X1 i_1_737_8 (.A(\out_as[7] [6]), .B(n_1_737_1295), .CO(n_1_737_8), .S());
   HA_X1 i_1_737_9 (.A(\out_as[7] [6]), .B(n_1_737_1294), .CO(n_1_737_9), .S());
   HA_X1 i_1_737_10 (.A(\out_as[7] [6]), .B(n_1_737_1293), .CO(n_1_737_10), 
      .S());
   HA_X1 i_1_737_11 (.A(\out_as[7] [6]), .B(n_1_737_1292), .CO(n_1_737_11), 
      .S());
   HA_X1 i_1_737_12 (.A(\out_as[7] [6]), .B(n_1_737_1291), .CO(n_1_737_12), 
      .S());
   HA_X1 i_1_737_13 (.A(\out_as[7] [6]), .B(n_1_737_1290), .CO(n_1_737_13), 
      .S());
   HA_X1 i_1_737_14 (.A(\out_as[7] [6]), .B(n_1_737_5142), .CO(n_1_737_14), 
      .S());
   HA_X1 i_1_737_15 (.A(\out_as[7] [6]), .B(n_1_737_1289), .CO(n_1_737_15), 
      .S());
   HA_X1 i_1_737_16 (.A(\out_as[7] [6]), .B(n_1_737_1288), .CO(n_1_737_16), 
      .S());
   HA_X1 i_1_737_17 (.A(\out_as[7] [6]), .B(n_1_737_1287), .CO(n_1_737_17), 
      .S());
   HA_X1 i_1_737_18 (.A(\out_as[7] [6]), .B(n_1_737_1286), .CO(n_1_737_18), 
      .S());
   HA_X1 i_1_737_19 (.A(\out_as[7] [6]), .B(n_1_737_1285), .CO(n_1_737_19), 
      .S());
   HA_X1 i_1_737_20 (.A(\out_as[7] [6]), .B(n_1_737_1284), .CO(n_1_737_20), 
      .S());
   HA_X1 i_1_737_21 (.A(\out_as[7] [6]), .B(n_1_737_1283), .CO(n_1_737_21), 
      .S());
   HA_X1 i_1_737_22 (.A(\out_as[7] [6]), .B(n_1_737_1282), .CO(n_1_737_22), 
      .S());
   HA_X1 i_1_737_23 (.A(\out_as[7] [6]), .B(n_1_737_1281), .CO(n_1_737_23), 
      .S());
   HA_X1 i_1_737_24 (.A(\out_as[7] [6]), .B(n_1_737_1280), .CO(n_1_737_24), 
      .S());
   HA_X1 i_1_737_25 (.A(\out_as[7] [6]), .B(n_1_737_1279), .CO(n_1_737_25), 
      .S());
   HA_X1 i_1_737_26 (.A(\out_as[7] [6]), .B(n_1_737_1278), .CO(n_1_737_26), 
      .S());
   HA_X1 i_1_737_27 (.A(\out_as[7] [6]), .B(n_1_737_1277), .CO(n_1_737_27), 
      .S());
   HA_X1 i_1_737_28 (.A(\out_as[7] [6]), .B(n_1_737_1276), .CO(n_1_737_28), 
      .S());
   HA_X1 i_1_737_29 (.A(\out_as[7] [6]), .B(n_1_737_1275), .CO(n_1_737_29), 
      .S());
   HA_X1 i_1_737_30 (.A(\out_as[7] [6]), .B(\out_as[7] [5]), .CO(n_1_737_30), 
      .S());
   HA_X1 i_1_737_31 (.A(\out_as[7] [5]), .B(n_1_737_2020), .CO(n_1_737_31), 
      .S());
   HA_X1 i_1_737_32 (.A(\out_as[7] [6]), .B(n_1_737_31), .CO(n_1_737_32), .S());
   HA_X1 i_1_737_33 (.A(\out_as[7] [5]), .B(n_1_737_1302), .CO(n_1_737_33), 
      .S());
   HA_X1 i_1_737_34 (.A(\out_as[7] [6]), .B(n_1_737_33), .CO(n_1_737_34), .S());
   HA_X1 i_1_737_35 (.A(\out_as[7] [5]), .B(n_1_737_1274), .CO(n_1_737_35), 
      .S());
   HA_X1 i_1_737_36 (.A(\out_as[7] [6]), .B(n_1_737_35), .CO(n_1_737_36), .S());
   HA_X1 i_1_737_37 (.A(\out_as[7] [5]), .B(n_1_737_5143), .CO(n_1_737_37), 
      .S());
   HA_X1 i_1_737_38 (.A(\out_as[7] [6]), .B(n_1_737_37), .CO(n_1_737_38), .S());
   HA_X1 i_1_737_39 (.A(\out_as[7] [5]), .B(n_1_737_1273), .CO(n_1_737_39), 
      .S());
   HA_X1 i_1_737_40 (.A(\out_as[7] [6]), .B(n_1_737_39), .CO(n_1_737_40), .S());
   HA_X1 i_1_737_41 (.A(\out_as[7] [5]), .B(n_1_737_1272), .CO(n_1_737_41), 
      .S());
   HA_X1 i_1_737_42 (.A(\out_as[7] [6]), .B(n_1_737_41), .CO(n_1_737_42), .S());
   HA_X1 i_1_737_43 (.A(\out_as[7] [5]), .B(n_1_737_1271), .CO(n_1_737_43), 
      .S());
   HA_X1 i_1_737_44 (.A(\out_as[7] [6]), .B(n_1_737_43), .CO(n_1_737_44), .S());
   HA_X1 i_1_737_45 (.A(\out_as[7] [5]), .B(n_1_737_5144), .CO(n_1_737_45), 
      .S());
   HA_X1 i_1_737_46 (.A(\out_as[7] [6]), .B(n_1_737_45), .CO(n_1_737_46), .S());
   HA_X1 i_1_737_47 (.A(\out_as[7] [5]), .B(n_1_737_1270), .CO(n_1_737_47), 
      .S());
   HA_X1 i_1_737_48 (.A(\out_as[7] [6]), .B(n_1_737_47), .CO(n_1_737_48), .S());
   HA_X1 i_1_737_49 (.A(\out_as[7] [5]), .B(n_1_737_1269), .CO(n_1_737_49), 
      .S());
   HA_X1 i_1_737_50 (.A(\out_as[7] [6]), .B(n_1_737_49), .CO(n_1_737_50), .S());
   HA_X1 i_1_737_51 (.A(\out_as[7] [5]), .B(n_1_737_1268), .CO(n_1_737_51), 
      .S());
   HA_X1 i_1_737_52 (.A(\out_as[7] [6]), .B(n_1_737_51), .CO(n_1_737_52), .S());
   HA_X1 i_1_737_53 (.A(\out_as[7] [5]), .B(n_1_737_1267), .CO(n_1_737_53), 
      .S());
   HA_X1 i_1_737_54 (.A(\out_as[7] [6]), .B(n_1_737_53), .CO(n_1_737_54), .S());
   HA_X1 i_1_737_55 (.A(\out_as[7] [5]), .B(n_1_737_1266), .CO(n_1_737_55), 
      .S());
   HA_X1 i_1_737_56 (.A(\out_as[7] [6]), .B(n_1_737_55), .CO(n_1_737_56), .S());
   HA_X1 i_1_737_57 (.A(\out_as[7] [5]), .B(n_1_737_1265), .CO(n_1_737_57), 
      .S());
   HA_X1 i_1_737_58 (.A(\out_as[7] [6]), .B(n_1_737_57), .CO(n_1_737_58), .S());
   HA_X1 i_1_737_59 (.A(\out_as[7] [5]), .B(n_1_737_1264), .CO(n_1_737_59), 
      .S());
   HA_X1 i_1_737_60 (.A(\out_as[7] [6]), .B(n_1_737_59), .CO(n_1_737_60), .S());
   HA_X1 i_1_737_61 (.A(\out_as[7] [5]), .B(\out_as[7] [4]), .CO(n_1_737_61), 
      .S());
   HA_X1 i_1_737_62 (.A(\out_as[7] [6]), .B(n_1_737_61), .CO(n_1_737_62), .S());
   HA_X1 i_1_737_63 (.A(\out_as[7] [4]), .B(n_1_737_2021), .CO(n_1_737_63), 
      .S());
   HA_X1 i_1_737_64 (.A(\out_as[7] [5]), .B(n_1_737_63), .CO(n_1_737_64), .S());
   HA_X1 i_1_737_65 (.A(\out_as[7] [6]), .B(n_1_737_64), .CO(n_1_737_65), .S());
   HA_X1 i_1_737_66 (.A(\out_as[7] [4]), .B(n_1_737_2024), .CO(n_1_737_66), 
      .S());
   HA_X1 i_1_737_67 (.A(\out_as[7] [5]), .B(n_1_737_66), .CO(n_1_737_67), .S());
   HA_X1 i_1_737_68 (.A(\out_as[7] [6]), .B(n_1_737_67), .CO(n_1_737_68), .S());
   HA_X1 i_1_737_69 (.A(\out_as[7] [4]), .B(n_1_737_1263), .CO(n_1_737_69), 
      .S());
   HA_X1 i_1_737_70 (.A(\out_as[7] [5]), .B(n_1_737_69), .CO(n_1_737_70), .S());
   HA_X1 i_1_737_71 (.A(\out_as[7] [6]), .B(n_1_737_70), .CO(n_1_737_71), .S());
   HA_X1 i_1_737_72 (.A(\out_as[7] [4]), .B(n_1_737_5145), .CO(n_1_737_72), 
      .S());
   HA_X1 i_1_737_73 (.A(\out_as[7] [5]), .B(n_1_737_72), .CO(n_1_737_73), .S());
   HA_X1 i_1_737_74 (.A(\out_as[7] [6]), .B(n_1_737_73), .CO(n_1_737_74), .S());
   HA_X1 i_1_737_75 (.A(\out_as[7] [4]), .B(n_1_737_1262), .CO(n_1_737_75), 
      .S());
   HA_X1 i_1_737_76 (.A(\out_as[7] [5]), .B(n_1_737_75), .CO(n_1_737_76), .S());
   HA_X1 i_1_737_77 (.A(\out_as[7] [6]), .B(n_1_737_76), .CO(n_1_737_77), .S());
   HA_X1 i_1_737_78 (.A(\out_as[7] [4]), .B(n_1_737_1261), .CO(n_1_737_78), 
      .S());
   HA_X1 i_1_737_79 (.A(\out_as[7] [5]), .B(n_1_737_78), .CO(n_1_737_79), .S());
   HA_X1 i_1_737_80 (.A(\out_as[7] [6]), .B(n_1_737_79), .CO(n_1_737_80), .S());
   HA_X1 i_1_737_81 (.A(\out_as[7] [4]), .B(n_1_737_1260), .CO(n_1_737_81), 
      .S());
   HA_X1 i_1_737_82 (.A(\out_as[7] [5]), .B(n_1_737_81), .CO(n_1_737_82), .S());
   HA_X1 i_1_737_83 (.A(\out_as[7] [6]), .B(n_1_737_82), .CO(n_1_737_83), .S());
   HA_X1 i_1_737_84 (.A(\out_as[7] [4]), .B(\out_as[7] [3]), .CO(n_1_737_84), 
      .S());
   HA_X1 i_1_737_85 (.A(\out_as[7] [5]), .B(n_1_737_84), .CO(n_1_737_85), .S());
   HA_X1 i_1_737_86 (.A(\out_as[7] [6]), .B(n_1_737_85), .CO(n_1_737_86), .S());
   HA_X1 i_1_737_87 (.A(\out_as[7] [3]), .B(n_1_737_2022), .CO(n_1_737_87), 
      .S());
   HA_X1 i_1_737_88 (.A(\out_as[7] [4]), .B(n_1_737_87), .CO(n_1_737_88), .S());
   HA_X1 i_1_737_89 (.A(\out_as[7] [5]), .B(n_1_737_88), .CO(n_1_737_89), .S());
   HA_X1 i_1_737_90 (.A(\out_as[7] [6]), .B(n_1_737_89), .CO(n_1_737_90), .S());
   HA_X1 i_1_737_91 (.A(\out_as[7] [3]), .B(n_1_737_2025), .CO(n_1_737_91), 
      .S());
   HA_X1 i_1_737_92 (.A(\out_as[7] [4]), .B(n_1_737_91), .CO(n_1_737_92), .S());
   HA_X1 i_1_737_93 (.A(\out_as[7] [5]), .B(n_1_737_92), .CO(n_1_737_93), .S());
   HA_X1 i_1_737_94 (.A(\out_as[7] [6]), .B(n_1_737_93), .CO(n_1_737_94), .S());
   HA_X1 i_1_737_95 (.A(\out_as[7] [3]), .B(n_1_737_1259), .CO(n_1_737_95), 
      .S());
   HA_X1 i_1_737_96 (.A(\out_as[7] [4]), .B(n_1_737_95), .CO(n_1_737_96), .S());
   HA_X1 i_1_737_97 (.A(\out_as[7] [5]), .B(n_1_737_96), .CO(n_1_737_97), .S());
   HA_X1 i_1_737_98 (.A(\out_as[7] [6]), .B(n_1_737_97), .CO(n_1_737_98), .S());
   HA_X1 i_1_737_99 (.A(\out_as[7] [3]), .B(\out_as[7] [2]), .CO(n_1_737_99), 
      .S());
   HA_X1 i_1_737_100 (.A(\out_as[7] [4]), .B(n_1_737_99), .CO(n_1_737_100), 
      .S());
   HA_X1 i_1_737_101 (.A(\out_as[7] [5]), .B(n_1_737_100), .CO(n_1_737_101), 
      .S());
   HA_X1 i_1_737_102 (.A(\out_as[7] [6]), .B(n_1_737_101), .CO(n_1_737_102), 
      .S());
   HA_X1 i_1_737_103 (.A(\out_as[7] [2]), .B(n_1_737_2023), .CO(n_1_737_103), 
      .S());
   HA_X1 i_1_737_104 (.A(\out_as[7] [3]), .B(n_1_737_103), .CO(n_1_737_104), 
      .S());
   HA_X1 i_1_737_105 (.A(\out_as[7] [4]), .B(n_1_737_104), .CO(n_1_737_105), 
      .S());
   HA_X1 i_1_737_106 (.A(\out_as[7] [5]), .B(n_1_737_105), .CO(n_1_737_106), 
      .S());
   HA_X1 i_1_737_107 (.A(\out_as[7] [6]), .B(n_1_737_106), .CO(n_1_737_107), 
      .S());
   HA_X1 i_1_737_108 (.A(\out_as[7] [2]), .B(\out_as[7] [1]), .CO(n_1_737_108), 
      .S());
   HA_X1 i_1_737_109 (.A(\out_as[7] [3]), .B(n_1_737_108), .CO(n_1_737_109), 
      .S());
   HA_X1 i_1_737_110 (.A(\out_as[7] [4]), .B(n_1_737_109), .CO(n_1_737_110), 
      .S());
   HA_X1 i_1_737_111 (.A(\out_as[7] [5]), .B(n_1_737_110), .CO(n_1_737_111), 
      .S());
   HA_X1 i_1_737_112 (.A(\out_as[7] [6]), .B(n_1_737_111), .CO(n_1_737_112), 
      .S());
   HA_X1 i_1_737_113 (.A(\out_as[7] [1]), .B(\out_as[7] [0]), .CO(n_1_737_113), 
      .S());
   HA_X1 i_1_737_114 (.A(\out_as[7] [2]), .B(n_1_737_113), .CO(n_1_737_114), 
      .S());
   HA_X1 i_1_737_115 (.A(\out_as[7] [3]), .B(n_1_737_114), .CO(n_1_737_115), 
      .S());
   HA_X1 i_1_737_116 (.A(\out_as[7] [4]), .B(n_1_737_115), .CO(n_1_737_116), 
      .S());
   HA_X1 i_1_737_117 (.A(\out_as[7] [5]), .B(n_1_737_116), .CO(n_1_737_117), 
      .S());
   HA_X1 i_1_737_118 (.A(\out_as[7] [6]), .B(n_1_737_117), .CO(n_1_737_118), 
      .S());
   HA_X1 i_1_737_119 (.A(\out_as[0] [1]), .B(\out_as[0] [0]), .CO(n_1_737_119), 
      .S());
   HA_X1 i_1_737_120 (.A(\out_as[1] [1]), .B(\out_as[1] [0]), .CO(n_1_737_120), 
      .S());
   HA_X1 i_1_737_121 (.A(\out_as[2] [1]), .B(\out_as[2] [0]), .CO(n_1_737_121), 
      .S());
   HA_X1 i_1_737_122 (.A(\out_as[3] [1]), .B(\out_as[3] [0]), .CO(n_1_737_122), 
      .S());
   HA_X1 i_1_737_123 (.A(\out_as[4] [1]), .B(\out_as[4] [0]), .CO(n_1_737_123), 
      .S());
   HA_X1 i_1_737_124 (.A(\out_as[5] [1]), .B(\out_as[5] [0]), .CO(n_1_737_124), 
      .S());
   HA_X1 i_1_737_125 (.A(\out_as[6] [1]), .B(\out_as[6] [0]), .CO(n_1_737_125), 
      .S());
   HA_X1 i_1_737_126 (.A(\out_as[0] [2]), .B(n_1_737_2008), .CO(n_1_737_126), 
      .S());
   HA_X1 i_1_737_127 (.A(\out_as[1] [2]), .B(n_1_737_1997), .CO(n_1_737_127), 
      .S());
   HA_X1 i_1_737_128 (.A(\out_as[2] [2]), .B(n_1_737_1991), .CO(n_1_737_128), 
      .S());
   HA_X1 i_1_737_129 (.A(\out_as[3] [2]), .B(n_1_737_2019), .CO(n_1_737_129), 
      .S());
   HA_X1 i_1_737_130 (.A(\out_as[4] [2]), .B(n_1_737_2002), .CO(n_1_737_130), 
      .S());
   HA_X1 i_1_737_131 (.A(\out_as[5] [2]), .B(n_1_737_2013), .CO(n_1_737_131), 
      .S());
   HA_X1 i_1_737_132 (.A(\out_as[6] [2]), .B(n_1_737_1984), .CO(n_1_737_132), 
      .S());
   HA_X1 i_1_737_133 (.A(\out_as[0] [2]), .B(\out_as[0] [1]), .CO(n_1_737_133), 
      .S());
   HA_X1 i_1_737_134 (.A(\out_as[1] [2]), .B(\out_as[1] [1]), .CO(n_1_737_134), 
      .S());
   HA_X1 i_1_737_135 (.A(\out_as[2] [2]), .B(\out_as[2] [1]), .CO(n_1_737_135), 
      .S());
   HA_X1 i_1_737_136 (.A(\out_as[3] [2]), .B(\out_as[3] [1]), .CO(n_1_737_136), 
      .S());
   HA_X1 i_1_737_137 (.A(\out_as[4] [2]), .B(\out_as[4] [1]), .CO(n_1_737_137), 
      .S());
   HA_X1 i_1_737_138 (.A(\out_as[5] [2]), .B(\out_as[5] [1]), .CO(n_1_737_138), 
      .S());
   HA_X1 i_1_737_139 (.A(\out_as[6] [2]), .B(\out_as[6] [1]), .CO(n_1_737_139), 
      .S());
   HA_X1 i_1_737_140 (.A(\out_as[0] [2]), .B(n_1_737_119), .CO(n_1_737_140), 
      .S());
   HA_X1 i_1_737_141 (.A(\out_as[1] [2]), .B(n_1_737_120), .CO(n_1_737_141), 
      .S());
   HA_X1 i_1_737_142 (.A(\out_as[2] [2]), .B(n_1_737_121), .CO(n_1_737_142), 
      .S());
   HA_X1 i_1_737_143 (.A(\out_as[3] [2]), .B(n_1_737_122), .CO(n_1_737_143), 
      .S());
   HA_X1 i_1_737_144 (.A(\out_as[4] [2]), .B(n_1_737_123), .CO(n_1_737_144), 
      .S());
   HA_X1 i_1_737_145 (.A(\out_as[5] [2]), .B(n_1_737_124), .CO(n_1_737_145), 
      .S());
   HA_X1 i_1_737_146 (.A(\out_as[6] [2]), .B(n_1_737_125), .CO(n_1_737_146), 
      .S());
   HA_X1 i_1_737_147 (.A(\out_as[0] [3]), .B(n_1_737_2007), .CO(n_1_737_147), 
      .S());
   HA_X1 i_1_737_148 (.A(\out_as[1] [3]), .B(n_1_737_1996), .CO(n_1_737_148), 
      .S());
   HA_X1 i_1_737_149 (.A(\out_as[2] [3]), .B(n_1_737_1990), .CO(n_1_737_149), 
      .S());
   HA_X1 i_1_737_150 (.A(\out_as[3] [3]), .B(n_1_737_2018), .CO(n_1_737_150), 
      .S());
   HA_X1 i_1_737_151 (.A(\out_as[4] [3]), .B(n_1_737_2001), .CO(n_1_737_151), 
      .S());
   HA_X1 i_1_737_152 (.A(\out_as[5] [3]), .B(n_1_737_2012), .CO(n_1_737_152), 
      .S());
   HA_X1 i_1_737_153 (.A(\out_as[6] [3]), .B(n_1_737_1983), .CO(n_1_737_153), 
      .S());
   HA_X1 i_1_737_154 (.A(\out_as[0] [3]), .B(n_1_737_5361), .CO(n_1_737_154), 
      .S());
   HA_X1 i_1_737_155 (.A(\out_as[1] [3]), .B(n_1_737_5323), .CO(n_1_737_155), 
      .S());
   HA_X1 i_1_737_156 (.A(\out_as[2] [3]), .B(n_1_737_5277), .CO(n_1_737_156), 
      .S());
   HA_X1 i_1_737_157 (.A(\out_as[3] [3]), .B(n_1_737_5218), .CO(n_1_737_157), 
      .S());
   HA_X1 i_1_737_158 (.A(\out_as[4] [3]), .B(n_1_737_5389), .CO(n_1_737_158), 
      .S());
   HA_X1 i_1_737_159 (.A(\out_as[5] [3]), .B(n_1_737_5170), .CO(n_1_737_159), 
      .S());
   HA_X1 i_1_737_160 (.A(\out_as[6] [3]), .B(n_1_737_5157), .CO(n_1_737_160), 
      .S());
   HA_X1 i_1_737_161 (.A(\out_as[0] [3]), .B(n_1_737_1258), .CO(n_1_737_161), 
      .S());
   HA_X1 i_1_737_162 (.A(\out_as[1] [3]), .B(n_1_737_1257), .CO(n_1_737_162), 
      .S());
   HA_X1 i_1_737_163 (.A(\out_as[2] [3]), .B(n_1_737_1256), .CO(n_1_737_163), 
      .S());
   HA_X1 i_1_737_164 (.A(\out_as[3] [3]), .B(n_1_737_1255), .CO(n_1_737_164), 
      .S());
   HA_X1 i_1_737_165 (.A(\out_as[4] [3]), .B(n_1_737_1254), .CO(n_1_737_165), 
      .S());
   HA_X1 i_1_737_166 (.A(\out_as[5] [3]), .B(n_1_737_1253), .CO(n_1_737_166), 
      .S());
   HA_X1 i_1_737_167 (.A(\out_as[6] [3]), .B(n_1_737_1252), .CO(n_1_737_167), 
      .S());
   HA_X1 i_1_737_168 (.A(\out_as[0] [3]), .B(\out_as[0] [2]), .CO(n_1_737_168), 
      .S());
   HA_X1 i_1_737_169 (.A(\out_as[1] [3]), .B(\out_as[1] [2]), .CO(n_1_737_169), 
      .S());
   HA_X1 i_1_737_170 (.A(\out_as[2] [3]), .B(\out_as[2] [2]), .CO(n_1_737_170), 
      .S());
   HA_X1 i_1_737_171 (.A(\out_as[3] [3]), .B(\out_as[3] [2]), .CO(n_1_737_171), 
      .S());
   HA_X1 i_1_737_172 (.A(\out_as[4] [3]), .B(\out_as[4] [2]), .CO(n_1_737_172), 
      .S());
   HA_X1 i_1_737_173 (.A(\out_as[5] [3]), .B(\out_as[5] [2]), .CO(n_1_737_173), 
      .S());
   HA_X1 i_1_737_174 (.A(\out_as[6] [3]), .B(\out_as[6] [2]), .CO(n_1_737_174), 
      .S());
   HA_X1 i_1_737_175 (.A(\out_as[0] [3]), .B(n_1_737_126), .CO(n_1_737_175), 
      .S());
   HA_X1 i_1_737_176 (.A(\out_as[1] [3]), .B(n_1_737_127), .CO(n_1_737_176), 
      .S());
   HA_X1 i_1_737_177 (.A(\out_as[2] [3]), .B(n_1_737_128), .CO(n_1_737_177), 
      .S());
   HA_X1 i_1_737_178 (.A(\out_as[3] [3]), .B(n_1_737_129), .CO(n_1_737_178), 
      .S());
   HA_X1 i_1_737_179 (.A(\out_as[4] [3]), .B(n_1_737_130), .CO(n_1_737_179), 
      .S());
   HA_X1 i_1_737_180 (.A(\out_as[5] [3]), .B(n_1_737_131), .CO(n_1_737_180), 
      .S());
   HA_X1 i_1_737_181 (.A(\out_as[6] [3]), .B(n_1_737_132), .CO(n_1_737_181), 
      .S());
   HA_X1 i_1_737_182 (.A(\out_as[0] [3]), .B(n_1_737_133), .CO(n_1_737_182), 
      .S());
   HA_X1 i_1_737_183 (.A(\out_as[1] [3]), .B(n_1_737_134), .CO(n_1_737_183), 
      .S());
   HA_X1 i_1_737_184 (.A(\out_as[2] [3]), .B(n_1_737_135), .CO(n_1_737_184), 
      .S());
   HA_X1 i_1_737_185 (.A(\out_as[3] [3]), .B(n_1_737_136), .CO(n_1_737_185), 
      .S());
   HA_X1 i_1_737_186 (.A(\out_as[4] [3]), .B(n_1_737_137), .CO(n_1_737_186), 
      .S());
   HA_X1 i_1_737_187 (.A(\out_as[5] [3]), .B(n_1_737_138), .CO(n_1_737_187), 
      .S());
   HA_X1 i_1_737_188 (.A(\out_as[6] [3]), .B(n_1_737_139), .CO(n_1_737_188), 
      .S());
   HA_X1 i_1_737_189 (.A(\out_as[0] [3]), .B(n_1_737_140), .CO(n_1_737_189), 
      .S());
   HA_X1 i_1_737_190 (.A(\out_as[1] [3]), .B(n_1_737_141), .CO(n_1_737_190), 
      .S());
   HA_X1 i_1_737_191 (.A(\out_as[2] [3]), .B(n_1_737_142), .CO(n_1_737_191), 
      .S());
   HA_X1 i_1_737_192 (.A(\out_as[3] [3]), .B(n_1_737_143), .CO(n_1_737_192), 
      .S());
   HA_X1 i_1_737_193 (.A(\out_as[4] [3]), .B(n_1_737_144), .CO(n_1_737_193), 
      .S());
   HA_X1 i_1_737_194 (.A(\out_as[5] [3]), .B(n_1_737_145), .CO(n_1_737_194), 
      .S());
   HA_X1 i_1_737_195 (.A(\out_as[6] [3]), .B(n_1_737_146), .CO(n_1_737_195), 
      .S());
   HA_X1 i_1_737_196 (.A(\out_as[0] [4]), .B(n_1_737_2006), .CO(n_1_737_196), 
      .S());
   HA_X1 i_1_737_197 (.A(\out_as[1] [4]), .B(n_1_737_1995), .CO(n_1_737_197), 
      .S());
   HA_X1 i_1_737_198 (.A(\out_as[2] [4]), .B(n_1_737_1989), .CO(n_1_737_198), 
      .S());
   HA_X1 i_1_737_199 (.A(\out_as[3] [4]), .B(n_1_737_2017), .CO(n_1_737_199), 
      .S());
   HA_X1 i_1_737_200 (.A(\out_as[4] [4]), .B(n_1_737_2000), .CO(n_1_737_200), 
      .S());
   HA_X1 i_1_737_201 (.A(\out_as[5] [4]), .B(n_1_737_2011), .CO(n_1_737_201), 
      .S());
   HA_X1 i_1_737_202 (.A(\out_as[6] [4]), .B(n_1_737_1982), .CO(n_1_737_202), 
      .S());
   HA_X1 i_1_737_203 (.A(\out_as[0] [4]), .B(n_1_737_5350), .CO(n_1_737_203), 
      .S());
   HA_X1 i_1_737_204 (.A(\out_as[1] [4]), .B(n_1_737_5312), .CO(n_1_737_204), 
      .S());
   HA_X1 i_1_737_205 (.A(\out_as[2] [4]), .B(n_1_737_5268), .CO(n_1_737_205), 
      .S());
   HA_X1 i_1_737_206 (.A(\out_as[3] [4]), .B(n_1_737_5207), .CO(n_1_737_206), 
      .S());
   HA_X1 i_1_737_207 (.A(\out_as[4] [4]), .B(n_1_737_5380), .CO(n_1_737_207), 
      .S());
   HA_X1 i_1_737_208 (.A(\out_as[5] [4]), .B(n_1_737_5161), .CO(n_1_737_208), 
      .S());
   HA_X1 i_1_737_209 (.A(\out_as[6] [4]), .B(n_1_737_5149), .CO(n_1_737_209), 
      .S());
   HA_X1 i_1_737_210 (.A(\out_as[0] [4]), .B(n_1_737_1251), .CO(n_1_737_210), 
      .S());
   HA_X1 i_1_737_211 (.A(\out_as[1] [4]), .B(n_1_737_1250), .CO(n_1_737_211), 
      .S());
   HA_X1 i_1_737_212 (.A(\out_as[2] [4]), .B(n_1_737_1249), .CO(n_1_737_212), 
      .S());
   HA_X1 i_1_737_213 (.A(\out_as[3] [4]), .B(n_1_737_1248), .CO(n_1_737_213), 
      .S());
   HA_X1 i_1_737_214 (.A(\out_as[4] [4]), .B(n_1_737_1247), .CO(n_1_737_214), 
      .S());
   HA_X1 i_1_737_215 (.A(\out_as[5] [4]), .B(n_1_737_1246), .CO(n_1_737_215), 
      .S());
   HA_X1 i_1_737_216 (.A(\out_as[6] [4]), .B(n_1_737_1245), .CO(n_1_737_216), 
      .S());
   HA_X1 i_1_737_217 (.A(\out_as[0] [4]), .B(n_1_737_5351), .CO(n_1_737_217), 
      .S());
   HA_X1 i_1_737_218 (.A(\out_as[1] [4]), .B(n_1_737_5313), .CO(n_1_737_218), 
      .S());
   HA_X1 i_1_737_219 (.A(\out_as[2] [4]), .B(n_1_737_5269), .CO(n_1_737_219), 
      .S());
   HA_X1 i_1_737_220 (.A(\out_as[3] [4]), .B(n_1_737_5208), .CO(n_1_737_220), 
      .S());
   HA_X1 i_1_737_221 (.A(\out_as[4] [4]), .B(n_1_737_5381), .CO(n_1_737_221), 
      .S());
   HA_X1 i_1_737_222 (.A(\out_as[5] [4]), .B(n_1_737_5162), .CO(n_1_737_222), 
      .S());
   HA_X1 i_1_737_223 (.A(\out_as[6] [4]), .B(n_1_737_5150), .CO(n_1_737_223), 
      .S());
   HA_X1 i_1_737_224 (.A(\out_as[0] [4]), .B(n_1_737_1244), .CO(n_1_737_224), 
      .S());
   HA_X1 i_1_737_225 (.A(\out_as[1] [4]), .B(n_1_737_1243), .CO(n_1_737_225), 
      .S());
   HA_X1 i_1_737_226 (.A(\out_as[2] [4]), .B(n_1_737_1242), .CO(n_1_737_226), 
      .S());
   HA_X1 i_1_737_227 (.A(\out_as[3] [4]), .B(n_1_737_1241), .CO(n_1_737_227), 
      .S());
   HA_X1 i_1_737_228 (.A(\out_as[4] [4]), .B(n_1_737_1240), .CO(n_1_737_228), 
      .S());
   HA_X1 i_1_737_229 (.A(\out_as[5] [4]), .B(n_1_737_1239), .CO(n_1_737_229), 
      .S());
   HA_X1 i_1_737_230 (.A(\out_as[6] [4]), .B(n_1_737_1238), .CO(n_1_737_230), 
      .S());
   HA_X1 i_1_737_231 (.A(\out_as[0] [4]), .B(n_1_737_1237), .CO(n_1_737_231), 
      .S());
   HA_X1 i_1_737_232 (.A(\out_as[1] [4]), .B(n_1_737_1236), .CO(n_1_737_232), 
      .S());
   HA_X1 i_1_737_233 (.A(\out_as[2] [4]), .B(n_1_737_1235), .CO(n_1_737_233), 
      .S());
   HA_X1 i_1_737_234 (.A(\out_as[3] [4]), .B(n_1_737_1234), .CO(n_1_737_234), 
      .S());
   HA_X1 i_1_737_235 (.A(\out_as[4] [4]), .B(n_1_737_1233), .CO(n_1_737_235), 
      .S());
   HA_X1 i_1_737_236 (.A(\out_as[5] [4]), .B(n_1_737_1232), .CO(n_1_737_236), 
      .S());
   HA_X1 i_1_737_237 (.A(\out_as[6] [4]), .B(n_1_737_1231), .CO(n_1_737_237), 
      .S());
   HA_X1 i_1_737_238 (.A(\out_as[0] [4]), .B(n_1_737_1230), .CO(n_1_737_238), 
      .S());
   HA_X1 i_1_737_239 (.A(\out_as[1] [4]), .B(n_1_737_1229), .CO(n_1_737_239), 
      .S());
   HA_X1 i_1_737_240 (.A(\out_as[2] [4]), .B(n_1_737_1228), .CO(n_1_737_240), 
      .S());
   HA_X1 i_1_737_241 (.A(\out_as[3] [4]), .B(n_1_737_1227), .CO(n_1_737_241), 
      .S());
   HA_X1 i_1_737_242 (.A(\out_as[4] [4]), .B(n_1_737_1226), .CO(n_1_737_242), 
      .S());
   HA_X1 i_1_737_243 (.A(\out_as[5] [4]), .B(n_1_737_1225), .CO(n_1_737_243), 
      .S());
   HA_X1 i_1_737_244 (.A(\out_as[6] [4]), .B(n_1_737_1224), .CO(n_1_737_244), 
      .S());
   HA_X1 i_1_737_245 (.A(\out_as[0] [4]), .B(\out_as[0] [3]), .CO(n_1_737_245), 
      .S());
   HA_X1 i_1_737_246 (.A(\out_as[1] [4]), .B(\out_as[1] [3]), .CO(n_1_737_246), 
      .S());
   HA_X1 i_1_737_247 (.A(\out_as[2] [4]), .B(\out_as[2] [3]), .CO(n_1_737_247), 
      .S());
   HA_X1 i_1_737_248 (.A(\out_as[3] [4]), .B(\out_as[3] [3]), .CO(n_1_737_248), 
      .S());
   HA_X1 i_1_737_249 (.A(\out_as[4] [4]), .B(\out_as[4] [3]), .CO(n_1_737_249), 
      .S());
   HA_X1 i_1_737_250 (.A(\out_as[5] [4]), .B(\out_as[5] [3]), .CO(n_1_737_250), 
      .S());
   HA_X1 i_1_737_251 (.A(\out_as[6] [4]), .B(\out_as[6] [3]), .CO(n_1_737_251), 
      .S());
   HA_X1 i_1_737_252 (.A(\out_as[0] [4]), .B(n_1_737_147), .CO(n_1_737_252), 
      .S());
   HA_X1 i_1_737_253 (.A(\out_as[1] [4]), .B(n_1_737_148), .CO(n_1_737_253), 
      .S());
   HA_X1 i_1_737_254 (.A(\out_as[2] [4]), .B(n_1_737_149), .CO(n_1_737_254), 
      .S());
   HA_X1 i_1_737_255 (.A(\out_as[3] [4]), .B(n_1_737_150), .CO(n_1_737_255), 
      .S());
   HA_X1 i_1_737_256 (.A(\out_as[4] [4]), .B(n_1_737_151), .CO(n_1_737_256), 
      .S());
   HA_X1 i_1_737_257 (.A(\out_as[5] [4]), .B(n_1_737_152), .CO(n_1_737_257), 
      .S());
   HA_X1 i_1_737_258 (.A(\out_as[6] [4]), .B(n_1_737_153), .CO(n_1_737_258), 
      .S());
   HA_X1 i_1_737_259 (.A(\out_as[0] [4]), .B(n_1_737_154), .CO(n_1_737_259), 
      .S());
   HA_X1 i_1_737_260 (.A(\out_as[1] [4]), .B(n_1_737_155), .CO(n_1_737_260), 
      .S());
   HA_X1 i_1_737_261 (.A(\out_as[2] [4]), .B(n_1_737_156), .CO(n_1_737_261), 
      .S());
   HA_X1 i_1_737_262 (.A(\out_as[3] [4]), .B(n_1_737_157), .CO(n_1_737_262), 
      .S());
   HA_X1 i_1_737_263 (.A(\out_as[4] [4]), .B(n_1_737_158), .CO(n_1_737_263), 
      .S());
   HA_X1 i_1_737_264 (.A(\out_as[5] [4]), .B(n_1_737_159), .CO(n_1_737_264), 
      .S());
   HA_X1 i_1_737_265 (.A(\out_as[6] [4]), .B(n_1_737_160), .CO(n_1_737_265), 
      .S());
   HA_X1 i_1_737_266 (.A(\out_as[0] [4]), .B(n_1_737_161), .CO(n_1_737_266), 
      .S());
   HA_X1 i_1_737_267 (.A(\out_as[1] [4]), .B(n_1_737_162), .CO(n_1_737_267), 
      .S());
   HA_X1 i_1_737_268 (.A(\out_as[2] [4]), .B(n_1_737_163), .CO(n_1_737_268), 
      .S());
   HA_X1 i_1_737_269 (.A(\out_as[3] [4]), .B(n_1_737_164), .CO(n_1_737_269), 
      .S());
   HA_X1 i_1_737_270 (.A(\out_as[4] [4]), .B(n_1_737_165), .CO(n_1_737_270), 
      .S());
   HA_X1 i_1_737_271 (.A(\out_as[5] [4]), .B(n_1_737_166), .CO(n_1_737_271), 
      .S());
   HA_X1 i_1_737_272 (.A(\out_as[6] [4]), .B(n_1_737_167), .CO(n_1_737_272), 
      .S());
   HA_X1 i_1_737_273 (.A(\out_as[0] [4]), .B(n_1_737_168), .CO(n_1_737_273), 
      .S());
   HA_X1 i_1_737_274 (.A(\out_as[1] [4]), .B(n_1_737_169), .CO(n_1_737_274), 
      .S());
   HA_X1 i_1_737_275 (.A(\out_as[2] [4]), .B(n_1_737_170), .CO(n_1_737_275), 
      .S());
   HA_X1 i_1_737_276 (.A(\out_as[3] [4]), .B(n_1_737_171), .CO(n_1_737_276), 
      .S());
   HA_X1 i_1_737_277 (.A(\out_as[4] [4]), .B(n_1_737_172), .CO(n_1_737_277), 
      .S());
   HA_X1 i_1_737_278 (.A(\out_as[5] [4]), .B(n_1_737_173), .CO(n_1_737_278), 
      .S());
   HA_X1 i_1_737_279 (.A(\out_as[6] [4]), .B(n_1_737_174), .CO(n_1_737_279), 
      .S());
   HA_X1 i_1_737_280 (.A(\out_as[0] [4]), .B(n_1_737_175), .CO(n_1_737_280), 
      .S());
   HA_X1 i_1_737_281 (.A(\out_as[1] [4]), .B(n_1_737_176), .CO(n_1_737_281), 
      .S());
   HA_X1 i_1_737_282 (.A(\out_as[2] [4]), .B(n_1_737_177), .CO(n_1_737_282), 
      .S());
   HA_X1 i_1_737_283 (.A(\out_as[3] [4]), .B(n_1_737_178), .CO(n_1_737_283), 
      .S());
   HA_X1 i_1_737_284 (.A(\out_as[4] [4]), .B(n_1_737_179), .CO(n_1_737_284), 
      .S());
   HA_X1 i_1_737_285 (.A(\out_as[5] [4]), .B(n_1_737_180), .CO(n_1_737_285), 
      .S());
   HA_X1 i_1_737_286 (.A(\out_as[6] [4]), .B(n_1_737_181), .CO(n_1_737_286), 
      .S());
   HA_X1 i_1_737_287 (.A(\out_as[0] [4]), .B(n_1_737_182), .CO(n_1_737_287), 
      .S());
   HA_X1 i_1_737_288 (.A(\out_as[1] [4]), .B(n_1_737_183), .CO(n_1_737_288), 
      .S());
   HA_X1 i_1_737_289 (.A(\out_as[2] [4]), .B(n_1_737_184), .CO(n_1_737_289), 
      .S());
   HA_X1 i_1_737_290 (.A(\out_as[3] [4]), .B(n_1_737_185), .CO(n_1_737_290), 
      .S());
   HA_X1 i_1_737_291 (.A(\out_as[4] [4]), .B(n_1_737_186), .CO(n_1_737_291), 
      .S());
   HA_X1 i_1_737_292 (.A(\out_as[5] [4]), .B(n_1_737_187), .CO(n_1_737_292), 
      .S());
   HA_X1 i_1_737_293 (.A(\out_as[6] [4]), .B(n_1_737_188), .CO(n_1_737_293), 
      .S());
   HA_X1 i_1_737_294 (.A(\out_as[0] [4]), .B(n_1_737_189), .CO(n_1_737_294), 
      .S());
   HA_X1 i_1_737_295 (.A(\out_as[1] [4]), .B(n_1_737_190), .CO(n_1_737_295), 
      .S());
   HA_X1 i_1_737_296 (.A(\out_as[2] [4]), .B(n_1_737_191), .CO(n_1_737_296), 
      .S());
   HA_X1 i_1_737_297 (.A(\out_as[3] [4]), .B(n_1_737_192), .CO(n_1_737_297), 
      .S());
   HA_X1 i_1_737_298 (.A(\out_as[4] [4]), .B(n_1_737_193), .CO(n_1_737_298), 
      .S());
   HA_X1 i_1_737_299 (.A(\out_as[5] [4]), .B(n_1_737_194), .CO(n_1_737_299), 
      .S());
   HA_X1 i_1_737_300 (.A(\out_as[6] [4]), .B(n_1_737_195), .CO(n_1_737_300), 
      .S());
   HA_X1 i_1_737_301 (.A(\out_as[0] [5]), .B(n_1_737_2005), .CO(n_1_737_301), 
      .S());
   HA_X1 i_1_737_302 (.A(\out_as[1] [5]), .B(n_1_737_1994), .CO(n_1_737_302), 
      .S());
   HA_X1 i_1_737_303 (.A(\out_as[2] [5]), .B(n_1_737_1988), .CO(n_1_737_303), 
      .S());
   HA_X1 i_1_737_304 (.A(\out_as[3] [5]), .B(n_1_737_2016), .CO(n_1_737_304), 
      .S());
   HA_X1 i_1_737_305 (.A(\out_as[4] [5]), .B(n_1_737_1999), .CO(n_1_737_305), 
      .S());
   HA_X1 i_1_737_306 (.A(\out_as[5] [5]), .B(n_1_737_2010), .CO(n_1_737_306), 
      .S());
   HA_X1 i_1_737_307 (.A(\out_as[6] [5]), .B(n_1_737_1981), .CO(n_1_737_307), 
      .S());
   HA_X1 i_1_737_308 (.A(\out_as[0] [5]), .B(n_1_737_5348), .CO(n_1_737_308), 
      .S());
   HA_X1 i_1_737_309 (.A(\out_as[1] [5]), .B(n_1_737_5310), .CO(n_1_737_309), 
      .S());
   HA_X1 i_1_737_310 (.A(\out_as[2] [5]), .B(n_1_737_5266), .CO(n_1_737_310), 
      .S());
   HA_X1 i_1_737_311 (.A(\out_as[3] [5]), .B(n_1_737_5205), .CO(n_1_737_311), 
      .S());
   HA_X1 i_1_737_312 (.A(\out_as[4] [5]), .B(n_1_737_5378), .CO(n_1_737_312), 
      .S());
   HA_X1 i_1_737_313 (.A(\out_as[5] [5]), .B(n_1_737_5159), .CO(n_1_737_313), 
      .S());
   HA_X1 i_1_737_314 (.A(\out_as[6] [5]), .B(n_1_737_5147), .CO(n_1_737_314), 
      .S());
   HA_X1 i_1_737_315 (.A(\out_as[0] [5]), .B(n_1_737_1223), .CO(n_1_737_315), 
      .S());
   HA_X1 i_1_737_316 (.A(\out_as[1] [5]), .B(n_1_737_1222), .CO(n_1_737_316), 
      .S());
   HA_X1 i_1_737_317 (.A(\out_as[2] [5]), .B(n_1_737_1221), .CO(n_1_737_317), 
      .S());
   HA_X1 i_1_737_318 (.A(\out_as[3] [5]), .B(n_1_737_1220), .CO(n_1_737_318), 
      .S());
   HA_X1 i_1_737_319 (.A(\out_as[4] [5]), .B(n_1_737_1219), .CO(n_1_737_319), 
      .S());
   HA_X1 i_1_737_320 (.A(\out_as[5] [5]), .B(n_1_737_1218), .CO(n_1_737_320), 
      .S());
   HA_X1 i_1_737_321 (.A(\out_as[6] [5]), .B(n_1_737_1217), .CO(n_1_737_321), 
      .S());
   HA_X1 i_1_737_322 (.A(\out_as[0] [5]), .B(n_1_737_5349), .CO(n_1_737_322), 
      .S());
   HA_X1 i_1_737_323 (.A(\out_as[1] [5]), .B(n_1_737_5311), .CO(n_1_737_323), 
      .S());
   HA_X1 i_1_737_324 (.A(\out_as[2] [5]), .B(n_1_737_5267), .CO(n_1_737_324), 
      .S());
   HA_X1 i_1_737_325 (.A(\out_as[3] [5]), .B(n_1_737_5206), .CO(n_1_737_325), 
      .S());
   HA_X1 i_1_737_326 (.A(\out_as[4] [5]), .B(n_1_737_5379), .CO(n_1_737_326), 
      .S());
   HA_X1 i_1_737_327 (.A(\out_as[5] [5]), .B(n_1_737_5160), .CO(n_1_737_327), 
      .S());
   HA_X1 i_1_737_328 (.A(\out_as[6] [5]), .B(n_1_737_5148), .CO(n_1_737_328), 
      .S());
   HA_X1 i_1_737_329 (.A(\out_as[0] [5]), .B(n_1_737_1216), .CO(n_1_737_329), 
      .S());
   HA_X1 i_1_737_330 (.A(\out_as[1] [5]), .B(n_1_737_1215), .CO(n_1_737_330), 
      .S());
   HA_X1 i_1_737_331 (.A(\out_as[2] [5]), .B(n_1_737_1214), .CO(n_1_737_331), 
      .S());
   HA_X1 i_1_737_332 (.A(\out_as[3] [5]), .B(n_1_737_1213), .CO(n_1_737_332), 
      .S());
   HA_X1 i_1_737_333 (.A(\out_as[4] [5]), .B(n_1_737_1212), .CO(n_1_737_333), 
      .S());
   HA_X1 i_1_737_334 (.A(\out_as[5] [5]), .B(n_1_737_1211), .CO(n_1_737_334), 
      .S());
   HA_X1 i_1_737_335 (.A(\out_as[6] [5]), .B(n_1_737_1210), .CO(n_1_737_335), 
      .S());
   HA_X1 i_1_737_336 (.A(\out_as[0] [5]), .B(n_1_737_1209), .CO(n_1_737_336), 
      .S());
   HA_X1 i_1_737_337 (.A(\out_as[1] [5]), .B(n_1_737_1208), .CO(n_1_737_337), 
      .S());
   HA_X1 i_1_737_338 (.A(\out_as[2] [5]), .B(n_1_737_1207), .CO(n_1_737_338), 
      .S());
   HA_X1 i_1_737_339 (.A(\out_as[3] [5]), .B(n_1_737_1206), .CO(n_1_737_339), 
      .S());
   HA_X1 i_1_737_340 (.A(\out_as[4] [5]), .B(n_1_737_1205), .CO(n_1_737_340), 
      .S());
   HA_X1 i_1_737_341 (.A(\out_as[5] [5]), .B(n_1_737_1204), .CO(n_1_737_341), 
      .S());
   HA_X1 i_1_737_342 (.A(\out_as[6] [5]), .B(n_1_737_1203), .CO(n_1_737_342), 
      .S());
   HA_X1 i_1_737_343 (.A(\out_as[0] [5]), .B(n_1_737_1202), .CO(n_1_737_343), 
      .S());
   HA_X1 i_1_737_344 (.A(\out_as[1] [5]), .B(n_1_737_1201), .CO(n_1_737_344), 
      .S());
   HA_X1 i_1_737_345 (.A(\out_as[2] [5]), .B(n_1_737_1200), .CO(n_1_737_345), 
      .S());
   HA_X1 i_1_737_346 (.A(\out_as[3] [5]), .B(n_1_737_1199), .CO(n_1_737_346), 
      .S());
   HA_X1 i_1_737_347 (.A(\out_as[4] [5]), .B(n_1_737_1198), .CO(n_1_737_347), 
      .S());
   HA_X1 i_1_737_348 (.A(\out_as[5] [5]), .B(n_1_737_1197), .CO(n_1_737_348), 
      .S());
   HA_X1 i_1_737_349 (.A(\out_as[6] [5]), .B(n_1_737_1196), .CO(n_1_737_349), 
      .S());
   HA_X1 i_1_737_350 (.A(\out_as[0] [5]), .B(n_1_737_5355), .CO(n_1_737_350), 
      .S());
   HA_X1 i_1_737_351 (.A(\out_as[1] [5]), .B(n_1_737_5317), .CO(n_1_737_351), 
      .S());
   HA_X1 i_1_737_352 (.A(\out_as[2] [5]), .B(n_1_737_5272), .CO(n_1_737_352), 
      .S());
   HA_X1 i_1_737_353 (.A(\out_as[3] [5]), .B(n_1_737_5212), .CO(n_1_737_353), 
      .S());
   HA_X1 i_1_737_354 (.A(\out_as[4] [5]), .B(n_1_737_5384), .CO(n_1_737_354), 
      .S());
   HA_X1 i_1_737_355 (.A(\out_as[5] [5]), .B(n_1_737_5165), .CO(n_1_737_355), 
      .S());
   HA_X1 i_1_737_356 (.A(\out_as[6] [5]), .B(n_1_737_5153), .CO(n_1_737_356), 
      .S());
   HA_X1 i_1_737_357 (.A(\out_as[0] [5]), .B(n_1_737_1195), .CO(n_1_737_357), 
      .S());
   HA_X1 i_1_737_358 (.A(\out_as[1] [5]), .B(n_1_737_1194), .CO(n_1_737_358), 
      .S());
   HA_X1 i_1_737_359 (.A(\out_as[2] [5]), .B(n_1_737_1193), .CO(n_1_737_359), 
      .S());
   HA_X1 i_1_737_360 (.A(\out_as[3] [5]), .B(n_1_737_1192), .CO(n_1_737_360), 
      .S());
   HA_X1 i_1_737_361 (.A(\out_as[4] [5]), .B(n_1_737_1191), .CO(n_1_737_361), 
      .S());
   HA_X1 i_1_737_362 (.A(\out_as[5] [5]), .B(n_1_737_1190), .CO(n_1_737_362), 
      .S());
   HA_X1 i_1_737_363 (.A(\out_as[6] [5]), .B(n_1_737_1189), .CO(n_1_737_363), 
      .S());
   HA_X1 i_1_737_364 (.A(\out_as[0] [5]), .B(n_1_737_1188), .CO(n_1_737_364), 
      .S());
   HA_X1 i_1_737_365 (.A(\out_as[1] [5]), .B(n_1_737_1187), .CO(n_1_737_365), 
      .S());
   HA_X1 i_1_737_366 (.A(\out_as[2] [5]), .B(n_1_737_1186), .CO(n_1_737_366), 
      .S());
   HA_X1 i_1_737_367 (.A(\out_as[3] [5]), .B(n_1_737_1185), .CO(n_1_737_367), 
      .S());
   HA_X1 i_1_737_368 (.A(\out_as[4] [5]), .B(n_1_737_1184), .CO(n_1_737_368), 
      .S());
   HA_X1 i_1_737_369 (.A(\out_as[5] [5]), .B(n_1_737_1183), .CO(n_1_737_369), 
      .S());
   HA_X1 i_1_737_370 (.A(\out_as[6] [5]), .B(n_1_737_1182), .CO(n_1_737_370), 
      .S());
   HA_X1 i_1_737_371 (.A(\out_as[0] [5]), .B(n_1_737_1181), .CO(n_1_737_371), 
      .S());
   HA_X1 i_1_737_372 (.A(\out_as[1] [5]), .B(n_1_737_1180), .CO(n_1_737_372), 
      .S());
   HA_X1 i_1_737_373 (.A(\out_as[2] [5]), .B(n_1_737_1179), .CO(n_1_737_373), 
      .S());
   HA_X1 i_1_737_374 (.A(\out_as[3] [5]), .B(n_1_737_1178), .CO(n_1_737_374), 
      .S());
   HA_X1 i_1_737_375 (.A(\out_as[4] [5]), .B(n_1_737_1177), .CO(n_1_737_375), 
      .S());
   HA_X1 i_1_737_376 (.A(\out_as[5] [5]), .B(n_1_737_1176), .CO(n_1_737_376), 
      .S());
   HA_X1 i_1_737_377 (.A(\out_as[6] [5]), .B(n_1_737_1175), .CO(n_1_737_377), 
      .S());
   HA_X1 i_1_737_378 (.A(\out_as[0] [5]), .B(n_1_737_1174), .CO(n_1_737_378), 
      .S());
   HA_X1 i_1_737_379 (.A(\out_as[1] [5]), .B(n_1_737_1173), .CO(n_1_737_379), 
      .S());
   HA_X1 i_1_737_380 (.A(\out_as[2] [5]), .B(n_1_737_1172), .CO(n_1_737_380), 
      .S());
   HA_X1 i_1_737_381 (.A(\out_as[3] [5]), .B(n_1_737_1171), .CO(n_1_737_381), 
      .S());
   HA_X1 i_1_737_382 (.A(\out_as[4] [5]), .B(n_1_737_1170), .CO(n_1_737_382), 
      .S());
   HA_X1 i_1_737_383 (.A(\out_as[5] [5]), .B(n_1_737_1169), .CO(n_1_737_383), 
      .S());
   HA_X1 i_1_737_384 (.A(\out_as[6] [5]), .B(n_1_737_1168), .CO(n_1_737_384), 
      .S());
   HA_X1 i_1_737_385 (.A(\out_as[0] [5]), .B(n_1_737_1167), .CO(n_1_737_385), 
      .S());
   HA_X1 i_1_737_386 (.A(\out_as[1] [5]), .B(n_1_737_1166), .CO(n_1_737_386), 
      .S());
   HA_X1 i_1_737_387 (.A(\out_as[2] [5]), .B(n_1_737_1165), .CO(n_1_737_387), 
      .S());
   HA_X1 i_1_737_388 (.A(\out_as[3] [5]), .B(n_1_737_1164), .CO(n_1_737_388), 
      .S());
   HA_X1 i_1_737_389 (.A(\out_as[4] [5]), .B(n_1_737_1163), .CO(n_1_737_389), 
      .S());
   HA_X1 i_1_737_390 (.A(\out_as[5] [5]), .B(n_1_737_1162), .CO(n_1_737_390), 
      .S());
   HA_X1 i_1_737_391 (.A(\out_as[6] [5]), .B(n_1_737_1161), .CO(n_1_737_391), 
      .S());
   HA_X1 i_1_737_392 (.A(\out_as[0] [5]), .B(n_1_737_1160), .CO(n_1_737_392), 
      .S());
   HA_X1 i_1_737_393 (.A(\out_as[1] [5]), .B(n_1_737_1159), .CO(n_1_737_393), 
      .S());
   HA_X1 i_1_737_394 (.A(\out_as[2] [5]), .B(n_1_737_1158), .CO(n_1_737_394), 
      .S());
   HA_X1 i_1_737_395 (.A(\out_as[3] [5]), .B(n_1_737_1157), .CO(n_1_737_395), 
      .S());
   HA_X1 i_1_737_396 (.A(\out_as[4] [5]), .B(n_1_737_1156), .CO(n_1_737_396), 
      .S());
   HA_X1 i_1_737_397 (.A(\out_as[5] [5]), .B(n_1_737_1155), .CO(n_1_737_397), 
      .S());
   HA_X1 i_1_737_398 (.A(\out_as[6] [5]), .B(n_1_737_1154), .CO(n_1_737_398), 
      .S());
   HA_X1 i_1_737_399 (.A(\out_as[0] [5]), .B(n_1_737_1153), .CO(n_1_737_399), 
      .S());
   HA_X1 i_1_737_400 (.A(\out_as[1] [5]), .B(n_1_737_1152), .CO(n_1_737_400), 
      .S());
   HA_X1 i_1_737_401 (.A(\out_as[2] [5]), .B(n_1_737_1151), .CO(n_1_737_401), 
      .S());
   HA_X1 i_1_737_402 (.A(\out_as[3] [5]), .B(n_1_737_1150), .CO(n_1_737_402), 
      .S());
   HA_X1 i_1_737_403 (.A(\out_as[4] [5]), .B(n_1_737_1149), .CO(n_1_737_403), 
      .S());
   HA_X1 i_1_737_404 (.A(\out_as[5] [5]), .B(n_1_737_1148), .CO(n_1_737_404), 
      .S());
   HA_X1 i_1_737_405 (.A(\out_as[6] [5]), .B(n_1_737_1147), .CO(n_1_737_405), 
      .S());
   HA_X1 i_1_737_406 (.A(\out_as[0] [5]), .B(\out_as[0] [4]), .CO(n_1_737_406), 
      .S());
   HA_X1 i_1_737_407 (.A(\out_as[1] [5]), .B(\out_as[1] [4]), .CO(n_1_737_407), 
      .S());
   HA_X1 i_1_737_408 (.A(\out_as[2] [5]), .B(\out_as[2] [4]), .CO(n_1_737_408), 
      .S());
   HA_X1 i_1_737_409 (.A(\out_as[3] [5]), .B(\out_as[3] [4]), .CO(n_1_737_409), 
      .S());
   HA_X1 i_1_737_410 (.A(\out_as[4] [5]), .B(\out_as[4] [4]), .CO(n_1_737_410), 
      .S());
   HA_X1 i_1_737_411 (.A(\out_as[5] [5]), .B(\out_as[5] [4]), .CO(n_1_737_411), 
      .S());
   HA_X1 i_1_737_412 (.A(\out_as[6] [5]), .B(\out_as[6] [4]), .CO(n_1_737_412), 
      .S());
   HA_X1 i_1_737_413 (.A(\out_as[0] [5]), .B(n_1_737_196), .CO(n_1_737_413), 
      .S());
   HA_X1 i_1_737_414 (.A(\out_as[1] [5]), .B(n_1_737_197), .CO(n_1_737_414), 
      .S());
   HA_X1 i_1_737_415 (.A(\out_as[2] [5]), .B(n_1_737_198), .CO(n_1_737_415), 
      .S());
   HA_X1 i_1_737_416 (.A(\out_as[3] [5]), .B(n_1_737_199), .CO(n_1_737_416), 
      .S());
   HA_X1 i_1_737_417 (.A(\out_as[4] [5]), .B(n_1_737_200), .CO(n_1_737_417), 
      .S());
   HA_X1 i_1_737_418 (.A(\out_as[5] [5]), .B(n_1_737_201), .CO(n_1_737_418), 
      .S());
   HA_X1 i_1_737_419 (.A(\out_as[6] [5]), .B(n_1_737_202), .CO(n_1_737_419), 
      .S());
   HA_X1 i_1_737_420 (.A(\out_as[0] [5]), .B(n_1_737_203), .CO(n_1_737_420), 
      .S());
   HA_X1 i_1_737_421 (.A(\out_as[1] [5]), .B(n_1_737_204), .CO(n_1_737_421), 
      .S());
   HA_X1 i_1_737_422 (.A(\out_as[2] [5]), .B(n_1_737_205), .CO(n_1_737_422), 
      .S());
   HA_X1 i_1_737_423 (.A(\out_as[3] [5]), .B(n_1_737_206), .CO(n_1_737_423), 
      .S());
   HA_X1 i_1_737_424 (.A(\out_as[4] [5]), .B(n_1_737_207), .CO(n_1_737_424), 
      .S());
   HA_X1 i_1_737_425 (.A(\out_as[5] [5]), .B(n_1_737_208), .CO(n_1_737_425), 
      .S());
   HA_X1 i_1_737_426 (.A(\out_as[6] [5]), .B(n_1_737_209), .CO(n_1_737_426), 
      .S());
   HA_X1 i_1_737_427 (.A(\out_as[0] [5]), .B(n_1_737_210), .CO(n_1_737_427), 
      .S());
   HA_X1 i_1_737_428 (.A(\out_as[1] [5]), .B(n_1_737_211), .CO(n_1_737_428), 
      .S());
   HA_X1 i_1_737_429 (.A(\out_as[2] [5]), .B(n_1_737_212), .CO(n_1_737_429), 
      .S());
   HA_X1 i_1_737_430 (.A(\out_as[3] [5]), .B(n_1_737_213), .CO(n_1_737_430), 
      .S());
   HA_X1 i_1_737_431 (.A(\out_as[4] [5]), .B(n_1_737_214), .CO(n_1_737_431), 
      .S());
   HA_X1 i_1_737_432 (.A(\out_as[5] [5]), .B(n_1_737_215), .CO(n_1_737_432), 
      .S());
   HA_X1 i_1_737_433 (.A(\out_as[6] [5]), .B(n_1_737_216), .CO(n_1_737_433), 
      .S());
   HA_X1 i_1_737_434 (.A(\out_as[0] [5]), .B(n_1_737_217), .CO(n_1_737_434), 
      .S());
   HA_X1 i_1_737_435 (.A(\out_as[1] [5]), .B(n_1_737_218), .CO(n_1_737_435), 
      .S());
   HA_X1 i_1_737_436 (.A(\out_as[2] [5]), .B(n_1_737_219), .CO(n_1_737_436), 
      .S());
   HA_X1 i_1_737_437 (.A(\out_as[3] [5]), .B(n_1_737_220), .CO(n_1_737_437), 
      .S());
   HA_X1 i_1_737_438 (.A(\out_as[4] [5]), .B(n_1_737_221), .CO(n_1_737_438), 
      .S());
   HA_X1 i_1_737_439 (.A(\out_as[5] [5]), .B(n_1_737_222), .CO(n_1_737_439), 
      .S());
   HA_X1 i_1_737_440 (.A(\out_as[6] [5]), .B(n_1_737_223), .CO(n_1_737_440), 
      .S());
   HA_X1 i_1_737_441 (.A(\out_as[0] [5]), .B(n_1_737_224), .CO(n_1_737_441), 
      .S());
   HA_X1 i_1_737_442 (.A(\out_as[1] [5]), .B(n_1_737_225), .CO(n_1_737_442), 
      .S());
   HA_X1 i_1_737_443 (.A(\out_as[2] [5]), .B(n_1_737_226), .CO(n_1_737_443), 
      .S());
   HA_X1 i_1_737_444 (.A(\out_as[3] [5]), .B(n_1_737_227), .CO(n_1_737_444), 
      .S());
   HA_X1 i_1_737_445 (.A(\out_as[4] [5]), .B(n_1_737_228), .CO(n_1_737_445), 
      .S());
   HA_X1 i_1_737_446 (.A(\out_as[5] [5]), .B(n_1_737_229), .CO(n_1_737_446), 
      .S());
   HA_X1 i_1_737_447 (.A(\out_as[6] [5]), .B(n_1_737_230), .CO(n_1_737_447), 
      .S());
   HA_X1 i_1_737_448 (.A(\out_as[0] [5]), .B(n_1_737_231), .CO(n_1_737_448), 
      .S());
   HA_X1 i_1_737_449 (.A(\out_as[1] [5]), .B(n_1_737_232), .CO(n_1_737_449), 
      .S());
   HA_X1 i_1_737_450 (.A(\out_as[2] [5]), .B(n_1_737_233), .CO(n_1_737_450), 
      .S());
   HA_X1 i_1_737_451 (.A(\out_as[3] [5]), .B(n_1_737_234), .CO(n_1_737_451), 
      .S());
   HA_X1 i_1_737_452 (.A(\out_as[4] [5]), .B(n_1_737_235), .CO(n_1_737_452), 
      .S());
   HA_X1 i_1_737_453 (.A(\out_as[5] [5]), .B(n_1_737_236), .CO(n_1_737_453), 
      .S());
   HA_X1 i_1_737_454 (.A(\out_as[6] [5]), .B(n_1_737_237), .CO(n_1_737_454), 
      .S());
   HA_X1 i_1_737_455 (.A(\out_as[0] [5]), .B(n_1_737_238), .CO(n_1_737_455), 
      .S());
   HA_X1 i_1_737_456 (.A(\out_as[1] [5]), .B(n_1_737_239), .CO(n_1_737_456), 
      .S());
   HA_X1 i_1_737_457 (.A(\out_as[2] [5]), .B(n_1_737_240), .CO(n_1_737_457), 
      .S());
   HA_X1 i_1_737_458 (.A(\out_as[3] [5]), .B(n_1_737_241), .CO(n_1_737_458), 
      .S());
   HA_X1 i_1_737_459 (.A(\out_as[4] [5]), .B(n_1_737_242), .CO(n_1_737_459), 
      .S());
   HA_X1 i_1_737_460 (.A(\out_as[5] [5]), .B(n_1_737_243), .CO(n_1_737_460), 
      .S());
   HA_X1 i_1_737_461 (.A(\out_as[6] [5]), .B(n_1_737_244), .CO(n_1_737_461), 
      .S());
   HA_X1 i_1_737_462 (.A(\out_as[0] [5]), .B(n_1_737_245), .CO(n_1_737_462), 
      .S());
   HA_X1 i_1_737_463 (.A(\out_as[1] [5]), .B(n_1_737_246), .CO(n_1_737_463), 
      .S());
   HA_X1 i_1_737_464 (.A(\out_as[2] [5]), .B(n_1_737_247), .CO(n_1_737_464), 
      .S());
   HA_X1 i_1_737_465 (.A(\out_as[3] [5]), .B(n_1_737_248), .CO(n_1_737_465), 
      .S());
   HA_X1 i_1_737_466 (.A(\out_as[4] [5]), .B(n_1_737_249), .CO(n_1_737_466), 
      .S());
   HA_X1 i_1_737_467 (.A(\out_as[5] [5]), .B(n_1_737_250), .CO(n_1_737_467), 
      .S());
   HA_X1 i_1_737_468 (.A(\out_as[6] [5]), .B(n_1_737_251), .CO(n_1_737_468), 
      .S());
   HA_X1 i_1_737_469 (.A(\out_as[0] [5]), .B(n_1_737_252), .CO(n_1_737_469), 
      .S());
   HA_X1 i_1_737_470 (.A(\out_as[1] [5]), .B(n_1_737_253), .CO(n_1_737_470), 
      .S());
   HA_X1 i_1_737_471 (.A(\out_as[2] [5]), .B(n_1_737_254), .CO(n_1_737_471), 
      .S());
   HA_X1 i_1_737_472 (.A(\out_as[3] [5]), .B(n_1_737_255), .CO(n_1_737_472), 
      .S());
   HA_X1 i_1_737_473 (.A(\out_as[4] [5]), .B(n_1_737_256), .CO(n_1_737_473), 
      .S());
   HA_X1 i_1_737_474 (.A(\out_as[5] [5]), .B(n_1_737_257), .CO(n_1_737_474), 
      .S());
   HA_X1 i_1_737_475 (.A(\out_as[6] [5]), .B(n_1_737_258), .CO(n_1_737_475), 
      .S());
   HA_X1 i_1_737_476 (.A(\out_as[0] [5]), .B(n_1_737_259), .CO(n_1_737_476), 
      .S());
   HA_X1 i_1_737_477 (.A(\out_as[1] [5]), .B(n_1_737_260), .CO(n_1_737_477), 
      .S());
   HA_X1 i_1_737_478 (.A(\out_as[2] [5]), .B(n_1_737_261), .CO(n_1_737_478), 
      .S());
   HA_X1 i_1_737_479 (.A(\out_as[3] [5]), .B(n_1_737_262), .CO(n_1_737_479), 
      .S());
   HA_X1 i_1_737_480 (.A(\out_as[4] [5]), .B(n_1_737_263), .CO(n_1_737_480), 
      .S());
   HA_X1 i_1_737_481 (.A(\out_as[5] [5]), .B(n_1_737_264), .CO(n_1_737_481), 
      .S());
   HA_X1 i_1_737_482 (.A(\out_as[6] [5]), .B(n_1_737_265), .CO(n_1_737_482), 
      .S());
   HA_X1 i_1_737_483 (.A(\out_as[0] [5]), .B(n_1_737_266), .CO(n_1_737_483), 
      .S());
   HA_X1 i_1_737_484 (.A(\out_as[1] [5]), .B(n_1_737_267), .CO(n_1_737_484), 
      .S());
   HA_X1 i_1_737_485 (.A(\out_as[2] [5]), .B(n_1_737_268), .CO(n_1_737_485), 
      .S());
   HA_X1 i_1_737_486 (.A(\out_as[3] [5]), .B(n_1_737_269), .CO(n_1_737_486), 
      .S());
   HA_X1 i_1_737_487 (.A(\out_as[4] [5]), .B(n_1_737_270), .CO(n_1_737_487), 
      .S());
   HA_X1 i_1_737_488 (.A(\out_as[5] [5]), .B(n_1_737_271), .CO(n_1_737_488), 
      .S());
   HA_X1 i_1_737_489 (.A(\out_as[6] [5]), .B(n_1_737_272), .CO(n_1_737_489), 
      .S());
   HA_X1 i_1_737_490 (.A(\out_as[0] [5]), .B(n_1_737_273), .CO(n_1_737_490), 
      .S());
   HA_X1 i_1_737_491 (.A(\out_as[1] [5]), .B(n_1_737_274), .CO(n_1_737_491), 
      .S());
   HA_X1 i_1_737_492 (.A(\out_as[2] [5]), .B(n_1_737_275), .CO(n_1_737_492), 
      .S());
   HA_X1 i_1_737_493 (.A(\out_as[3] [5]), .B(n_1_737_276), .CO(n_1_737_493), 
      .S());
   HA_X1 i_1_737_494 (.A(\out_as[4] [5]), .B(n_1_737_277), .CO(n_1_737_494), 
      .S());
   HA_X1 i_1_737_495 (.A(\out_as[5] [5]), .B(n_1_737_278), .CO(n_1_737_495), 
      .S());
   HA_X1 i_1_737_496 (.A(\out_as[6] [5]), .B(n_1_737_279), .CO(n_1_737_496), 
      .S());
   HA_X1 i_1_737_497 (.A(\out_as[0] [5]), .B(n_1_737_280), .CO(n_1_737_497), 
      .S());
   HA_X1 i_1_737_498 (.A(\out_as[1] [5]), .B(n_1_737_281), .CO(n_1_737_498), 
      .S());
   HA_X1 i_1_737_499 (.A(\out_as[2] [5]), .B(n_1_737_282), .CO(n_1_737_499), 
      .S());
   HA_X1 i_1_737_500 (.A(\out_as[3] [5]), .B(n_1_737_283), .CO(n_1_737_500), 
      .S());
   HA_X1 i_1_737_501 (.A(\out_as[4] [5]), .B(n_1_737_284), .CO(n_1_737_501), 
      .S());
   HA_X1 i_1_737_502 (.A(\out_as[5] [5]), .B(n_1_737_285), .CO(n_1_737_502), 
      .S());
   HA_X1 i_1_737_503 (.A(\out_as[6] [5]), .B(n_1_737_286), .CO(n_1_737_503), 
      .S());
   HA_X1 i_1_737_504 (.A(\out_as[0] [5]), .B(n_1_737_287), .CO(n_1_737_504), 
      .S());
   HA_X1 i_1_737_505 (.A(\out_as[1] [5]), .B(n_1_737_288), .CO(n_1_737_505), 
      .S());
   HA_X1 i_1_737_506 (.A(\out_as[2] [5]), .B(n_1_737_289), .CO(n_1_737_506), 
      .S());
   HA_X1 i_1_737_507 (.A(\out_as[3] [5]), .B(n_1_737_290), .CO(n_1_737_507), 
      .S());
   HA_X1 i_1_737_508 (.A(\out_as[4] [5]), .B(n_1_737_291), .CO(n_1_737_508), 
      .S());
   HA_X1 i_1_737_509 (.A(\out_as[5] [5]), .B(n_1_737_292), .CO(n_1_737_509), 
      .S());
   HA_X1 i_1_737_510 (.A(\out_as[6] [5]), .B(n_1_737_293), .CO(n_1_737_510), 
      .S());
   HA_X1 i_1_737_511 (.A(\out_as[0] [5]), .B(n_1_737_294), .CO(n_1_737_511), 
      .S());
   HA_X1 i_1_737_512 (.A(\out_as[1] [5]), .B(n_1_737_295), .CO(n_1_737_512), 
      .S());
   HA_X1 i_1_737_513 (.A(\out_as[2] [5]), .B(n_1_737_296), .CO(n_1_737_513), 
      .S());
   HA_X1 i_1_737_514 (.A(\out_as[3] [5]), .B(n_1_737_297), .CO(n_1_737_514), 
      .S());
   HA_X1 i_1_737_515 (.A(\out_as[4] [5]), .B(n_1_737_298), .CO(n_1_737_515), 
      .S());
   HA_X1 i_1_737_516 (.A(\out_as[5] [5]), .B(n_1_737_299), .CO(n_1_737_516), 
      .S());
   HA_X1 i_1_737_517 (.A(\out_as[6] [5]), .B(n_1_737_300), .CO(n_1_737_517), 
      .S());
   HA_X1 i_1_737_518 (.A(\out_as[0] [6]), .B(n_1_737_1146), .CO(n_1_737_518), 
      .S());
   HA_X1 i_1_737_519 (.A(\out_as[1] [6]), .B(n_1_737_1145), .CO(n_1_737_519), 
      .S());
   HA_X1 i_1_737_520 (.A(\out_as[2] [6]), .B(n_1_737_1144), .CO(n_1_737_520), 
      .S());
   HA_X1 i_1_737_521 (.A(\out_as[3] [6]), .B(n_1_737_1143), .CO(n_1_737_521), 
      .S());
   HA_X1 i_1_737_522 (.A(\out_as[4] [6]), .B(n_1_737_1142), .CO(n_1_737_522), 
      .S());
   HA_X1 i_1_737_523 (.A(\out_as[5] [6]), .B(n_1_737_1141), .CO(n_1_737_523), 
      .S());
   HA_X1 i_1_737_524 (.A(\out_as[6] [6]), .B(n_1_737_1980), .CO(n_1_737_524), 
      .S());
   HA_X1 i_1_737_525 (.A(\out_as[0] [6]), .B(n_1_737_5347), .CO(n_1_737_525), 
      .S());
   HA_X1 i_1_737_526 (.A(\out_as[1] [6]), .B(n_1_737_5309), .CO(n_1_737_526), 
      .S());
   HA_X1 i_1_737_527 (.A(\out_as[2] [6]), .B(n_1_737_5265), .CO(n_1_737_527), 
      .S());
   HA_X1 i_1_737_528 (.A(\out_as[3] [6]), .B(n_1_737_5204), .CO(n_1_737_528), 
      .S());
   HA_X1 i_1_737_529 (.A(\out_as[4] [6]), .B(n_1_737_5377), .CO(n_1_737_529), 
      .S());
   HA_X1 i_1_737_530 (.A(\out_as[5] [6]), .B(n_1_737_5158), .CO(n_1_737_530), 
      .S());
   HA_X1 i_1_737_531 (.A(\out_as[6] [6]), .B(n_1_737_5146), .CO(n_1_737_531), 
      .S());
   HA_X1 i_1_737_532 (.A(\out_as[0] [6]), .B(n_1_737_1140), .CO(n_1_737_532), 
      .S());
   HA_X1 i_1_737_533 (.A(\out_as[1] [6]), .B(n_1_737_1139), .CO(n_1_737_533), 
      .S());
   HA_X1 i_1_737_534 (.A(\out_as[2] [6]), .B(n_1_737_1138), .CO(n_1_737_534), 
      .S());
   HA_X1 i_1_737_535 (.A(\out_as[3] [6]), .B(n_1_737_1137), .CO(n_1_737_535), 
      .S());
   HA_X1 i_1_737_536 (.A(\out_as[4] [6]), .B(n_1_737_1136), .CO(n_1_737_536), 
      .S());
   HA_X1 i_1_737_537 (.A(\out_as[5] [6]), .B(n_1_737_1135), .CO(n_1_737_537), 
      .S());
   HA_X1 i_1_737_538 (.A(\out_as[6] [6]), .B(n_1_737_1134), .CO(n_1_737_538), 
      .S());
   HA_X1 i_1_737_539 (.A(\out_as[0] [6]), .B(n_1_737_5088), .CO(n_1_737_539), 
      .S());
   HA_X1 i_1_737_540 (.A(\out_as[1] [6]), .B(n_1_737_5108), .CO(n_1_737_540), 
      .S());
   HA_X1 i_1_737_541 (.A(\out_as[2] [6]), .B(n_1_737_5101), .CO(n_1_737_541), 
      .S());
   HA_X1 i_1_737_542 (.A(\out_as[3] [6]), .B(n_1_737_5118), .CO(n_1_737_542), 
      .S());
   HA_X1 i_1_737_543 (.A(\out_as[4] [6]), .B(n_1_737_5136), .CO(n_1_737_543), 
      .S());
   HA_X1 i_1_737_544 (.A(\out_as[5] [6]), .B(n_1_737_5070), .CO(n_1_737_544), 
      .S());
   HA_X1 i_1_737_545 (.A(\out_as[6] [6]), .B(n_1_737_5067), .CO(n_1_737_545), 
      .S());
   HA_X1 i_1_737_546 (.A(\out_as[0] [6]), .B(n_1_737_1133), .CO(n_1_737_546), 
      .S());
   HA_X1 i_1_737_547 (.A(\out_as[1] [6]), .B(n_1_737_1132), .CO(n_1_737_547), 
      .S());
   HA_X1 i_1_737_548 (.A(\out_as[2] [6]), .B(n_1_737_1131), .CO(n_1_737_548), 
      .S());
   HA_X1 i_1_737_549 (.A(\out_as[3] [6]), .B(n_1_737_1130), .CO(n_1_737_549), 
      .S());
   HA_X1 i_1_737_550 (.A(\out_as[4] [6]), .B(n_1_737_1129), .CO(n_1_737_550), 
      .S());
   HA_X1 i_1_737_551 (.A(\out_as[5] [6]), .B(n_1_737_1128), .CO(n_1_737_551), 
      .S());
   HA_X1 i_1_737_552 (.A(\out_as[6] [6]), .B(n_1_737_1127), .CO(n_1_737_552), 
      .S());
   HA_X1 i_1_737_553 (.A(\out_as[0] [6]), .B(n_1_737_1126), .CO(n_1_737_553), 
      .S());
   HA_X1 i_1_737_554 (.A(\out_as[1] [6]), .B(n_1_737_1125), .CO(n_1_737_554), 
      .S());
   HA_X1 i_1_737_555 (.A(\out_as[2] [6]), .B(n_1_737_1124), .CO(n_1_737_555), 
      .S());
   HA_X1 i_1_737_556 (.A(\out_as[3] [6]), .B(n_1_737_1123), .CO(n_1_737_556), 
      .S());
   HA_X1 i_1_737_557 (.A(\out_as[4] [6]), .B(n_1_737_1122), .CO(n_1_737_557), 
      .S());
   HA_X1 i_1_737_558 (.A(\out_as[5] [6]), .B(n_1_737_1121), .CO(n_1_737_558), 
      .S());
   HA_X1 i_1_737_559 (.A(\out_as[6] [6]), .B(n_1_737_1120), .CO(n_1_737_559), 
      .S());
   HA_X1 i_1_737_560 (.A(\out_as[0] [6]), .B(n_1_737_1119), .CO(n_1_737_560), 
      .S());
   HA_X1 i_1_737_561 (.A(\out_as[1] [6]), .B(n_1_737_1118), .CO(n_1_737_561), 
      .S());
   HA_X1 i_1_737_562 (.A(\out_as[2] [6]), .B(n_1_737_1117), .CO(n_1_737_562), 
      .S());
   HA_X1 i_1_737_563 (.A(\out_as[3] [6]), .B(n_1_737_1116), .CO(n_1_737_563), 
      .S());
   HA_X1 i_1_737_564 (.A(\out_as[4] [6]), .B(n_1_737_1115), .CO(n_1_737_564), 
      .S());
   HA_X1 i_1_737_565 (.A(\out_as[5] [6]), .B(n_1_737_1114), .CO(n_1_737_565), 
      .S());
   HA_X1 i_1_737_566 (.A(\out_as[6] [6]), .B(n_1_737_1113), .CO(n_1_737_566), 
      .S());
   HA_X1 i_1_737_567 (.A(\out_as[0] [6]), .B(n_1_737_5354), .CO(n_1_737_567), 
      .S());
   HA_X1 i_1_737_568 (.A(\out_as[1] [6]), .B(n_1_737_5316), .CO(n_1_737_568), 
      .S());
   HA_X1 i_1_737_569 (.A(\out_as[2] [6]), .B(n_1_737_5271), .CO(n_1_737_569), 
      .S());
   HA_X1 i_1_737_570 (.A(\out_as[3] [6]), .B(n_1_737_5211), .CO(n_1_737_570), 
      .S());
   HA_X1 i_1_737_571 (.A(\out_as[4] [6]), .B(n_1_737_5383), .CO(n_1_737_571), 
      .S());
   HA_X1 i_1_737_572 (.A(\out_as[5] [6]), .B(n_1_737_5164), .CO(n_1_737_572), 
      .S());
   HA_X1 i_1_737_573 (.A(\out_as[6] [6]), .B(n_1_737_5152), .CO(n_1_737_573), 
      .S());
   HA_X1 i_1_737_574 (.A(\out_as[0] [6]), .B(n_1_737_1112), .CO(n_1_737_574), 
      .S());
   HA_X1 i_1_737_575 (.A(\out_as[1] [6]), .B(n_1_737_1111), .CO(n_1_737_575), 
      .S());
   HA_X1 i_1_737_576 (.A(\out_as[2] [6]), .B(n_1_737_1110), .CO(n_1_737_576), 
      .S());
   HA_X1 i_1_737_577 (.A(\out_as[3] [6]), .B(n_1_737_1109), .CO(n_1_737_577), 
      .S());
   HA_X1 i_1_737_578 (.A(\out_as[4] [6]), .B(n_1_737_1108), .CO(n_1_737_578), 
      .S());
   HA_X1 i_1_737_579 (.A(\out_as[5] [6]), .B(n_1_737_1107), .CO(n_1_737_579), 
      .S());
   HA_X1 i_1_737_580 (.A(\out_as[6] [6]), .B(n_1_737_1106), .CO(n_1_737_580), 
      .S());
   HA_X1 i_1_737_581 (.A(\out_as[0] [6]), .B(n_1_737_1105), .CO(n_1_737_581), 
      .S());
   HA_X1 i_1_737_582 (.A(\out_as[1] [6]), .B(n_1_737_1104), .CO(n_1_737_582), 
      .S());
   HA_X1 i_1_737_583 (.A(\out_as[2] [6]), .B(n_1_737_1103), .CO(n_1_737_583), 
      .S());
   HA_X1 i_1_737_584 (.A(\out_as[3] [6]), .B(n_1_737_1102), .CO(n_1_737_584), 
      .S());
   HA_X1 i_1_737_585 (.A(\out_as[4] [6]), .B(n_1_737_1101), .CO(n_1_737_585), 
      .S());
   HA_X1 i_1_737_586 (.A(\out_as[5] [6]), .B(n_1_737_1100), .CO(n_1_737_586), 
      .S());
   HA_X1 i_1_737_587 (.A(\out_as[6] [6]), .B(n_1_737_1099), .CO(n_1_737_587), 
      .S());
   HA_X1 i_1_737_588 (.A(\out_as[0] [6]), .B(n_1_737_1098), .CO(n_1_737_588), 
      .S());
   HA_X1 i_1_737_589 (.A(\out_as[1] [6]), .B(n_1_737_1097), .CO(n_1_737_589), 
      .S());
   HA_X1 i_1_737_590 (.A(\out_as[2] [6]), .B(n_1_737_1096), .CO(n_1_737_590), 
      .S());
   HA_X1 i_1_737_591 (.A(\out_as[3] [6]), .B(n_1_737_1095), .CO(n_1_737_591), 
      .S());
   HA_X1 i_1_737_592 (.A(\out_as[4] [6]), .B(n_1_737_1094), .CO(n_1_737_592), 
      .S());
   HA_X1 i_1_737_593 (.A(\out_as[5] [6]), .B(n_1_737_1093), .CO(n_1_737_593), 
      .S());
   HA_X1 i_1_737_594 (.A(\out_as[6] [6]), .B(n_1_737_1092), .CO(n_1_737_594), 
      .S());
   HA_X1 i_1_737_595 (.A(\out_as[0] [6]), .B(n_1_737_1091), .CO(n_1_737_595), 
      .S());
   HA_X1 i_1_737_596 (.A(\out_as[1] [6]), .B(n_1_737_1090), .CO(n_1_737_596), 
      .S());
   HA_X1 i_1_737_597 (.A(\out_as[2] [6]), .B(n_1_737_1089), .CO(n_1_737_597), 
      .S());
   HA_X1 i_1_737_598 (.A(\out_as[3] [6]), .B(n_1_737_1088), .CO(n_1_737_598), 
      .S());
   HA_X1 i_1_737_599 (.A(\out_as[4] [6]), .B(n_1_737_1087), .CO(n_1_737_599), 
      .S());
   HA_X1 i_1_737_600 (.A(\out_as[5] [6]), .B(n_1_737_1086), .CO(n_1_737_600), 
      .S());
   HA_X1 i_1_737_601 (.A(\out_as[6] [6]), .B(n_1_737_1085), .CO(n_1_737_601), 
      .S());
   HA_X1 i_1_737_602 (.A(\out_as[0] [6]), .B(n_1_737_1084), .CO(n_1_737_602), 
      .S());
   HA_X1 i_1_737_603 (.A(\out_as[1] [6]), .B(n_1_737_1083), .CO(n_1_737_603), 
      .S());
   HA_X1 i_1_737_604 (.A(\out_as[2] [6]), .B(n_1_737_1082), .CO(n_1_737_604), 
      .S());
   HA_X1 i_1_737_605 (.A(\out_as[3] [6]), .B(n_1_737_1081), .CO(n_1_737_605), 
      .S());
   HA_X1 i_1_737_606 (.A(\out_as[4] [6]), .B(n_1_737_1080), .CO(n_1_737_606), 
      .S());
   HA_X1 i_1_737_607 (.A(\out_as[5] [6]), .B(n_1_737_1079), .CO(n_1_737_607), 
      .S());
   HA_X1 i_1_737_608 (.A(\out_as[6] [6]), .B(n_1_737_1078), .CO(n_1_737_608), 
      .S());
   HA_X1 i_1_737_609 (.A(\out_as[0] [6]), .B(n_1_737_1077), .CO(n_1_737_609), 
      .S());
   HA_X1 i_1_737_610 (.A(\out_as[1] [6]), .B(n_1_737_1076), .CO(n_1_737_610), 
      .S());
   HA_X1 i_1_737_611 (.A(\out_as[2] [6]), .B(n_1_737_1075), .CO(n_1_737_611), 
      .S());
   HA_X1 i_1_737_612 (.A(\out_as[3] [6]), .B(n_1_737_1074), .CO(n_1_737_612), 
      .S());
   HA_X1 i_1_737_613 (.A(\out_as[4] [6]), .B(n_1_737_1073), .CO(n_1_737_613), 
      .S());
   HA_X1 i_1_737_614 (.A(\out_as[5] [6]), .B(n_1_737_1072), .CO(n_1_737_614), 
      .S());
   HA_X1 i_1_737_615 (.A(\out_as[6] [6]), .B(n_1_737_1071), .CO(n_1_737_615), 
      .S());
   HA_X1 i_1_737_616 (.A(\out_as[0] [6]), .B(n_1_737_1070), .CO(n_1_737_616), 
      .S());
   HA_X1 i_1_737_617 (.A(\out_as[1] [6]), .B(n_1_737_1069), .CO(n_1_737_617), 
      .S());
   HA_X1 i_1_737_618 (.A(\out_as[2] [6]), .B(n_1_737_1068), .CO(n_1_737_618), 
      .S());
   HA_X1 i_1_737_619 (.A(\out_as[3] [6]), .B(n_1_737_1067), .CO(n_1_737_619), 
      .S());
   HA_X1 i_1_737_620 (.A(\out_as[4] [6]), .B(n_1_737_1066), .CO(n_1_737_620), 
      .S());
   HA_X1 i_1_737_621 (.A(\out_as[5] [6]), .B(n_1_737_1065), .CO(n_1_737_621), 
      .S());
   HA_X1 i_1_737_622 (.A(\out_as[6] [6]), .B(n_1_737_1064), .CO(n_1_737_622), 
      .S());
   HA_X1 i_1_737_623 (.A(\out_as[0] [6]), .B(n_1_737_5360), .CO(n_1_737_623), 
      .S());
   HA_X1 i_1_737_624 (.A(\out_as[1] [6]), .B(n_1_737_5322), .CO(n_1_737_624), 
      .S());
   HA_X1 i_1_737_625 (.A(\out_as[2] [6]), .B(n_1_737_5276), .CO(n_1_737_625), 
      .S());
   HA_X1 i_1_737_626 (.A(\out_as[3] [6]), .B(n_1_737_5217), .CO(n_1_737_626), 
      .S());
   HA_X1 i_1_737_627 (.A(\out_as[4] [6]), .B(n_1_737_5388), .CO(n_1_737_627), 
      .S());
   HA_X1 i_1_737_628 (.A(\out_as[5] [6]), .B(n_1_737_5169), .CO(n_1_737_628), 
      .S());
   HA_X1 i_1_737_629 (.A(\out_as[6] [6]), .B(n_1_737_5156), .CO(n_1_737_629), 
      .S());
   HA_X1 i_1_737_630 (.A(\out_as[0] [6]), .B(n_1_737_1063), .CO(n_1_737_630), 
      .S());
   HA_X1 i_1_737_631 (.A(\out_as[1] [6]), .B(n_1_737_1062), .CO(n_1_737_631), 
      .S());
   HA_X1 i_1_737_632 (.A(\out_as[2] [6]), .B(n_1_737_1061), .CO(n_1_737_632), 
      .S());
   HA_X1 i_1_737_633 (.A(\out_as[3] [6]), .B(n_1_737_1060), .CO(n_1_737_633), 
      .S());
   HA_X1 i_1_737_634 (.A(\out_as[4] [6]), .B(n_1_737_1059), .CO(n_1_737_634), 
      .S());
   HA_X1 i_1_737_635 (.A(\out_as[5] [6]), .B(n_1_737_1058), .CO(n_1_737_635), 
      .S());
   HA_X1 i_1_737_636 (.A(\out_as[6] [6]), .B(n_1_737_1057), .CO(n_1_737_636), 
      .S());
   HA_X1 i_1_737_637 (.A(\out_as[0] [6]), .B(n_1_737_1056), .CO(n_1_737_637), 
      .S());
   HA_X1 i_1_737_638 (.A(\out_as[1] [6]), .B(n_1_737_1055), .CO(n_1_737_638), 
      .S());
   HA_X1 i_1_737_639 (.A(\out_as[2] [6]), .B(n_1_737_1054), .CO(n_1_737_639), 
      .S());
   HA_X1 i_1_737_640 (.A(\out_as[3] [6]), .B(n_1_737_1053), .CO(n_1_737_640), 
      .S());
   HA_X1 i_1_737_641 (.A(\out_as[4] [6]), .B(n_1_737_1052), .CO(n_1_737_641), 
      .S());
   HA_X1 i_1_737_642 (.A(\out_as[5] [6]), .B(n_1_737_1051), .CO(n_1_737_642), 
      .S());
   HA_X1 i_1_737_643 (.A(\out_as[6] [6]), .B(n_1_737_1050), .CO(n_1_737_643), 
      .S());
   HA_X1 i_1_737_644 (.A(\out_as[0] [6]), .B(n_1_737_1049), .CO(n_1_737_644), 
      .S());
   HA_X1 i_1_737_645 (.A(\out_as[1] [6]), .B(n_1_737_1048), .CO(n_1_737_645), 
      .S());
   HA_X1 i_1_737_646 (.A(\out_as[2] [6]), .B(n_1_737_1047), .CO(n_1_737_646), 
      .S());
   HA_X1 i_1_737_647 (.A(\out_as[3] [6]), .B(n_1_737_1046), .CO(n_1_737_647), 
      .S());
   HA_X1 i_1_737_648 (.A(\out_as[4] [6]), .B(n_1_737_1045), .CO(n_1_737_648), 
      .S());
   HA_X1 i_1_737_649 (.A(\out_as[5] [6]), .B(n_1_737_1044), .CO(n_1_737_649), 
      .S());
   HA_X1 i_1_737_650 (.A(\out_as[6] [6]), .B(n_1_737_1043), .CO(n_1_737_650), 
      .S());
   HA_X1 i_1_737_651 (.A(\out_as[0] [6]), .B(n_1_737_1042), .CO(n_1_737_651), 
      .S());
   HA_X1 i_1_737_652 (.A(\out_as[1] [6]), .B(n_1_737_1041), .CO(n_1_737_652), 
      .S());
   HA_X1 i_1_737_653 (.A(\out_as[2] [6]), .B(n_1_737_1040), .CO(n_1_737_653), 
      .S());
   HA_X1 i_1_737_654 (.A(\out_as[3] [6]), .B(n_1_737_1039), .CO(n_1_737_654), 
      .S());
   HA_X1 i_1_737_655 (.A(\out_as[4] [6]), .B(n_1_737_1038), .CO(n_1_737_655), 
      .S());
   HA_X1 i_1_737_656 (.A(\out_as[5] [6]), .B(n_1_737_1037), .CO(n_1_737_656), 
      .S());
   HA_X1 i_1_737_657 (.A(\out_as[6] [6]), .B(n_1_737_1036), .CO(n_1_737_657), 
      .S());
   HA_X1 i_1_737_658 (.A(\out_as[0] [6]), .B(n_1_737_1035), .CO(n_1_737_658), 
      .S());
   HA_X1 i_1_737_659 (.A(\out_as[1] [6]), .B(n_1_737_1034), .CO(n_1_737_659), 
      .S());
   HA_X1 i_1_737_660 (.A(\out_as[2] [6]), .B(n_1_737_1033), .CO(n_1_737_660), 
      .S());
   HA_X1 i_1_737_661 (.A(\out_as[3] [6]), .B(n_1_737_1032), .CO(n_1_737_661), 
      .S());
   HA_X1 i_1_737_662 (.A(\out_as[4] [6]), .B(n_1_737_1031), .CO(n_1_737_662), 
      .S());
   HA_X1 i_1_737_663 (.A(\out_as[5] [6]), .B(n_1_737_1030), .CO(n_1_737_663), 
      .S());
   HA_X1 i_1_737_664 (.A(\out_as[6] [6]), .B(n_1_737_1029), .CO(n_1_737_664), 
      .S());
   HA_X1 i_1_737_665 (.A(\out_as[0] [6]), .B(n_1_737_1028), .CO(n_1_737_665), 
      .S());
   HA_X1 i_1_737_666 (.A(\out_as[1] [6]), .B(n_1_737_1027), .CO(n_1_737_666), 
      .S());
   HA_X1 i_1_737_667 (.A(\out_as[2] [6]), .B(n_1_737_1026), .CO(n_1_737_667), 
      .S());
   HA_X1 i_1_737_668 (.A(\out_as[3] [6]), .B(n_1_737_1025), .CO(n_1_737_668), 
      .S());
   HA_X1 i_1_737_669 (.A(\out_as[4] [6]), .B(n_1_737_1024), .CO(n_1_737_669), 
      .S());
   HA_X1 i_1_737_670 (.A(\out_as[5] [6]), .B(n_1_737_1023), .CO(n_1_737_670), 
      .S());
   HA_X1 i_1_737_671 (.A(\out_as[6] [6]), .B(n_1_737_1022), .CO(n_1_737_671), 
      .S());
   HA_X1 i_1_737_672 (.A(\out_as[0] [6]), .B(n_1_737_1021), .CO(n_1_737_672), 
      .S());
   HA_X1 i_1_737_673 (.A(\out_as[1] [6]), .B(n_1_737_1020), .CO(n_1_737_673), 
      .S());
   HA_X1 i_1_737_674 (.A(\out_as[2] [6]), .B(n_1_737_1019), .CO(n_1_737_674), 
      .S());
   HA_X1 i_1_737_675 (.A(\out_as[3] [6]), .B(n_1_737_1018), .CO(n_1_737_675), 
      .S());
   HA_X1 i_1_737_676 (.A(\out_as[4] [6]), .B(n_1_737_1017), .CO(n_1_737_676), 
      .S());
   HA_X1 i_1_737_677 (.A(\out_as[5] [6]), .B(n_1_737_1016), .CO(n_1_737_677), 
      .S());
   HA_X1 i_1_737_678 (.A(\out_as[6] [6]), .B(n_1_737_1015), .CO(n_1_737_678), 
      .S());
   HA_X1 i_1_737_679 (.A(\out_as[0] [6]), .B(n_1_737_1014), .CO(n_1_737_679), 
      .S());
   HA_X1 i_1_737_680 (.A(\out_as[1] [6]), .B(n_1_737_1013), .CO(n_1_737_680), 
      .S());
   HA_X1 i_1_737_681 (.A(\out_as[2] [6]), .B(n_1_737_1012), .CO(n_1_737_681), 
      .S());
   HA_X1 i_1_737_682 (.A(\out_as[3] [6]), .B(n_1_737_1011), .CO(n_1_737_682), 
      .S());
   HA_X1 i_1_737_683 (.A(\out_as[4] [6]), .B(n_1_737_1010), .CO(n_1_737_683), 
      .S());
   HA_X1 i_1_737_684 (.A(\out_as[5] [6]), .B(n_1_737_1009), .CO(n_1_737_684), 
      .S());
   HA_X1 i_1_737_685 (.A(\out_as[6] [6]), .B(n_1_737_1008), .CO(n_1_737_685), 
      .S());
   HA_X1 i_1_737_686 (.A(\out_as[0] [6]), .B(n_1_737_1007), .CO(n_1_737_686), 
      .S());
   HA_X1 i_1_737_687 (.A(\out_as[1] [6]), .B(n_1_737_1006), .CO(n_1_737_687), 
      .S());
   HA_X1 i_1_737_688 (.A(\out_as[2] [6]), .B(n_1_737_1005), .CO(n_1_737_688), 
      .S());
   HA_X1 i_1_737_689 (.A(\out_as[3] [6]), .B(n_1_737_1004), .CO(n_1_737_689), 
      .S());
   HA_X1 i_1_737_690 (.A(\out_as[4] [6]), .B(n_1_737_1003), .CO(n_1_737_690), 
      .S());
   HA_X1 i_1_737_691 (.A(\out_as[5] [6]), .B(n_1_737_1002), .CO(n_1_737_691), 
      .S());
   HA_X1 i_1_737_692 (.A(\out_as[6] [6]), .B(n_1_737_1001), .CO(n_1_737_692), 
      .S());
   HA_X1 i_1_737_693 (.A(\out_as[0] [6]), .B(n_1_737_1000), .CO(n_1_737_693), 
      .S());
   HA_X1 i_1_737_694 (.A(\out_as[1] [6]), .B(n_1_737_999), .CO(n_1_737_694), 
      .S());
   HA_X1 i_1_737_695 (.A(\out_as[2] [6]), .B(n_1_737_998), .CO(n_1_737_695), 
      .S());
   HA_X1 i_1_737_696 (.A(\out_as[3] [6]), .B(n_1_737_997), .CO(n_1_737_696), 
      .S());
   HA_X1 i_1_737_697 (.A(\out_as[4] [6]), .B(n_1_737_996), .CO(n_1_737_697), 
      .S());
   HA_X1 i_1_737_698 (.A(\out_as[5] [6]), .B(n_1_737_995), .CO(n_1_737_698), 
      .S());
   HA_X1 i_1_737_699 (.A(\out_as[6] [6]), .B(n_1_737_994), .CO(n_1_737_699), 
      .S());
   HA_X1 i_1_737_700 (.A(\out_as[0] [6]), .B(n_1_737_993), .CO(n_1_737_700), 
      .S());
   HA_X1 i_1_737_701 (.A(\out_as[1] [6]), .B(n_1_737_992), .CO(n_1_737_701), 
      .S());
   HA_X1 i_1_737_702 (.A(\out_as[2] [6]), .B(n_1_737_991), .CO(n_1_737_702), 
      .S());
   HA_X1 i_1_737_703 (.A(\out_as[3] [6]), .B(n_1_737_990), .CO(n_1_737_703), 
      .S());
   HA_X1 i_1_737_704 (.A(\out_as[4] [6]), .B(n_1_737_989), .CO(n_1_737_704), 
      .S());
   HA_X1 i_1_737_705 (.A(\out_as[5] [6]), .B(n_1_737_988), .CO(n_1_737_705), 
      .S());
   HA_X1 i_1_737_706 (.A(\out_as[6] [6]), .B(n_1_737_987), .CO(n_1_737_706), 
      .S());
   HA_X1 i_1_737_707 (.A(\out_as[0] [6]), .B(n_1_737_986), .CO(n_1_737_707), 
      .S());
   HA_X1 i_1_737_708 (.A(\out_as[1] [6]), .B(n_1_737_985), .CO(n_1_737_708), 
      .S());
   HA_X1 i_1_737_709 (.A(\out_as[2] [6]), .B(n_1_737_984), .CO(n_1_737_709), 
      .S());
   HA_X1 i_1_737_710 (.A(\out_as[3] [6]), .B(n_1_737_983), .CO(n_1_737_710), 
      .S());
   HA_X1 i_1_737_711 (.A(\out_as[4] [6]), .B(n_1_737_982), .CO(n_1_737_711), 
      .S());
   HA_X1 i_1_737_712 (.A(\out_as[5] [6]), .B(n_1_737_981), .CO(n_1_737_712), 
      .S());
   HA_X1 i_1_737_713 (.A(\out_as[6] [6]), .B(n_1_737_980), .CO(n_1_737_713), 
      .S());
   HA_X1 i_1_737_714 (.A(\out_as[0] [6]), .B(n_1_737_979), .CO(n_1_737_714), 
      .S());
   HA_X1 i_1_737_715 (.A(\out_as[1] [6]), .B(n_1_737_978), .CO(n_1_737_715), 
      .S());
   HA_X1 i_1_737_716 (.A(\out_as[2] [6]), .B(n_1_737_977), .CO(n_1_737_716), 
      .S());
   HA_X1 i_1_737_717 (.A(\out_as[3] [6]), .B(n_1_737_976), .CO(n_1_737_717), 
      .S());
   HA_X1 i_1_737_718 (.A(\out_as[4] [6]), .B(n_1_737_975), .CO(n_1_737_718), 
      .S());
   HA_X1 i_1_737_719 (.A(\out_as[5] [6]), .B(n_1_737_974), .CO(n_1_737_719), 
      .S());
   HA_X1 i_1_737_720 (.A(\out_as[6] [6]), .B(n_1_737_973), .CO(n_1_737_720), 
      .S());
   HA_X1 i_1_737_721 (.A(\out_as[0] [6]), .B(n_1_737_972), .CO(n_1_737_721), 
      .S());
   HA_X1 i_1_737_722 (.A(\out_as[1] [6]), .B(n_1_737_971), .CO(n_1_737_722), 
      .S());
   HA_X1 i_1_737_723 (.A(\out_as[2] [6]), .B(n_1_737_970), .CO(n_1_737_723), 
      .S());
   HA_X1 i_1_737_724 (.A(\out_as[3] [6]), .B(n_1_737_969), .CO(n_1_737_724), 
      .S());
   HA_X1 i_1_737_725 (.A(\out_as[4] [6]), .B(n_1_737_968), .CO(n_1_737_725), 
      .S());
   HA_X1 i_1_737_726 (.A(\out_as[5] [6]), .B(n_1_737_967), .CO(n_1_737_726), 
      .S());
   HA_X1 i_1_737_727 (.A(\out_as[6] [6]), .B(n_1_737_966), .CO(n_1_737_727), 
      .S());
   HA_X1 i_1_737_728 (.A(\out_as[0] [6]), .B(n_1_737_965), .CO(n_1_737_728), 
      .S());
   HA_X1 i_1_737_729 (.A(\out_as[1] [6]), .B(n_1_737_964), .CO(n_1_737_729), 
      .S());
   HA_X1 i_1_737_730 (.A(\out_as[2] [6]), .B(n_1_737_963), .CO(n_1_737_730), 
      .S());
   HA_X1 i_1_737_731 (.A(\out_as[3] [6]), .B(n_1_737_962), .CO(n_1_737_731), 
      .S());
   HA_X1 i_1_737_732 (.A(\out_as[4] [6]), .B(n_1_737_961), .CO(n_1_737_732), 
      .S());
   HA_X1 i_1_737_733 (.A(\out_as[5] [6]), .B(n_1_737_960), .CO(n_1_737_733), 
      .S());
   HA_X1 i_1_737_734 (.A(\out_as[6] [6]), .B(n_1_737_959), .CO(n_1_737_734), 
      .S());
   HA_X1 i_1_737_735 (.A(\out_as[0] [6]), .B(\out_as[0] [5]), .CO(n_1_737_735), 
      .S());
   HA_X1 i_1_737_736 (.A(\out_as[1] [6]), .B(\out_as[1] [5]), .CO(n_1_737_736), 
      .S());
   HA_X1 i_1_737_737 (.A(\out_as[2] [6]), .B(\out_as[2] [5]), .CO(n_1_737_737), 
      .S());
   HA_X1 i_1_737_738 (.A(\out_as[3] [6]), .B(\out_as[3] [5]), .CO(n_1_737_738), 
      .S());
   HA_X1 i_1_737_739 (.A(\out_as[4] [6]), .B(\out_as[4] [5]), .CO(n_1_737_739), 
      .S());
   HA_X1 i_1_737_740 (.A(\out_as[5] [6]), .B(\out_as[5] [5]), .CO(n_1_737_740), 
      .S());
   HA_X1 i_1_737_741 (.A(\out_as[6] [6]), .B(\out_as[6] [5]), .CO(n_1_737_741), 
      .S());
   HA_X1 i_1_737_742 (.A(\out_as[0] [6]), .B(n_1_737_301), .CO(n_1_737_742), 
      .S());
   HA_X1 i_1_737_743 (.A(\out_as[1] [6]), .B(n_1_737_302), .CO(n_1_737_743), 
      .S());
   HA_X1 i_1_737_744 (.A(\out_as[2] [6]), .B(n_1_737_303), .CO(n_1_737_744), 
      .S());
   HA_X1 i_1_737_745 (.A(\out_as[3] [6]), .B(n_1_737_304), .CO(n_1_737_745), 
      .S());
   HA_X1 i_1_737_746 (.A(\out_as[4] [6]), .B(n_1_737_305), .CO(n_1_737_746), 
      .S());
   HA_X1 i_1_737_747 (.A(\out_as[5] [6]), .B(n_1_737_306), .CO(n_1_737_747), 
      .S());
   HA_X1 i_1_737_748 (.A(\out_as[6] [6]), .B(n_1_737_307), .CO(n_1_737_748), 
      .S());
   HA_X1 i_1_737_749 (.A(\out_as[0] [6]), .B(n_1_737_308), .CO(n_1_737_749), 
      .S());
   HA_X1 i_1_737_750 (.A(\out_as[1] [6]), .B(n_1_737_309), .CO(n_1_737_750), 
      .S());
   HA_X1 i_1_737_751 (.A(\out_as[2] [6]), .B(n_1_737_310), .CO(n_1_737_751), 
      .S());
   HA_X1 i_1_737_752 (.A(\out_as[3] [6]), .B(n_1_737_311), .CO(n_1_737_752), 
      .S());
   HA_X1 i_1_737_753 (.A(\out_as[4] [6]), .B(n_1_737_312), .CO(n_1_737_753), 
      .S());
   HA_X1 i_1_737_754 (.A(\out_as[5] [6]), .B(n_1_737_313), .CO(n_1_737_754), 
      .S());
   HA_X1 i_1_737_755 (.A(\out_as[6] [6]), .B(n_1_737_314), .CO(n_1_737_755), 
      .S());
   HA_X1 i_1_737_756 (.A(\out_as[0] [6]), .B(n_1_737_315), .CO(n_1_737_756), 
      .S());
   HA_X1 i_1_737_757 (.A(\out_as[1] [6]), .B(n_1_737_316), .CO(n_1_737_757), 
      .S());
   HA_X1 i_1_737_758 (.A(\out_as[2] [6]), .B(n_1_737_317), .CO(n_1_737_758), 
      .S());
   HA_X1 i_1_737_759 (.A(\out_as[3] [6]), .B(n_1_737_318), .CO(n_1_737_759), 
      .S());
   HA_X1 i_1_737_760 (.A(\out_as[4] [6]), .B(n_1_737_319), .CO(n_1_737_760), 
      .S());
   HA_X1 i_1_737_761 (.A(\out_as[5] [6]), .B(n_1_737_320), .CO(n_1_737_761), 
      .S());
   HA_X1 i_1_737_762 (.A(\out_as[6] [6]), .B(n_1_737_321), .CO(n_1_737_762), 
      .S());
   HA_X1 i_1_737_763 (.A(\out_as[0] [6]), .B(n_1_737_322), .CO(n_1_737_763), 
      .S());
   HA_X1 i_1_737_764 (.A(\out_as[1] [6]), .B(n_1_737_323), .CO(n_1_737_764), 
      .S());
   HA_X1 i_1_737_765 (.A(\out_as[2] [6]), .B(n_1_737_324), .CO(n_1_737_765), 
      .S());
   HA_X1 i_1_737_766 (.A(\out_as[3] [6]), .B(n_1_737_325), .CO(n_1_737_766), 
      .S());
   HA_X1 i_1_737_767 (.A(\out_as[4] [6]), .B(n_1_737_326), .CO(n_1_737_767), 
      .S());
   HA_X1 i_1_737_768 (.A(\out_as[5] [6]), .B(n_1_737_327), .CO(n_1_737_768), 
      .S());
   HA_X1 i_1_737_769 (.A(\out_as[6] [6]), .B(n_1_737_328), .CO(n_1_737_769), 
      .S());
   HA_X1 i_1_737_770 (.A(\out_as[0] [6]), .B(n_1_737_329), .CO(n_1_737_770), 
      .S());
   HA_X1 i_1_737_771 (.A(\out_as[1] [6]), .B(n_1_737_330), .CO(n_1_737_771), 
      .S());
   HA_X1 i_1_737_772 (.A(\out_as[2] [6]), .B(n_1_737_331), .CO(n_1_737_772), 
      .S());
   HA_X1 i_1_737_773 (.A(\out_as[3] [6]), .B(n_1_737_332), .CO(n_1_737_773), 
      .S());
   HA_X1 i_1_737_774 (.A(\out_as[4] [6]), .B(n_1_737_333), .CO(n_1_737_774), 
      .S());
   HA_X1 i_1_737_775 (.A(\out_as[5] [6]), .B(n_1_737_334), .CO(n_1_737_775), 
      .S());
   HA_X1 i_1_737_776 (.A(\out_as[6] [6]), .B(n_1_737_335), .CO(n_1_737_776), 
      .S());
   HA_X1 i_1_737_777 (.A(\out_as[0] [6]), .B(n_1_737_336), .CO(n_1_737_777), 
      .S());
   HA_X1 i_1_737_778 (.A(\out_as[1] [6]), .B(n_1_737_337), .CO(n_1_737_778), 
      .S());
   HA_X1 i_1_737_779 (.A(\out_as[2] [6]), .B(n_1_737_338), .CO(n_1_737_779), 
      .S());
   HA_X1 i_1_737_780 (.A(\out_as[3] [6]), .B(n_1_737_339), .CO(n_1_737_780), 
      .S());
   HA_X1 i_1_737_781 (.A(\out_as[4] [6]), .B(n_1_737_340), .CO(n_1_737_781), 
      .S());
   HA_X1 i_1_737_782 (.A(\out_as[5] [6]), .B(n_1_737_341), .CO(n_1_737_782), 
      .S());
   HA_X1 i_1_737_783 (.A(\out_as[6] [6]), .B(n_1_737_342), .CO(n_1_737_783), 
      .S());
   HA_X1 i_1_737_784 (.A(\out_as[0] [6]), .B(n_1_737_343), .CO(n_1_737_784), 
      .S());
   HA_X1 i_1_737_785 (.A(\out_as[1] [6]), .B(n_1_737_344), .CO(n_1_737_785), 
      .S());
   HA_X1 i_1_737_786 (.A(\out_as[2] [6]), .B(n_1_737_345), .CO(n_1_737_786), 
      .S());
   HA_X1 i_1_737_787 (.A(\out_as[3] [6]), .B(n_1_737_346), .CO(n_1_737_787), 
      .S());
   HA_X1 i_1_737_788 (.A(\out_as[4] [6]), .B(n_1_737_347), .CO(n_1_737_788), 
      .S());
   HA_X1 i_1_737_789 (.A(\out_as[5] [6]), .B(n_1_737_348), .CO(n_1_737_789), 
      .S());
   HA_X1 i_1_737_790 (.A(\out_as[6] [6]), .B(n_1_737_349), .CO(n_1_737_790), 
      .S());
   HA_X1 i_1_737_791 (.A(\out_as[0] [6]), .B(n_1_737_350), .CO(n_1_737_791), 
      .S());
   HA_X1 i_1_737_792 (.A(\out_as[1] [6]), .B(n_1_737_351), .CO(n_1_737_792), 
      .S());
   HA_X1 i_1_737_793 (.A(\out_as[2] [6]), .B(n_1_737_352), .CO(n_1_737_793), 
      .S());
   HA_X1 i_1_737_794 (.A(\out_as[3] [6]), .B(n_1_737_353), .CO(n_1_737_794), 
      .S());
   HA_X1 i_1_737_795 (.A(\out_as[4] [6]), .B(n_1_737_354), .CO(n_1_737_795), 
      .S());
   HA_X1 i_1_737_796 (.A(\out_as[5] [6]), .B(n_1_737_355), .CO(n_1_737_796), 
      .S());
   HA_X1 i_1_737_797 (.A(\out_as[6] [6]), .B(n_1_737_356), .CO(n_1_737_797), 
      .S());
   HA_X1 i_1_737_798 (.A(\out_as[0] [6]), .B(n_1_737_357), .CO(n_1_737_798), 
      .S());
   HA_X1 i_1_737_799 (.A(\out_as[1] [6]), .B(n_1_737_358), .CO(n_1_737_799), 
      .S());
   HA_X1 i_1_737_800 (.A(\out_as[2] [6]), .B(n_1_737_359), .CO(n_1_737_800), 
      .S());
   HA_X1 i_1_737_801 (.A(\out_as[3] [6]), .B(n_1_737_360), .CO(n_1_737_801), 
      .S());
   HA_X1 i_1_737_802 (.A(\out_as[4] [6]), .B(n_1_737_361), .CO(n_1_737_802), 
      .S());
   HA_X1 i_1_737_803 (.A(\out_as[5] [6]), .B(n_1_737_362), .CO(n_1_737_803), 
      .S());
   HA_X1 i_1_737_804 (.A(\out_as[6] [6]), .B(n_1_737_363), .CO(n_1_737_804), 
      .S());
   HA_X1 i_1_737_805 (.A(\out_as[0] [6]), .B(n_1_737_364), .CO(n_1_737_805), 
      .S());
   HA_X1 i_1_737_806 (.A(\out_as[1] [6]), .B(n_1_737_365), .CO(n_1_737_806), 
      .S());
   HA_X1 i_1_737_807 (.A(\out_as[2] [6]), .B(n_1_737_366), .CO(n_1_737_807), 
      .S());
   HA_X1 i_1_737_808 (.A(\out_as[3] [6]), .B(n_1_737_367), .CO(n_1_737_808), 
      .S());
   HA_X1 i_1_737_809 (.A(\out_as[4] [6]), .B(n_1_737_368), .CO(n_1_737_809), 
      .S());
   HA_X1 i_1_737_810 (.A(\out_as[5] [6]), .B(n_1_737_369), .CO(n_1_737_810), 
      .S());
   HA_X1 i_1_737_811 (.A(\out_as[6] [6]), .B(n_1_737_370), .CO(n_1_737_811), 
      .S());
   HA_X1 i_1_737_812 (.A(\out_as[0] [6]), .B(n_1_737_371), .CO(n_1_737_812), 
      .S());
   HA_X1 i_1_737_813 (.A(\out_as[1] [6]), .B(n_1_737_372), .CO(n_1_737_813), 
      .S());
   HA_X1 i_1_737_814 (.A(\out_as[2] [6]), .B(n_1_737_373), .CO(n_1_737_814), 
      .S());
   HA_X1 i_1_737_815 (.A(\out_as[3] [6]), .B(n_1_737_374), .CO(n_1_737_815), 
      .S());
   HA_X1 i_1_737_816 (.A(\out_as[4] [6]), .B(n_1_737_375), .CO(n_1_737_816), 
      .S());
   HA_X1 i_1_737_817 (.A(\out_as[5] [6]), .B(n_1_737_376), .CO(n_1_737_817), 
      .S());
   HA_X1 i_1_737_818 (.A(\out_as[6] [6]), .B(n_1_737_377), .CO(n_1_737_818), 
      .S());
   HA_X1 i_1_737_819 (.A(\out_as[0] [6]), .B(n_1_737_378), .CO(n_1_737_819), 
      .S());
   HA_X1 i_1_737_820 (.A(\out_as[1] [6]), .B(n_1_737_379), .CO(n_1_737_820), 
      .S());
   HA_X1 i_1_737_821 (.A(\out_as[2] [6]), .B(n_1_737_380), .CO(n_1_737_821), 
      .S());
   HA_X1 i_1_737_822 (.A(\out_as[3] [6]), .B(n_1_737_381), .CO(n_1_737_822), 
      .S());
   HA_X1 i_1_737_823 (.A(\out_as[4] [6]), .B(n_1_737_382), .CO(n_1_737_823), 
      .S());
   HA_X1 i_1_737_824 (.A(\out_as[5] [6]), .B(n_1_737_383), .CO(n_1_737_824), 
      .S());
   HA_X1 i_1_737_825 (.A(\out_as[6] [6]), .B(n_1_737_384), .CO(n_1_737_825), 
      .S());
   HA_X1 i_1_737_826 (.A(\out_as[0] [6]), .B(n_1_737_385), .CO(n_1_737_826), 
      .S());
   HA_X1 i_1_737_827 (.A(\out_as[1] [6]), .B(n_1_737_386), .CO(n_1_737_827), 
      .S());
   HA_X1 i_1_737_828 (.A(\out_as[2] [6]), .B(n_1_737_387), .CO(n_1_737_828), 
      .S());
   HA_X1 i_1_737_829 (.A(\out_as[3] [6]), .B(n_1_737_388), .CO(n_1_737_829), 
      .S());
   HA_X1 i_1_737_830 (.A(\out_as[4] [6]), .B(n_1_737_389), .CO(n_1_737_830), 
      .S());
   HA_X1 i_1_737_831 (.A(\out_as[5] [6]), .B(n_1_737_390), .CO(n_1_737_831), 
      .S());
   HA_X1 i_1_737_832 (.A(\out_as[6] [6]), .B(n_1_737_391), .CO(n_1_737_832), 
      .S());
   HA_X1 i_1_737_833 (.A(\out_as[0] [6]), .B(n_1_737_392), .CO(n_1_737_833), 
      .S());
   HA_X1 i_1_737_834 (.A(\out_as[1] [6]), .B(n_1_737_393), .CO(n_1_737_834), 
      .S());
   HA_X1 i_1_737_835 (.A(\out_as[2] [6]), .B(n_1_737_394), .CO(n_1_737_835), 
      .S());
   HA_X1 i_1_737_836 (.A(\out_as[3] [6]), .B(n_1_737_395), .CO(n_1_737_836), 
      .S());
   HA_X1 i_1_737_837 (.A(\out_as[4] [6]), .B(n_1_737_396), .CO(n_1_737_837), 
      .S());
   HA_X1 i_1_737_838 (.A(\out_as[5] [6]), .B(n_1_737_397), .CO(n_1_737_838), 
      .S());
   HA_X1 i_1_737_839 (.A(\out_as[6] [6]), .B(n_1_737_398), .CO(n_1_737_839), 
      .S());
   HA_X1 i_1_737_840 (.A(\out_as[0] [6]), .B(n_1_737_399), .CO(n_1_737_840), 
      .S());
   HA_X1 i_1_737_841 (.A(\out_as[1] [6]), .B(n_1_737_400), .CO(n_1_737_841), 
      .S());
   HA_X1 i_1_737_842 (.A(\out_as[2] [6]), .B(n_1_737_401), .CO(n_1_737_842), 
      .S());
   HA_X1 i_1_737_843 (.A(\out_as[3] [6]), .B(n_1_737_402), .CO(n_1_737_843), 
      .S());
   HA_X1 i_1_737_844 (.A(\out_as[4] [6]), .B(n_1_737_403), .CO(n_1_737_844), 
      .S());
   HA_X1 i_1_737_845 (.A(\out_as[5] [6]), .B(n_1_737_404), .CO(n_1_737_845), 
      .S());
   HA_X1 i_1_737_846 (.A(\out_as[6] [6]), .B(n_1_737_405), .CO(n_1_737_846), 
      .S());
   HA_X1 i_1_737_847 (.A(\out_as[0] [6]), .B(n_1_737_406), .CO(n_1_737_847), 
      .S());
   HA_X1 i_1_737_848 (.A(\out_as[1] [6]), .B(n_1_737_407), .CO(n_1_737_848), 
      .S());
   HA_X1 i_1_737_849 (.A(\out_as[2] [6]), .B(n_1_737_408), .CO(n_1_737_849), 
      .S());
   HA_X1 i_1_737_850 (.A(\out_as[3] [6]), .B(n_1_737_409), .CO(n_1_737_850), 
      .S());
   HA_X1 i_1_737_851 (.A(\out_as[4] [6]), .B(n_1_737_410), .CO(n_1_737_851), 
      .S());
   HA_X1 i_1_737_852 (.A(\out_as[5] [6]), .B(n_1_737_411), .CO(n_1_737_852), 
      .S());
   HA_X1 i_1_737_853 (.A(\out_as[6] [6]), .B(n_1_737_412), .CO(n_1_737_853), 
      .S());
   HA_X1 i_1_737_854 (.A(\out_as[0] [6]), .B(n_1_737_413), .CO(n_1_737_854), 
      .S());
   HA_X1 i_1_737_855 (.A(\out_as[1] [6]), .B(n_1_737_414), .CO(n_1_737_855), 
      .S());
   HA_X1 i_1_737_856 (.A(\out_as[2] [6]), .B(n_1_737_415), .CO(n_1_737_856), 
      .S());
   HA_X1 i_1_737_857 (.A(\out_as[3] [6]), .B(n_1_737_416), .CO(n_1_737_857), 
      .S());
   HA_X1 i_1_737_858 (.A(\out_as[4] [6]), .B(n_1_737_417), .CO(n_1_737_858), 
      .S());
   HA_X1 i_1_737_859 (.A(\out_as[5] [6]), .B(n_1_737_418), .CO(n_1_737_859), 
      .S());
   HA_X1 i_1_737_860 (.A(\out_as[6] [6]), .B(n_1_737_419), .CO(n_1_737_860), 
      .S());
   HA_X1 i_1_737_861 (.A(\out_as[0] [6]), .B(n_1_737_420), .CO(n_1_737_861), 
      .S());
   HA_X1 i_1_737_862 (.A(\out_as[1] [6]), .B(n_1_737_421), .CO(n_1_737_862), 
      .S());
   HA_X1 i_1_737_863 (.A(\out_as[2] [6]), .B(n_1_737_422), .CO(n_1_737_863), 
      .S());
   HA_X1 i_1_737_864 (.A(\out_as[3] [6]), .B(n_1_737_423), .CO(n_1_737_864), 
      .S());
   HA_X1 i_1_737_865 (.A(\out_as[4] [6]), .B(n_1_737_424), .CO(n_1_737_865), 
      .S());
   HA_X1 i_1_737_866 (.A(\out_as[5] [6]), .B(n_1_737_425), .CO(n_1_737_866), 
      .S());
   HA_X1 i_1_737_867 (.A(\out_as[6] [6]), .B(n_1_737_426), .CO(n_1_737_867), 
      .S());
   HA_X1 i_1_737_868 (.A(\out_as[0] [6]), .B(n_1_737_427), .CO(n_1_737_868), 
      .S());
   HA_X1 i_1_737_869 (.A(\out_as[1] [6]), .B(n_1_737_428), .CO(n_1_737_869), 
      .S());
   HA_X1 i_1_737_870 (.A(\out_as[2] [6]), .B(n_1_737_429), .CO(n_1_737_870), 
      .S());
   HA_X1 i_1_737_871 (.A(\out_as[3] [6]), .B(n_1_737_430), .CO(n_1_737_871), 
      .S());
   HA_X1 i_1_737_872 (.A(\out_as[4] [6]), .B(n_1_737_431), .CO(n_1_737_872), 
      .S());
   HA_X1 i_1_737_873 (.A(\out_as[5] [6]), .B(n_1_737_432), .CO(n_1_737_873), 
      .S());
   HA_X1 i_1_737_874 (.A(\out_as[6] [6]), .B(n_1_737_433), .CO(n_1_737_874), 
      .S());
   HA_X1 i_1_737_875 (.A(\out_as[0] [6]), .B(n_1_737_434), .CO(n_1_737_875), 
      .S());
   HA_X1 i_1_737_876 (.A(\out_as[1] [6]), .B(n_1_737_435), .CO(n_1_737_876), 
      .S());
   HA_X1 i_1_737_877 (.A(\out_as[2] [6]), .B(n_1_737_436), .CO(n_1_737_877), 
      .S());
   HA_X1 i_1_737_878 (.A(\out_as[3] [6]), .B(n_1_737_437), .CO(n_1_737_878), 
      .S());
   HA_X1 i_1_737_879 (.A(\out_as[4] [6]), .B(n_1_737_438), .CO(n_1_737_879), 
      .S());
   HA_X1 i_1_737_880 (.A(\out_as[5] [6]), .B(n_1_737_439), .CO(n_1_737_880), 
      .S());
   HA_X1 i_1_737_881 (.A(\out_as[6] [6]), .B(n_1_737_440), .CO(n_1_737_881), 
      .S());
   HA_X1 i_1_737_882 (.A(\out_as[0] [6]), .B(n_1_737_441), .CO(n_1_737_882), 
      .S());
   HA_X1 i_1_737_883 (.A(\out_as[1] [6]), .B(n_1_737_442), .CO(n_1_737_883), 
      .S());
   HA_X1 i_1_737_884 (.A(\out_as[2] [6]), .B(n_1_737_443), .CO(n_1_737_884), 
      .S());
   HA_X1 i_1_737_885 (.A(\out_as[3] [6]), .B(n_1_737_444), .CO(n_1_737_885), 
      .S());
   HA_X1 i_1_737_886 (.A(\out_as[4] [6]), .B(n_1_737_445), .CO(n_1_737_886), 
      .S());
   HA_X1 i_1_737_887 (.A(\out_as[5] [6]), .B(n_1_737_446), .CO(n_1_737_887), 
      .S());
   HA_X1 i_1_737_888 (.A(\out_as[6] [6]), .B(n_1_737_447), .CO(n_1_737_888), 
      .S());
   HA_X1 i_1_737_889 (.A(\out_as[0] [6]), .B(n_1_737_448), .CO(n_1_737_889), 
      .S());
   HA_X1 i_1_737_890 (.A(\out_as[1] [6]), .B(n_1_737_449), .CO(n_1_737_890), 
      .S());
   HA_X1 i_1_737_891 (.A(\out_as[2] [6]), .B(n_1_737_450), .CO(n_1_737_891), 
      .S());
   HA_X1 i_1_737_892 (.A(\out_as[3] [6]), .B(n_1_737_451), .CO(n_1_737_892), 
      .S());
   HA_X1 i_1_737_893 (.A(\out_as[4] [6]), .B(n_1_737_452), .CO(n_1_737_893), 
      .S());
   HA_X1 i_1_737_894 (.A(\out_as[5] [6]), .B(n_1_737_453), .CO(n_1_737_894), 
      .S());
   HA_X1 i_1_737_895 (.A(\out_as[6] [6]), .B(n_1_737_454), .CO(n_1_737_895), 
      .S());
   HA_X1 i_1_737_896 (.A(\out_as[0] [6]), .B(n_1_737_455), .CO(n_1_737_896), 
      .S());
   HA_X1 i_1_737_897 (.A(\out_as[1] [6]), .B(n_1_737_456), .CO(n_1_737_897), 
      .S());
   HA_X1 i_1_737_898 (.A(\out_as[2] [6]), .B(n_1_737_457), .CO(n_1_737_898), 
      .S());
   HA_X1 i_1_737_899 (.A(\out_as[3] [6]), .B(n_1_737_458), .CO(n_1_737_899), 
      .S());
   HA_X1 i_1_737_900 (.A(\out_as[4] [6]), .B(n_1_737_459), .CO(n_1_737_900), 
      .S());
   HA_X1 i_1_737_901 (.A(\out_as[5] [6]), .B(n_1_737_460), .CO(n_1_737_901), 
      .S());
   HA_X1 i_1_737_902 (.A(\out_as[6] [6]), .B(n_1_737_461), .CO(n_1_737_902), 
      .S());
   HA_X1 i_1_737_903 (.A(\out_as[0] [6]), .B(n_1_737_462), .CO(n_1_737_903), 
      .S());
   HA_X1 i_1_737_904 (.A(\out_as[1] [6]), .B(n_1_737_463), .CO(n_1_737_904), 
      .S());
   HA_X1 i_1_737_905 (.A(\out_as[2] [6]), .B(n_1_737_464), .CO(n_1_737_905), 
      .S());
   HA_X1 i_1_737_906 (.A(\out_as[3] [6]), .B(n_1_737_465), .CO(n_1_737_906), 
      .S());
   HA_X1 i_1_737_907 (.A(\out_as[4] [6]), .B(n_1_737_466), .CO(n_1_737_907), 
      .S());
   HA_X1 i_1_737_908 (.A(\out_as[5] [6]), .B(n_1_737_467), .CO(n_1_737_908), 
      .S());
   HA_X1 i_1_737_909 (.A(\out_as[6] [6]), .B(n_1_737_468), .CO(n_1_737_909), 
      .S());
   HA_X1 i_1_737_910 (.A(\out_as[0] [6]), .B(n_1_737_469), .CO(n_1_737_910), 
      .S());
   HA_X1 i_1_737_911 (.A(\out_as[1] [6]), .B(n_1_737_470), .CO(n_1_737_911), 
      .S());
   HA_X1 i_1_737_912 (.A(\out_as[2] [6]), .B(n_1_737_471), .CO(n_1_737_912), 
      .S());
   HA_X1 i_1_737_913 (.A(\out_as[3] [6]), .B(n_1_737_472), .CO(n_1_737_913), 
      .S());
   HA_X1 i_1_737_914 (.A(\out_as[4] [6]), .B(n_1_737_473), .CO(n_1_737_914), 
      .S());
   HA_X1 i_1_737_915 (.A(\out_as[5] [6]), .B(n_1_737_474), .CO(n_1_737_915), 
      .S());
   HA_X1 i_1_737_916 (.A(\out_as[6] [6]), .B(n_1_737_475), .CO(n_1_737_916), 
      .S());
   HA_X1 i_1_737_917 (.A(\out_as[0] [6]), .B(n_1_737_476), .CO(n_1_737_917), 
      .S());
   HA_X1 i_1_737_918 (.A(\out_as[1] [6]), .B(n_1_737_477), .CO(n_1_737_918), 
      .S());
   HA_X1 i_1_737_919 (.A(\out_as[2] [6]), .B(n_1_737_478), .CO(n_1_737_919), 
      .S());
   HA_X1 i_1_737_920 (.A(\out_as[3] [6]), .B(n_1_737_479), .CO(n_1_737_920), 
      .S());
   HA_X1 i_1_737_921 (.A(\out_as[4] [6]), .B(n_1_737_480), .CO(n_1_737_921), 
      .S());
   HA_X1 i_1_737_922 (.A(\out_as[5] [6]), .B(n_1_737_481), .CO(n_1_737_922), 
      .S());
   HA_X1 i_1_737_923 (.A(\out_as[6] [6]), .B(n_1_737_482), .CO(n_1_737_923), 
      .S());
   HA_X1 i_1_737_924 (.A(\out_as[0] [6]), .B(n_1_737_483), .CO(n_1_737_924), 
      .S());
   HA_X1 i_1_737_925 (.A(\out_as[1] [6]), .B(n_1_737_484), .CO(n_1_737_925), 
      .S());
   HA_X1 i_1_737_926 (.A(\out_as[2] [6]), .B(n_1_737_485), .CO(n_1_737_926), 
      .S());
   HA_X1 i_1_737_927 (.A(\out_as[3] [6]), .B(n_1_737_486), .CO(n_1_737_927), 
      .S());
   HA_X1 i_1_737_928 (.A(\out_as[4] [6]), .B(n_1_737_487), .CO(n_1_737_928), 
      .S());
   HA_X1 i_1_737_929 (.A(\out_as[5] [6]), .B(n_1_737_488), .CO(n_1_737_929), 
      .S());
   HA_X1 i_1_737_930 (.A(\out_as[6] [6]), .B(n_1_737_489), .CO(n_1_737_930), 
      .S());
   HA_X1 i_1_737_931 (.A(\out_as[0] [6]), .B(n_1_737_490), .CO(n_1_737_931), 
      .S());
   HA_X1 i_1_737_932 (.A(\out_as[1] [6]), .B(n_1_737_491), .CO(n_1_737_932), 
      .S());
   HA_X1 i_1_737_933 (.A(\out_as[2] [6]), .B(n_1_737_492), .CO(n_1_737_933), 
      .S());
   HA_X1 i_1_737_934 (.A(\out_as[3] [6]), .B(n_1_737_493), .CO(n_1_737_934), 
      .S());
   HA_X1 i_1_737_935 (.A(\out_as[4] [6]), .B(n_1_737_494), .CO(n_1_737_935), 
      .S());
   HA_X1 i_1_737_936 (.A(\out_as[5] [6]), .B(n_1_737_495), .CO(n_1_737_936), 
      .S());
   HA_X1 i_1_737_937 (.A(\out_as[6] [6]), .B(n_1_737_496), .CO(n_1_737_937), 
      .S());
   HA_X1 i_1_737_938 (.A(\out_as[0] [6]), .B(n_1_737_497), .CO(n_1_737_938), 
      .S());
   HA_X1 i_1_737_939 (.A(\out_as[1] [6]), .B(n_1_737_498), .CO(n_1_737_939), 
      .S());
   HA_X1 i_1_737_940 (.A(\out_as[2] [6]), .B(n_1_737_499), .CO(n_1_737_940), 
      .S());
   HA_X1 i_1_737_941 (.A(\out_as[3] [6]), .B(n_1_737_500), .CO(n_1_737_941), 
      .S());
   HA_X1 i_1_737_942 (.A(\out_as[4] [6]), .B(n_1_737_501), .CO(n_1_737_942), 
      .S());
   HA_X1 i_1_737_943 (.A(\out_as[5] [6]), .B(n_1_737_502), .CO(n_1_737_943), 
      .S());
   HA_X1 i_1_737_944 (.A(\out_as[6] [6]), .B(n_1_737_503), .CO(n_1_737_944), 
      .S());
   HA_X1 i_1_737_945 (.A(\out_as[0] [6]), .B(n_1_737_504), .CO(n_1_737_945), 
      .S());
   HA_X1 i_1_737_946 (.A(\out_as[1] [6]), .B(n_1_737_505), .CO(n_1_737_946), 
      .S());
   HA_X1 i_1_737_947 (.A(\out_as[2] [6]), .B(n_1_737_506), .CO(n_1_737_947), 
      .S());
   HA_X1 i_1_737_948 (.A(\out_as[3] [6]), .B(n_1_737_507), .CO(n_1_737_948), 
      .S());
   HA_X1 i_1_737_949 (.A(\out_as[4] [6]), .B(n_1_737_508), .CO(n_1_737_949), 
      .S());
   HA_X1 i_1_737_950 (.A(\out_as[5] [6]), .B(n_1_737_509), .CO(n_1_737_950), 
      .S());
   HA_X1 i_1_737_951 (.A(\out_as[6] [6]), .B(n_1_737_510), .CO(n_1_737_951), 
      .S());
   HA_X1 i_1_737_952 (.A(\out_as[0] [6]), .B(n_1_737_511), .CO(n_1_737_952), 
      .S());
   HA_X1 i_1_737_953 (.A(\out_as[1] [6]), .B(n_1_737_512), .CO(n_1_737_953), 
      .S());
   HA_X1 i_1_737_954 (.A(\out_as[2] [6]), .B(n_1_737_513), .CO(n_1_737_954), 
      .S());
   HA_X1 i_1_737_955 (.A(\out_as[3] [6]), .B(n_1_737_514), .CO(n_1_737_955), 
      .S());
   HA_X1 i_1_737_956 (.A(\out_as[4] [6]), .B(n_1_737_515), .CO(n_1_737_956), 
      .S());
   HA_X1 i_1_737_957 (.A(\out_as[5] [6]), .B(n_1_737_516), .CO(n_1_737_957), 
      .S());
   HA_X1 i_1_737_958 (.A(\out_as[6] [6]), .B(n_1_737_517), .CO(n_1_737_958), 
      .S());
   OR2_X1 i_1_737_959 (.A1(\out_as[6] [5]), .A2(n_1_737_300), .ZN(n_1_737_959));
   OR2_X1 i_1_737_960 (.A1(\out_as[5] [5]), .A2(n_1_737_299), .ZN(n_1_737_960));
   OR2_X1 i_1_737_961 (.A1(\out_as[4] [5]), .A2(n_1_737_298), .ZN(n_1_737_961));
   OR2_X1 i_1_737_962 (.A1(\out_as[3] [5]), .A2(n_1_737_297), .ZN(n_1_737_962));
   OR2_X1 i_1_737_963 (.A1(\out_as[2] [5]), .A2(n_1_737_296), .ZN(n_1_737_963));
   OR2_X1 i_1_737_964 (.A1(\out_as[1] [5]), .A2(n_1_737_295), .ZN(n_1_737_964));
   OR2_X1 i_1_737_965 (.A1(\out_as[0] [5]), .A2(n_1_737_294), .ZN(n_1_737_965));
   OR2_X1 i_1_737_966 (.A1(\out_as[6] [5]), .A2(n_1_737_293), .ZN(n_1_737_966));
   OR2_X1 i_1_737_967 (.A1(\out_as[5] [5]), .A2(n_1_737_292), .ZN(n_1_737_967));
   OR2_X1 i_1_737_968 (.A1(\out_as[4] [5]), .A2(n_1_737_291), .ZN(n_1_737_968));
   OR2_X1 i_1_737_969 (.A1(\out_as[3] [5]), .A2(n_1_737_290), .ZN(n_1_737_969));
   OR2_X1 i_1_737_970 (.A1(\out_as[2] [5]), .A2(n_1_737_289), .ZN(n_1_737_970));
   OR2_X1 i_1_737_971 (.A1(\out_as[1] [5]), .A2(n_1_737_288), .ZN(n_1_737_971));
   OR2_X1 i_1_737_972 (.A1(\out_as[0] [5]), .A2(n_1_737_287), .ZN(n_1_737_972));
   OR2_X1 i_1_737_973 (.A1(\out_as[6] [5]), .A2(n_1_737_286), .ZN(n_1_737_973));
   OR2_X1 i_1_737_974 (.A1(\out_as[5] [5]), .A2(n_1_737_285), .ZN(n_1_737_974));
   OR2_X1 i_1_737_975 (.A1(\out_as[4] [5]), .A2(n_1_737_284), .ZN(n_1_737_975));
   OR2_X1 i_1_737_976 (.A1(\out_as[3] [5]), .A2(n_1_737_283), .ZN(n_1_737_976));
   OR2_X1 i_1_737_977 (.A1(\out_as[2] [5]), .A2(n_1_737_282), .ZN(n_1_737_977));
   OR2_X1 i_1_737_978 (.A1(\out_as[1] [5]), .A2(n_1_737_281), .ZN(n_1_737_978));
   OR2_X1 i_1_737_979 (.A1(\out_as[0] [5]), .A2(n_1_737_280), .ZN(n_1_737_979));
   OR2_X1 i_1_737_980 (.A1(\out_as[6] [5]), .A2(n_1_737_279), .ZN(n_1_737_980));
   OR2_X1 i_1_737_981 (.A1(\out_as[5] [5]), .A2(n_1_737_278), .ZN(n_1_737_981));
   OR2_X1 i_1_737_982 (.A1(\out_as[4] [5]), .A2(n_1_737_277), .ZN(n_1_737_982));
   OR2_X1 i_1_737_983 (.A1(\out_as[3] [5]), .A2(n_1_737_276), .ZN(n_1_737_983));
   OR2_X1 i_1_737_984 (.A1(\out_as[2] [5]), .A2(n_1_737_275), .ZN(n_1_737_984));
   OR2_X1 i_1_737_985 (.A1(\out_as[1] [5]), .A2(n_1_737_274), .ZN(n_1_737_985));
   OR2_X1 i_1_737_986 (.A1(\out_as[0] [5]), .A2(n_1_737_273), .ZN(n_1_737_986));
   OR2_X1 i_1_737_987 (.A1(\out_as[6] [5]), .A2(n_1_737_272), .ZN(n_1_737_987));
   OR2_X1 i_1_737_988 (.A1(\out_as[5] [5]), .A2(n_1_737_271), .ZN(n_1_737_988));
   OR2_X1 i_1_737_989 (.A1(\out_as[4] [5]), .A2(n_1_737_270), .ZN(n_1_737_989));
   OR2_X1 i_1_737_990 (.A1(\out_as[3] [5]), .A2(n_1_737_269), .ZN(n_1_737_990));
   OR2_X1 i_1_737_991 (.A1(\out_as[2] [5]), .A2(n_1_737_268), .ZN(n_1_737_991));
   OR2_X1 i_1_737_992 (.A1(\out_as[1] [5]), .A2(n_1_737_267), .ZN(n_1_737_992));
   OR2_X1 i_1_737_993 (.A1(\out_as[0] [5]), .A2(n_1_737_266), .ZN(n_1_737_993));
   OR2_X1 i_1_737_994 (.A1(\out_as[6] [5]), .A2(n_1_737_265), .ZN(n_1_737_994));
   OR2_X1 i_1_737_995 (.A1(\out_as[5] [5]), .A2(n_1_737_264), .ZN(n_1_737_995));
   OR2_X1 i_1_737_996 (.A1(\out_as[4] [5]), .A2(n_1_737_263), .ZN(n_1_737_996));
   OR2_X1 i_1_737_997 (.A1(\out_as[3] [5]), .A2(n_1_737_262), .ZN(n_1_737_997));
   OR2_X1 i_1_737_998 (.A1(\out_as[2] [5]), .A2(n_1_737_261), .ZN(n_1_737_998));
   OR2_X1 i_1_737_999 (.A1(\out_as[1] [5]), .A2(n_1_737_260), .ZN(n_1_737_999));
   OR2_X1 i_1_737_1000 (.A1(\out_as[0] [5]), .A2(n_1_737_259), .ZN(n_1_737_1000));
   OR2_X1 i_1_737_1001 (.A1(\out_as[6] [5]), .A2(n_1_737_258), .ZN(n_1_737_1001));
   OR2_X1 i_1_737_1002 (.A1(\out_as[5] [5]), .A2(n_1_737_257), .ZN(n_1_737_1002));
   OR2_X1 i_1_737_1003 (.A1(\out_as[4] [5]), .A2(n_1_737_256), .ZN(n_1_737_1003));
   OR2_X1 i_1_737_1004 (.A1(\out_as[3] [5]), .A2(n_1_737_255), .ZN(n_1_737_1004));
   OR2_X1 i_1_737_1005 (.A1(\out_as[2] [5]), .A2(n_1_737_254), .ZN(n_1_737_1005));
   OR2_X1 i_1_737_1006 (.A1(\out_as[1] [5]), .A2(n_1_737_253), .ZN(n_1_737_1006));
   OR2_X1 i_1_737_1007 (.A1(\out_as[0] [5]), .A2(n_1_737_252), .ZN(n_1_737_1007));
   OR2_X1 i_1_737_1008 (.A1(\out_as[6] [5]), .A2(n_1_737_251), .ZN(n_1_737_1008));
   OR2_X1 i_1_737_1009 (.A1(\out_as[5] [5]), .A2(n_1_737_250), .ZN(n_1_737_1009));
   OR2_X1 i_1_737_1010 (.A1(\out_as[4] [5]), .A2(n_1_737_249), .ZN(n_1_737_1010));
   OR2_X1 i_1_737_1011 (.A1(\out_as[3] [5]), .A2(n_1_737_248), .ZN(n_1_737_1011));
   OR2_X1 i_1_737_1012 (.A1(\out_as[2] [5]), .A2(n_1_737_247), .ZN(n_1_737_1012));
   OR2_X1 i_1_737_1013 (.A1(\out_as[1] [5]), .A2(n_1_737_246), .ZN(n_1_737_1013));
   OR2_X1 i_1_737_1014 (.A1(\out_as[0] [5]), .A2(n_1_737_245), .ZN(n_1_737_1014));
   OR2_X1 i_1_737_1015 (.A1(\out_as[6] [5]), .A2(n_1_737_244), .ZN(n_1_737_1015));
   OR2_X1 i_1_737_1016 (.A1(\out_as[5] [5]), .A2(n_1_737_243), .ZN(n_1_737_1016));
   OR2_X1 i_1_737_1017 (.A1(\out_as[4] [5]), .A2(n_1_737_242), .ZN(n_1_737_1017));
   OR2_X1 i_1_737_1018 (.A1(\out_as[3] [5]), .A2(n_1_737_241), .ZN(n_1_737_1018));
   OR2_X1 i_1_737_1019 (.A1(\out_as[2] [5]), .A2(n_1_737_240), .ZN(n_1_737_1019));
   OR2_X1 i_1_737_1020 (.A1(\out_as[1] [5]), .A2(n_1_737_239), .ZN(n_1_737_1020));
   OR2_X1 i_1_737_1021 (.A1(\out_as[0] [5]), .A2(n_1_737_238), .ZN(n_1_737_1021));
   OR2_X1 i_1_737_1022 (.A1(\out_as[6] [5]), .A2(n_1_737_237), .ZN(n_1_737_1022));
   OR2_X1 i_1_737_1023 (.A1(\out_as[5] [5]), .A2(n_1_737_236), .ZN(n_1_737_1023));
   OR2_X1 i_1_737_1024 (.A1(\out_as[4] [5]), .A2(n_1_737_235), .ZN(n_1_737_1024));
   OR2_X1 i_1_737_1025 (.A1(\out_as[3] [5]), .A2(n_1_737_234), .ZN(n_1_737_1025));
   OR2_X1 i_1_737_1026 (.A1(\out_as[2] [5]), .A2(n_1_737_233), .ZN(n_1_737_1026));
   OR2_X1 i_1_737_1027 (.A1(\out_as[1] [5]), .A2(n_1_737_232), .ZN(n_1_737_1027));
   OR2_X1 i_1_737_1028 (.A1(\out_as[0] [5]), .A2(n_1_737_231), .ZN(n_1_737_1028));
   OR2_X1 i_1_737_1029 (.A1(\out_as[6] [5]), .A2(n_1_737_230), .ZN(n_1_737_1029));
   OR2_X1 i_1_737_1030 (.A1(\out_as[5] [5]), .A2(n_1_737_229), .ZN(n_1_737_1030));
   OR2_X1 i_1_737_1031 (.A1(\out_as[4] [5]), .A2(n_1_737_228), .ZN(n_1_737_1031));
   OR2_X1 i_1_737_1032 (.A1(\out_as[3] [5]), .A2(n_1_737_227), .ZN(n_1_737_1032));
   OR2_X1 i_1_737_1033 (.A1(\out_as[2] [5]), .A2(n_1_737_226), .ZN(n_1_737_1033));
   OR2_X1 i_1_737_1034 (.A1(\out_as[1] [5]), .A2(n_1_737_225), .ZN(n_1_737_1034));
   OR2_X1 i_1_737_1035 (.A1(\out_as[0] [5]), .A2(n_1_737_224), .ZN(n_1_737_1035));
   OR2_X1 i_1_737_1036 (.A1(\out_as[6] [5]), .A2(n_1_737_223), .ZN(n_1_737_1036));
   OR2_X1 i_1_737_1037 (.A1(\out_as[5] [5]), .A2(n_1_737_222), .ZN(n_1_737_1037));
   OR2_X1 i_1_737_1038 (.A1(\out_as[4] [5]), .A2(n_1_737_221), .ZN(n_1_737_1038));
   OR2_X1 i_1_737_1039 (.A1(\out_as[3] [5]), .A2(n_1_737_220), .ZN(n_1_737_1039));
   OR2_X1 i_1_737_1040 (.A1(\out_as[2] [5]), .A2(n_1_737_219), .ZN(n_1_737_1040));
   OR2_X1 i_1_737_1041 (.A1(\out_as[1] [5]), .A2(n_1_737_218), .ZN(n_1_737_1041));
   OR2_X1 i_1_737_1042 (.A1(\out_as[0] [5]), .A2(n_1_737_217), .ZN(n_1_737_1042));
   OR2_X1 i_1_737_1043 (.A1(\out_as[6] [5]), .A2(n_1_737_216), .ZN(n_1_737_1043));
   OR2_X1 i_1_737_1044 (.A1(\out_as[5] [5]), .A2(n_1_737_215), .ZN(n_1_737_1044));
   OR2_X1 i_1_737_1045 (.A1(\out_as[4] [5]), .A2(n_1_737_214), .ZN(n_1_737_1045));
   OR2_X1 i_1_737_1046 (.A1(\out_as[3] [5]), .A2(n_1_737_213), .ZN(n_1_737_1046));
   OR2_X1 i_1_737_1047 (.A1(\out_as[2] [5]), .A2(n_1_737_212), .ZN(n_1_737_1047));
   OR2_X1 i_1_737_1048 (.A1(\out_as[1] [5]), .A2(n_1_737_211), .ZN(n_1_737_1048));
   OR2_X1 i_1_737_1049 (.A1(\out_as[0] [5]), .A2(n_1_737_210), .ZN(n_1_737_1049));
   OR2_X1 i_1_737_1050 (.A1(\out_as[6] [5]), .A2(n_1_737_209), .ZN(n_1_737_1050));
   OR2_X1 i_1_737_1051 (.A1(\out_as[5] [5]), .A2(n_1_737_208), .ZN(n_1_737_1051));
   OR2_X1 i_1_737_1052 (.A1(\out_as[4] [5]), .A2(n_1_737_207), .ZN(n_1_737_1052));
   OR2_X1 i_1_737_1053 (.A1(\out_as[3] [5]), .A2(n_1_737_206), .ZN(n_1_737_1053));
   OR2_X1 i_1_737_1054 (.A1(\out_as[2] [5]), .A2(n_1_737_205), .ZN(n_1_737_1054));
   OR2_X1 i_1_737_1055 (.A1(\out_as[1] [5]), .A2(n_1_737_204), .ZN(n_1_737_1055));
   OR2_X1 i_1_737_1056 (.A1(\out_as[0] [5]), .A2(n_1_737_203), .ZN(n_1_737_1056));
   OR2_X1 i_1_737_1057 (.A1(\out_as[6] [5]), .A2(n_1_737_202), .ZN(n_1_737_1057));
   OR2_X1 i_1_737_1058 (.A1(\out_as[5] [5]), .A2(n_1_737_201), .ZN(n_1_737_1058));
   OR2_X1 i_1_737_1059 (.A1(\out_as[4] [5]), .A2(n_1_737_200), .ZN(n_1_737_1059));
   OR2_X1 i_1_737_1060 (.A1(\out_as[3] [5]), .A2(n_1_737_199), .ZN(n_1_737_1060));
   OR2_X1 i_1_737_1061 (.A1(\out_as[2] [5]), .A2(n_1_737_198), .ZN(n_1_737_1061));
   OR2_X1 i_1_737_1062 (.A1(\out_as[1] [5]), .A2(n_1_737_197), .ZN(n_1_737_1062));
   OR2_X1 i_1_737_1063 (.A1(\out_as[0] [5]), .A2(n_1_737_196), .ZN(n_1_737_1063));
   OR2_X1 i_1_737_1064 (.A1(n_1_737_195), .A2(n_1_737_5156), .ZN(n_1_737_1064));
   OR2_X1 i_1_737_1065 (.A1(n_1_737_194), .A2(n_1_737_5169), .ZN(n_1_737_1065));
   OR2_X1 i_1_737_1066 (.A1(n_1_737_193), .A2(n_1_737_5388), .ZN(n_1_737_1066));
   OR2_X1 i_1_737_1067 (.A1(n_1_737_192), .A2(n_1_737_5217), .ZN(n_1_737_1067));
   OR2_X1 i_1_737_1068 (.A1(n_1_737_191), .A2(n_1_737_5276), .ZN(n_1_737_1068));
   OR2_X1 i_1_737_1069 (.A1(n_1_737_190), .A2(n_1_737_5322), .ZN(n_1_737_1069));
   OR2_X1 i_1_737_1070 (.A1(n_1_737_189), .A2(n_1_737_5360), .ZN(n_1_737_1070));
   OR2_X1 i_1_737_1071 (.A1(n_1_737_188), .A2(n_1_737_5156), .ZN(n_1_737_1071));
   OR2_X1 i_1_737_1072 (.A1(n_1_737_187), .A2(n_1_737_5169), .ZN(n_1_737_1072));
   OR2_X1 i_1_737_1073 (.A1(n_1_737_186), .A2(n_1_737_5388), .ZN(n_1_737_1073));
   OR2_X1 i_1_737_1074 (.A1(n_1_737_185), .A2(n_1_737_5217), .ZN(n_1_737_1074));
   OR2_X1 i_1_737_1075 (.A1(n_1_737_184), .A2(n_1_737_5276), .ZN(n_1_737_1075));
   OR2_X1 i_1_737_1076 (.A1(n_1_737_183), .A2(n_1_737_5322), .ZN(n_1_737_1076));
   OR2_X1 i_1_737_1077 (.A1(n_1_737_182), .A2(n_1_737_5360), .ZN(n_1_737_1077));
   OR2_X1 i_1_737_1078 (.A1(n_1_737_181), .A2(n_1_737_5156), .ZN(n_1_737_1078));
   OR2_X1 i_1_737_1079 (.A1(n_1_737_180), .A2(n_1_737_5169), .ZN(n_1_737_1079));
   OR2_X1 i_1_737_1080 (.A1(n_1_737_179), .A2(n_1_737_5388), .ZN(n_1_737_1080));
   OR2_X1 i_1_737_1081 (.A1(n_1_737_178), .A2(n_1_737_5217), .ZN(n_1_737_1081));
   OR2_X1 i_1_737_1082 (.A1(n_1_737_177), .A2(n_1_737_5276), .ZN(n_1_737_1082));
   OR2_X1 i_1_737_1083 (.A1(n_1_737_176), .A2(n_1_737_5322), .ZN(n_1_737_1083));
   OR2_X1 i_1_737_1084 (.A1(n_1_737_175), .A2(n_1_737_5360), .ZN(n_1_737_1084));
   OR2_X1 i_1_737_1085 (.A1(n_1_737_174), .A2(n_1_737_5156), .ZN(n_1_737_1085));
   OR2_X1 i_1_737_1086 (.A1(n_1_737_173), .A2(n_1_737_5169), .ZN(n_1_737_1086));
   OR2_X1 i_1_737_1087 (.A1(n_1_737_172), .A2(n_1_737_5388), .ZN(n_1_737_1087));
   OR2_X1 i_1_737_1088 (.A1(n_1_737_171), .A2(n_1_737_5217), .ZN(n_1_737_1088));
   OR2_X1 i_1_737_1089 (.A1(n_1_737_170), .A2(n_1_737_5276), .ZN(n_1_737_1089));
   OR2_X1 i_1_737_1090 (.A1(n_1_737_169), .A2(n_1_737_5322), .ZN(n_1_737_1090));
   OR2_X1 i_1_737_1091 (.A1(n_1_737_168), .A2(n_1_737_5360), .ZN(n_1_737_1091));
   OR2_X1 i_1_737_1092 (.A1(n_1_737_167), .A2(n_1_737_5156), .ZN(n_1_737_1092));
   OR2_X1 i_1_737_1093 (.A1(n_1_737_166), .A2(n_1_737_5169), .ZN(n_1_737_1093));
   OR2_X1 i_1_737_1094 (.A1(n_1_737_165), .A2(n_1_737_5388), .ZN(n_1_737_1094));
   OR2_X1 i_1_737_1095 (.A1(n_1_737_164), .A2(n_1_737_5217), .ZN(n_1_737_1095));
   OR2_X1 i_1_737_1096 (.A1(n_1_737_163), .A2(n_1_737_5276), .ZN(n_1_737_1096));
   OR2_X1 i_1_737_1097 (.A1(n_1_737_162), .A2(n_1_737_5322), .ZN(n_1_737_1097));
   OR2_X1 i_1_737_1098 (.A1(n_1_737_161), .A2(n_1_737_5360), .ZN(n_1_737_1098));
   OR2_X1 i_1_737_1099 (.A1(n_1_737_160), .A2(n_1_737_5156), .ZN(n_1_737_1099));
   OR2_X1 i_1_737_1100 (.A1(n_1_737_159), .A2(n_1_737_5169), .ZN(n_1_737_1100));
   OR2_X1 i_1_737_1101 (.A1(n_1_737_158), .A2(n_1_737_5388), .ZN(n_1_737_1101));
   OR2_X1 i_1_737_1102 (.A1(n_1_737_157), .A2(n_1_737_5217), .ZN(n_1_737_1102));
   OR2_X1 i_1_737_1103 (.A1(n_1_737_156), .A2(n_1_737_5276), .ZN(n_1_737_1103));
   OR2_X1 i_1_737_1104 (.A1(n_1_737_155), .A2(n_1_737_5322), .ZN(n_1_737_1104));
   OR2_X1 i_1_737_1105 (.A1(n_1_737_154), .A2(n_1_737_5360), .ZN(n_1_737_1105));
   OR2_X1 i_1_737_1106 (.A1(n_1_737_153), .A2(n_1_737_5156), .ZN(n_1_737_1106));
   OR2_X1 i_1_737_1107 (.A1(n_1_737_152), .A2(n_1_737_5169), .ZN(n_1_737_1107));
   OR2_X1 i_1_737_1108 (.A1(n_1_737_151), .A2(n_1_737_5388), .ZN(n_1_737_1108));
   OR2_X1 i_1_737_1109 (.A1(n_1_737_150), .A2(n_1_737_5217), .ZN(n_1_737_1109));
   OR2_X1 i_1_737_1110 (.A1(n_1_737_149), .A2(n_1_737_5276), .ZN(n_1_737_1110));
   OR2_X1 i_1_737_1111 (.A1(n_1_737_148), .A2(n_1_737_5322), .ZN(n_1_737_1111));
   OR2_X1 i_1_737_1112 (.A1(n_1_737_147), .A2(n_1_737_5360), .ZN(n_1_737_1112));
   OR2_X1 i_1_737_1113 (.A1(n_1_737_146), .A2(n_1_737_5152), .ZN(n_1_737_1113));
   OR2_X1 i_1_737_1114 (.A1(n_1_737_145), .A2(n_1_737_5164), .ZN(n_1_737_1114));
   OR2_X1 i_1_737_1115 (.A1(n_1_737_144), .A2(n_1_737_5383), .ZN(n_1_737_1115));
   OR2_X1 i_1_737_1116 (.A1(n_1_737_143), .A2(n_1_737_5211), .ZN(n_1_737_1116));
   OR2_X1 i_1_737_1117 (.A1(n_1_737_142), .A2(n_1_737_5271), .ZN(n_1_737_1117));
   OR2_X1 i_1_737_1118 (.A1(n_1_737_141), .A2(n_1_737_5316), .ZN(n_1_737_1118));
   OR2_X1 i_1_737_1119 (.A1(n_1_737_140), .A2(n_1_737_5354), .ZN(n_1_737_1119));
   OR2_X1 i_1_737_1120 (.A1(n_1_737_139), .A2(n_1_737_5152), .ZN(n_1_737_1120));
   OR2_X1 i_1_737_1121 (.A1(n_1_737_138), .A2(n_1_737_5164), .ZN(n_1_737_1121));
   OR2_X1 i_1_737_1122 (.A1(n_1_737_137), .A2(n_1_737_5383), .ZN(n_1_737_1122));
   OR2_X1 i_1_737_1123 (.A1(n_1_737_136), .A2(n_1_737_5211), .ZN(n_1_737_1123));
   OR2_X1 i_1_737_1124 (.A1(n_1_737_135), .A2(n_1_737_5271), .ZN(n_1_737_1124));
   OR2_X1 i_1_737_1125 (.A1(n_1_737_134), .A2(n_1_737_5316), .ZN(n_1_737_1125));
   OR2_X1 i_1_737_1126 (.A1(n_1_737_133), .A2(n_1_737_5354), .ZN(n_1_737_1126));
   OR2_X1 i_1_737_1127 (.A1(n_1_737_132), .A2(n_1_737_5152), .ZN(n_1_737_1127));
   OR2_X1 i_1_737_1128 (.A1(n_1_737_131), .A2(n_1_737_5164), .ZN(n_1_737_1128));
   OR2_X1 i_1_737_1129 (.A1(n_1_737_130), .A2(n_1_737_5383), .ZN(n_1_737_1129));
   OR2_X1 i_1_737_1130 (.A1(n_1_737_129), .A2(n_1_737_5211), .ZN(n_1_737_1130));
   OR2_X1 i_1_737_1131 (.A1(n_1_737_128), .A2(n_1_737_5271), .ZN(n_1_737_1131));
   OR2_X1 i_1_737_1132 (.A1(n_1_737_127), .A2(n_1_737_5316), .ZN(n_1_737_1132));
   OR2_X1 i_1_737_1133 (.A1(n_1_737_126), .A2(n_1_737_5354), .ZN(n_1_737_1133));
   OR2_X1 i_1_737_1134 (.A1(n_1_737_125), .A2(n_1_737_5067), .ZN(n_1_737_1134));
   OR2_X1 i_1_737_1135 (.A1(n_1_737_124), .A2(n_1_737_5070), .ZN(n_1_737_1135));
   OR2_X1 i_1_737_1136 (.A1(n_1_737_123), .A2(n_1_737_5136), .ZN(n_1_737_1136));
   OR2_X1 i_1_737_1137 (.A1(n_1_737_122), .A2(n_1_737_5118), .ZN(n_1_737_1137));
   OR2_X1 i_1_737_1138 (.A1(n_1_737_121), .A2(n_1_737_5101), .ZN(n_1_737_1138));
   OR2_X1 i_1_737_1139 (.A1(n_1_737_120), .A2(n_1_737_5108), .ZN(n_1_737_1139));
   OR2_X1 i_1_737_1140 (.A1(n_1_737_119), .A2(n_1_737_5088), .ZN(n_1_737_1140));
   OR2_X1 i_1_737_1141 (.A1(n_1_737_5070), .A2(n_1_737_2013), .ZN(n_1_737_1141));
   OR2_X1 i_1_737_1142 (.A1(\out_as[4] [5]), .A2(n_1_737_1999), .ZN(n_1_737_1142));
   OR2_X1 i_1_737_1143 (.A1(\out_as[3] [5]), .A2(n_1_737_2016), .ZN(n_1_737_1143));
   OR2_X1 i_1_737_1144 (.A1(\out_as[2] [5]), .A2(n_1_737_1988), .ZN(n_1_737_1144));
   OR2_X1 i_1_737_1145 (.A1(\out_as[1] [5]), .A2(n_1_737_1994), .ZN(n_1_737_1145));
   OR2_X1 i_1_737_1146 (.A1(\out_as[0] [5]), .A2(n_1_737_2005), .ZN(n_1_737_1146));
   OR2_X1 i_1_737_1147 (.A1(\out_as[6] [4]), .A2(n_1_737_195), .ZN(n_1_737_1147));
   OR2_X1 i_1_737_1148 (.A1(\out_as[5] [4]), .A2(n_1_737_194), .ZN(n_1_737_1148));
   OR2_X1 i_1_737_1149 (.A1(\out_as[4] [4]), .A2(n_1_737_193), .ZN(n_1_737_1149));
   OR2_X1 i_1_737_1150 (.A1(\out_as[3] [4]), .A2(n_1_737_192), .ZN(n_1_737_1150));
   OR2_X1 i_1_737_1151 (.A1(\out_as[2] [4]), .A2(n_1_737_191), .ZN(n_1_737_1151));
   OR2_X1 i_1_737_1152 (.A1(\out_as[1] [4]), .A2(n_1_737_190), .ZN(n_1_737_1152));
   OR2_X1 i_1_737_1153 (.A1(\out_as[0] [4]), .A2(n_1_737_189), .ZN(n_1_737_1153));
   OR2_X1 i_1_737_1154 (.A1(\out_as[6] [4]), .A2(n_1_737_188), .ZN(n_1_737_1154));
   OR2_X1 i_1_737_1155 (.A1(\out_as[5] [4]), .A2(n_1_737_187), .ZN(n_1_737_1155));
   OR2_X1 i_1_737_1156 (.A1(\out_as[4] [4]), .A2(n_1_737_186), .ZN(n_1_737_1156));
   OR2_X1 i_1_737_1157 (.A1(\out_as[3] [4]), .A2(n_1_737_185), .ZN(n_1_737_1157));
   OR2_X1 i_1_737_1158 (.A1(\out_as[2] [4]), .A2(n_1_737_184), .ZN(n_1_737_1158));
   OR2_X1 i_1_737_1159 (.A1(\out_as[1] [4]), .A2(n_1_737_183), .ZN(n_1_737_1159));
   OR2_X1 i_1_737_1160 (.A1(\out_as[0] [4]), .A2(n_1_737_182), .ZN(n_1_737_1160));
   OR2_X1 i_1_737_1161 (.A1(\out_as[6] [4]), .A2(n_1_737_181), .ZN(n_1_737_1161));
   OR2_X1 i_1_737_1162 (.A1(\out_as[5] [4]), .A2(n_1_737_180), .ZN(n_1_737_1162));
   OR2_X1 i_1_737_1163 (.A1(\out_as[4] [4]), .A2(n_1_737_179), .ZN(n_1_737_1163));
   OR2_X1 i_1_737_1164 (.A1(\out_as[3] [4]), .A2(n_1_737_178), .ZN(n_1_737_1164));
   OR2_X1 i_1_737_1165 (.A1(\out_as[2] [4]), .A2(n_1_737_177), .ZN(n_1_737_1165));
   OR2_X1 i_1_737_1166 (.A1(\out_as[1] [4]), .A2(n_1_737_176), .ZN(n_1_737_1166));
   OR2_X1 i_1_737_1167 (.A1(\out_as[0] [4]), .A2(n_1_737_175), .ZN(n_1_737_1167));
   OR2_X1 i_1_737_1168 (.A1(\out_as[6] [4]), .A2(n_1_737_174), .ZN(n_1_737_1168));
   OR2_X1 i_1_737_1169 (.A1(\out_as[5] [4]), .A2(n_1_737_173), .ZN(n_1_737_1169));
   OR2_X1 i_1_737_1170 (.A1(\out_as[4] [4]), .A2(n_1_737_172), .ZN(n_1_737_1170));
   OR2_X1 i_1_737_1171 (.A1(\out_as[3] [4]), .A2(n_1_737_171), .ZN(n_1_737_1171));
   OR2_X1 i_1_737_1172 (.A1(\out_as[2] [4]), .A2(n_1_737_170), .ZN(n_1_737_1172));
   OR2_X1 i_1_737_1173 (.A1(\out_as[1] [4]), .A2(n_1_737_169), .ZN(n_1_737_1173));
   OR2_X1 i_1_737_1174 (.A1(\out_as[0] [4]), .A2(n_1_737_168), .ZN(n_1_737_1174));
   OR2_X1 i_1_737_1175 (.A1(\out_as[6] [4]), .A2(n_1_737_167), .ZN(n_1_737_1175));
   OR2_X1 i_1_737_1176 (.A1(\out_as[5] [4]), .A2(n_1_737_166), .ZN(n_1_737_1176));
   OR2_X1 i_1_737_1177 (.A1(\out_as[4] [4]), .A2(n_1_737_165), .ZN(n_1_737_1177));
   OR2_X1 i_1_737_1178 (.A1(\out_as[3] [4]), .A2(n_1_737_164), .ZN(n_1_737_1178));
   OR2_X1 i_1_737_1179 (.A1(\out_as[2] [4]), .A2(n_1_737_163), .ZN(n_1_737_1179));
   OR2_X1 i_1_737_1180 (.A1(\out_as[1] [4]), .A2(n_1_737_162), .ZN(n_1_737_1180));
   OR2_X1 i_1_737_1181 (.A1(\out_as[0] [4]), .A2(n_1_737_161), .ZN(n_1_737_1181));
   OR2_X1 i_1_737_1182 (.A1(\out_as[6] [4]), .A2(n_1_737_160), .ZN(n_1_737_1182));
   OR2_X1 i_1_737_1183 (.A1(\out_as[5] [4]), .A2(n_1_737_159), .ZN(n_1_737_1183));
   OR2_X1 i_1_737_1184 (.A1(\out_as[4] [4]), .A2(n_1_737_158), .ZN(n_1_737_1184));
   OR2_X1 i_1_737_1185 (.A1(\out_as[3] [4]), .A2(n_1_737_157), .ZN(n_1_737_1185));
   OR2_X1 i_1_737_1186 (.A1(\out_as[2] [4]), .A2(n_1_737_156), .ZN(n_1_737_1186));
   OR2_X1 i_1_737_1187 (.A1(\out_as[1] [4]), .A2(n_1_737_155), .ZN(n_1_737_1187));
   OR2_X1 i_1_737_1188 (.A1(\out_as[0] [4]), .A2(n_1_737_154), .ZN(n_1_737_1188));
   OR2_X1 i_1_737_1189 (.A1(\out_as[6] [4]), .A2(n_1_737_153), .ZN(n_1_737_1189));
   OR2_X1 i_1_737_1190 (.A1(\out_as[5] [4]), .A2(n_1_737_152), .ZN(n_1_737_1190));
   OR2_X1 i_1_737_1191 (.A1(\out_as[4] [4]), .A2(n_1_737_151), .ZN(n_1_737_1191));
   OR2_X1 i_1_737_1192 (.A1(\out_as[3] [4]), .A2(n_1_737_150), .ZN(n_1_737_1192));
   OR2_X1 i_1_737_1193 (.A1(\out_as[2] [4]), .A2(n_1_737_149), .ZN(n_1_737_1193));
   OR2_X1 i_1_737_1194 (.A1(\out_as[1] [4]), .A2(n_1_737_148), .ZN(n_1_737_1194));
   OR2_X1 i_1_737_1195 (.A1(\out_as[0] [4]), .A2(n_1_737_147), .ZN(n_1_737_1195));
   OR2_X1 i_1_737_1196 (.A1(n_1_737_146), .A2(n_1_737_5153), .ZN(n_1_737_1196));
   OR2_X1 i_1_737_1197 (.A1(n_1_737_145), .A2(n_1_737_5165), .ZN(n_1_737_1197));
   OR2_X1 i_1_737_1198 (.A1(n_1_737_144), .A2(n_1_737_5384), .ZN(n_1_737_1198));
   OR2_X1 i_1_737_1199 (.A1(n_1_737_143), .A2(n_1_737_5212), .ZN(n_1_737_1199));
   OR2_X1 i_1_737_1200 (.A1(n_1_737_142), .A2(n_1_737_5272), .ZN(n_1_737_1200));
   OR2_X1 i_1_737_1201 (.A1(n_1_737_141), .A2(n_1_737_5317), .ZN(n_1_737_1201));
   OR2_X1 i_1_737_1202 (.A1(n_1_737_140), .A2(n_1_737_5355), .ZN(n_1_737_1202));
   OR2_X1 i_1_737_1203 (.A1(n_1_737_139), .A2(n_1_737_5153), .ZN(n_1_737_1203));
   OR2_X1 i_1_737_1204 (.A1(n_1_737_138), .A2(n_1_737_5165), .ZN(n_1_737_1204));
   OR2_X1 i_1_737_1205 (.A1(n_1_737_137), .A2(n_1_737_5384), .ZN(n_1_737_1205));
   OR2_X1 i_1_737_1206 (.A1(n_1_737_136), .A2(n_1_737_5212), .ZN(n_1_737_1206));
   OR2_X1 i_1_737_1207 (.A1(n_1_737_135), .A2(n_1_737_5272), .ZN(n_1_737_1207));
   OR2_X1 i_1_737_1208 (.A1(n_1_737_134), .A2(n_1_737_5317), .ZN(n_1_737_1208));
   OR2_X1 i_1_737_1209 (.A1(n_1_737_133), .A2(n_1_737_5355), .ZN(n_1_737_1209));
   OR2_X1 i_1_737_1210 (.A1(n_1_737_132), .A2(n_1_737_5153), .ZN(n_1_737_1210));
   OR2_X1 i_1_737_1211 (.A1(n_1_737_131), .A2(n_1_737_5165), .ZN(n_1_737_1211));
   OR2_X1 i_1_737_1212 (.A1(n_1_737_130), .A2(n_1_737_5384), .ZN(n_1_737_1212));
   OR2_X1 i_1_737_1213 (.A1(n_1_737_129), .A2(n_1_737_5212), .ZN(n_1_737_1213));
   OR2_X1 i_1_737_1214 (.A1(n_1_737_128), .A2(n_1_737_5272), .ZN(n_1_737_1214));
   OR2_X1 i_1_737_1215 (.A1(n_1_737_127), .A2(n_1_737_5317), .ZN(n_1_737_1215));
   OR2_X1 i_1_737_1216 (.A1(n_1_737_126), .A2(n_1_737_5355), .ZN(n_1_737_1216));
   OR2_X1 i_1_737_1217 (.A1(n_1_737_125), .A2(n_1_737_5148), .ZN(n_1_737_1217));
   OR2_X1 i_1_737_1218 (.A1(n_1_737_124), .A2(n_1_737_5160), .ZN(n_1_737_1218));
   OR2_X1 i_1_737_1219 (.A1(n_1_737_123), .A2(n_1_737_5379), .ZN(n_1_737_1219));
   OR2_X1 i_1_737_1220 (.A1(n_1_737_122), .A2(n_1_737_5206), .ZN(n_1_737_1220));
   OR2_X1 i_1_737_1221 (.A1(n_1_737_121), .A2(n_1_737_5267), .ZN(n_1_737_1221));
   OR2_X1 i_1_737_1222 (.A1(n_1_737_120), .A2(n_1_737_5311), .ZN(n_1_737_1222));
   OR2_X1 i_1_737_1223 (.A1(n_1_737_119), .A2(n_1_737_5349), .ZN(n_1_737_1223));
   OR2_X1 i_1_737_1224 (.A1(\out_as[6] [3]), .A2(n_1_737_146), .ZN(n_1_737_1224));
   OR2_X1 i_1_737_1225 (.A1(\out_as[5] [3]), .A2(n_1_737_145), .ZN(n_1_737_1225));
   OR2_X1 i_1_737_1226 (.A1(\out_as[4] [3]), .A2(n_1_737_144), .ZN(n_1_737_1226));
   OR2_X1 i_1_737_1227 (.A1(\out_as[3] [3]), .A2(n_1_737_143), .ZN(n_1_737_1227));
   OR2_X1 i_1_737_1228 (.A1(\out_as[2] [3]), .A2(n_1_737_142), .ZN(n_1_737_1228));
   OR2_X1 i_1_737_1229 (.A1(\out_as[1] [3]), .A2(n_1_737_141), .ZN(n_1_737_1229));
   OR2_X1 i_1_737_1230 (.A1(\out_as[0] [3]), .A2(n_1_737_140), .ZN(n_1_737_1230));
   OR2_X1 i_1_737_1231 (.A1(\out_as[6] [3]), .A2(n_1_737_139), .ZN(n_1_737_1231));
   OR2_X1 i_1_737_1232 (.A1(\out_as[5] [3]), .A2(n_1_737_138), .ZN(n_1_737_1232));
   OR2_X1 i_1_737_1233 (.A1(\out_as[4] [3]), .A2(n_1_737_137), .ZN(n_1_737_1233));
   OR2_X1 i_1_737_1234 (.A1(\out_as[3] [3]), .A2(n_1_737_136), .ZN(n_1_737_1234));
   OR2_X1 i_1_737_1235 (.A1(\out_as[2] [3]), .A2(n_1_737_135), .ZN(n_1_737_1235));
   OR2_X1 i_1_737_1236 (.A1(\out_as[1] [3]), .A2(n_1_737_134), .ZN(n_1_737_1236));
   OR2_X1 i_1_737_1237 (.A1(\out_as[0] [3]), .A2(n_1_737_133), .ZN(n_1_737_1237));
   OR2_X1 i_1_737_1238 (.A1(\out_as[6] [3]), .A2(n_1_737_132), .ZN(n_1_737_1238));
   OR2_X1 i_1_737_1239 (.A1(\out_as[5] [3]), .A2(n_1_737_131), .ZN(n_1_737_1239));
   OR2_X1 i_1_737_1240 (.A1(\out_as[4] [3]), .A2(n_1_737_130), .ZN(n_1_737_1240));
   OR2_X1 i_1_737_1241 (.A1(\out_as[3] [3]), .A2(n_1_737_129), .ZN(n_1_737_1241));
   OR2_X1 i_1_737_1242 (.A1(\out_as[2] [3]), .A2(n_1_737_128), .ZN(n_1_737_1242));
   OR2_X1 i_1_737_1243 (.A1(\out_as[1] [3]), .A2(n_1_737_127), .ZN(n_1_737_1243));
   OR2_X1 i_1_737_1244 (.A1(\out_as[0] [3]), .A2(n_1_737_126), .ZN(n_1_737_1244));
   OR2_X1 i_1_737_1245 (.A1(n_1_737_125), .A2(n_1_737_5150), .ZN(n_1_737_1245));
   OR2_X1 i_1_737_1246 (.A1(n_1_737_124), .A2(n_1_737_5162), .ZN(n_1_737_1246));
   OR2_X1 i_1_737_1247 (.A1(n_1_737_123), .A2(n_1_737_5381), .ZN(n_1_737_1247));
   OR2_X1 i_1_737_1248 (.A1(n_1_737_122), .A2(n_1_737_5208), .ZN(n_1_737_1248));
   OR2_X1 i_1_737_1249 (.A1(n_1_737_121), .A2(n_1_737_5269), .ZN(n_1_737_1249));
   OR2_X1 i_1_737_1250 (.A1(n_1_737_120), .A2(n_1_737_5313), .ZN(n_1_737_1250));
   OR2_X1 i_1_737_1251 (.A1(n_1_737_119), .A2(n_1_737_5351), .ZN(n_1_737_1251));
   OR2_X1 i_1_737_1252 (.A1(\out_as[6] [2]), .A2(n_1_737_125), .ZN(n_1_737_1252));
   OR2_X1 i_1_737_1253 (.A1(\out_as[5] [2]), .A2(n_1_737_124), .ZN(n_1_737_1253));
   OR2_X1 i_1_737_1254 (.A1(\out_as[4] [2]), .A2(n_1_737_123), .ZN(n_1_737_1254));
   OR2_X1 i_1_737_1255 (.A1(\out_as[3] [2]), .A2(n_1_737_122), .ZN(n_1_737_1255));
   OR2_X1 i_1_737_1256 (.A1(\out_as[2] [2]), .A2(n_1_737_121), .ZN(n_1_737_1256));
   OR2_X1 i_1_737_1257 (.A1(\out_as[1] [2]), .A2(n_1_737_120), .ZN(n_1_737_1257));
   OR2_X1 i_1_737_1258 (.A1(\out_as[0] [2]), .A2(n_1_737_119), .ZN(n_1_737_1258));
   OR2_X1 i_1_737_1259 (.A1(\out_as[7] [2]), .A2(n_1_737_113), .ZN(n_1_737_1259));
   OR2_X1 i_1_737_1260 (.A1(\out_as[7] [3]), .A2(n_1_737_114), .ZN(n_1_737_1260));
   OR2_X1 i_1_737_1261 (.A1(\out_as[7] [3]), .A2(n_1_737_108), .ZN(n_1_737_1261));
   OR2_X1 i_1_737_1262 (.A1(\out_as[7] [3]), .A2(n_1_737_103), .ZN(n_1_737_1262));
   OR2_X1 i_1_737_1263 (.A1(n_1_737_113), .A2(n_1_737_5145), .ZN(n_1_737_1263));
   OR2_X1 i_1_737_1264 (.A1(\out_as[7] [4]), .A2(n_1_737_115), .ZN(n_1_737_1264));
   OR2_X1 i_1_737_1265 (.A1(\out_as[7] [4]), .A2(n_1_737_109), .ZN(n_1_737_1265));
   OR2_X1 i_1_737_1266 (.A1(\out_as[7] [4]), .A2(n_1_737_104), .ZN(n_1_737_1266));
   OR2_X1 i_1_737_1267 (.A1(\out_as[7] [4]), .A2(n_1_737_99), .ZN(n_1_737_1267));
   OR2_X1 i_1_737_1268 (.A1(\out_as[7] [4]), .A2(n_1_737_95), .ZN(n_1_737_1268));
   OR2_X1 i_1_737_1269 (.A1(\out_as[7] [4]), .A2(n_1_737_91), .ZN(n_1_737_1269));
   OR2_X1 i_1_737_1270 (.A1(\out_as[7] [4]), .A2(n_1_737_87), .ZN(n_1_737_1270));
   OR2_X1 i_1_737_1271 (.A1(n_1_737_114), .A2(n_1_737_5144), .ZN(n_1_737_1271));
   OR2_X1 i_1_737_1272 (.A1(n_1_737_108), .A2(n_1_737_5144), .ZN(n_1_737_1272));
   OR2_X1 i_1_737_1273 (.A1(n_1_737_103), .A2(n_1_737_5144), .ZN(n_1_737_1273));
   OR2_X1 i_1_737_1274 (.A1(n_1_737_113), .A2(n_1_737_5143), .ZN(n_1_737_1274));
   OR2_X1 i_1_737_1275 (.A1(\out_as[7] [5]), .A2(n_1_737_116), .ZN(n_1_737_1275));
   OR2_X1 i_1_737_1276 (.A1(\out_as[7] [5]), .A2(n_1_737_110), .ZN(n_1_737_1276));
   OR2_X1 i_1_737_1277 (.A1(\out_as[7] [5]), .A2(n_1_737_105), .ZN(n_1_737_1277));
   OR2_X1 i_1_737_1278 (.A1(\out_as[7] [5]), .A2(n_1_737_100), .ZN(n_1_737_1278));
   OR2_X1 i_1_737_1279 (.A1(\out_as[7] [5]), .A2(n_1_737_96), .ZN(n_1_737_1279));
   OR2_X1 i_1_737_1280 (.A1(\out_as[7] [5]), .A2(n_1_737_92), .ZN(n_1_737_1280));
   OR2_X1 i_1_737_1281 (.A1(\out_as[7] [5]), .A2(n_1_737_88), .ZN(n_1_737_1281));
   OR2_X1 i_1_737_1282 (.A1(\out_as[7] [5]), .A2(n_1_737_84), .ZN(n_1_737_1282));
   OR2_X1 i_1_737_1283 (.A1(\out_as[7] [5]), .A2(n_1_737_81), .ZN(n_1_737_1283));
   OR2_X1 i_1_737_1284 (.A1(\out_as[7] [5]), .A2(n_1_737_78), .ZN(n_1_737_1284));
   OR2_X1 i_1_737_1285 (.A1(\out_as[7] [5]), .A2(n_1_737_75), .ZN(n_1_737_1285));
   OR2_X1 i_1_737_1286 (.A1(\out_as[7] [5]), .A2(n_1_737_72), .ZN(n_1_737_1286));
   OR2_X1 i_1_737_1287 (.A1(\out_as[7] [5]), .A2(n_1_737_69), .ZN(n_1_737_1287));
   OR2_X1 i_1_737_1288 (.A1(\out_as[7] [5]), .A2(n_1_737_66), .ZN(n_1_737_1288));
   OR2_X1 i_1_737_1289 (.A1(\out_as[7] [5]), .A2(n_1_737_63), .ZN(n_1_737_1289));
   OR2_X1 i_1_737_1290 (.A1(n_1_737_115), .A2(n_1_737_5142), .ZN(n_1_737_1290));
   OR2_X1 i_1_737_1291 (.A1(n_1_737_109), .A2(n_1_737_5142), .ZN(n_1_737_1291));
   OR2_X1 i_1_737_1292 (.A1(n_1_737_104), .A2(n_1_737_5142), .ZN(n_1_737_1292));
   OR2_X1 i_1_737_1293 (.A1(n_1_737_99), .A2(n_1_737_5142), .ZN(n_1_737_1293));
   OR2_X1 i_1_737_1294 (.A1(n_1_737_95), .A2(n_1_737_5142), .ZN(n_1_737_1294));
   OR2_X1 i_1_737_1295 (.A1(n_1_737_91), .A2(n_1_737_5142), .ZN(n_1_737_1295));
   OR2_X1 i_1_737_1296 (.A1(n_1_737_87), .A2(n_1_737_5142), .ZN(n_1_737_1296));
   OR2_X1 i_1_737_1297 (.A1(n_1_737_114), .A2(n_1_737_5138), .ZN(n_1_737_1297));
   OR2_X1 i_1_737_1298 (.A1(n_1_737_108), .A2(n_1_737_5138), .ZN(n_1_737_1298));
   OR2_X1 i_1_737_1299 (.A1(n_1_737_103), .A2(n_1_737_5138), .ZN(n_1_737_1299));
   OR2_X1 i_1_737_1300 (.A1(n_1_737_113), .A2(n_1_737_5141), .ZN(n_1_737_1300));
   OR2_X1 i_1_737_1301 (.A1(\out_as[7] [5]), .A2(n_1_737_1302), .ZN(n_1_737_1301));
   OR2_X1 i_1_737_1302 (.A1(\out_as[7] [4]), .A2(n_1_737_2024), .ZN(n_1_737_1302));
   OAI21_X1 i_1_737_1303 (.A(n_1_737_1303), .B1(n_1_737_5595), .B2(n_1_737_1308), 
      .ZN(n_2));
   OAI211_X1 i_1_737_1304 (.A(n_1_737_1308), .B(n_1_737_1304), .C1(in_data[8]), 
      .C2(n_1_737_1970), .ZN(n_1_737_1303));
   OAI221_X1 i_1_737_1305 (.A(n_1_737_1970), .B1(n_1_737_5597), .B2(n_1_737_1973), 
      .C1(n_1_737_1974), .C2(n_1_737_1305), .ZN(n_1_737_1304));
   AOI22_X1 i_1_737_1306 (.A1(n_1_737_1977), .A2(n_1_737_1306), .B1(in_data[16]), 
      .B2(n_1_737_1978), .ZN(n_1_737_1305));
   OAI21_X1 i_1_737_1307 (.A(n_1_737_1307), .B1(n_1_737_5599), .B2(n_1_737_1975), 
      .ZN(n_1_737_1306));
   OAI221_X1 i_1_737_1308 (.A(n_1_737_1975), .B1(in_data[28]), .B2(n_1_737_1972), 
      .C1(in_data[24]), .C2(n_1_737_1971), .ZN(n_1_737_1307));
   NOR2_X1 i_1_737_1309 (.A1(n_1_737_5594), .A2(n_129), .ZN(n_1_737_1308));
   AOI21_X1 i_1_737_1310 (.A(n_1_737_1309), .B1(n_1_737_5596), .B2(n_1_737_2009), 
      .ZN(n_3));
   AOI211_X1 i_1_737_1311 (.A(n_1_737_1310), .B(n_1_737_2009), .C1(in_data[12]), 
      .C2(n_1_737_1998), .ZN(n_1_737_1309));
   AOI211_X1 i_1_737_1312 (.A(n_1_737_1998), .B(n_1_737_1311), .C1(n_1_737_5598), 
      .C2(n_1_737_2015), .ZN(n_1_737_1310));
   AOI221_X1 i_1_737_1313 (.A(n_1_737_2015), .B1(n_1_737_1986), .B2(n_1_737_1312), 
      .C1(in_data[20]), .C2(n_1_737_1987), .ZN(n_1_737_1311));
   OAI22_X1 i_1_737_1314 (.A1(n_1_737_5600), .A2(n_1_737_1992), .B1(n_1_737_5601), 
      .B2(n_1_737_1993), .ZN(n_1_737_1312));
   AOI21_X1 i_1_737_1315 (.A(n_1_737_1313), .B1(n_1_737_5597), .B2(n_1_737_2087), 
      .ZN(n_4));
   AOI211_X1 i_1_737_1316 (.A(n_1_737_1314), .B(n_1_737_2087), .C1(in_data[16]), 
      .C2(n_1_737_2085), .ZN(n_1_737_1313));
   AOI221_X1 i_1_737_1317 (.A(n_1_737_2085), .B1(n_1_737_2078), .B2(n_1_737_1315), 
      .C1(n_1_737_5599), .C2(n_1_737_2077), .ZN(n_1_737_1314));
   OAI22_X1 i_1_737_1318 (.A1(in_data[24]), .A2(n_1_737_2083), .B1(in_data[28]), 
      .B2(n_1_737_2082), .ZN(n_1_737_1315));
   AOI21_X1 i_1_737_1319 (.A(n_1_737_1316), .B1(n_1_737_5597), .B2(n_1_737_2100), 
      .ZN(n_5));
   AOI221_X1 i_1_737_1320 (.A(n_1_737_2100), .B1(n_1_737_2095), .B2(n_1_737_1317), 
      .C1(in_data[16]), .C2(n_1_737_2094), .ZN(n_1_737_1316));
   AOI21_X1 i_1_737_1321 (.A(n_1_737_1318), .B1(n_1_737_5599), .B2(n_1_737_2097), 
      .ZN(n_1_737_1317));
   AOI221_X1 i_1_737_1322 (.A(n_1_737_2097), .B1(in_data[28]), .B2(n_1_737_2092), 
      .C1(in_data[24]), .C2(n_1_737_2091), .ZN(n_1_737_1318));
   OAI222_X1 i_1_737_1323 (.A1(n_1_737_5597), .A2(n_1_737_2140), .B1(
      n_1_737_2139), .B2(n_1_737_1321), .C1(n_1_737_2136), .C2(n_1_737_1319), 
      .ZN(n_6));
   OAI22_X1 i_1_737_1324 (.A1(n_1_737_2150), .A2(n_1_737_1320), .B1(in_data[20]), 
      .B2(n_1_737_2151), .ZN(n_1_737_1319));
   AOI22_X1 i_1_737_1325 (.A1(n_1_737_5601), .A2(n_1_737_2143), .B1(n_1_737_5600), 
      .B2(n_1_737_2144), .ZN(n_1_737_1320));
   OR2_X1 i_1_737_1326 (.A1(n_1_737_5598), .A2(n_1_737_2137), .ZN(n_1_737_1321));
   AOI22_X1 i_1_737_1327 (.A1(n_1_737_2281), .A2(n_1_737_1322), .B1(n_1_737_5597), 
      .B2(n_1_737_2280), .ZN(n_7));
   OAI22_X1 i_1_737_1328 (.A1(in_data[16]), .A2(n_1_737_2273), .B1(n_1_737_1324), 
      .B2(n_1_737_1323), .ZN(n_1_737_1322));
   OAI21_X1 i_1_737_1329 (.A(n_1_737_2273), .B1(n_1_737_5599), .B2(n_1_737_2276), 
      .ZN(n_1_737_1323));
   AOI21_X1 i_1_737_1330 (.A(n_1_737_1325), .B1(n_1_737_5601), .B2(n_1_737_2269), 
      .ZN(n_1_737_1324));
   OAI21_X1 i_1_737_1331 (.A(n_1_737_2276), .B1(in_data[24]), .B2(n_1_737_2269), 
      .ZN(n_1_737_1325));
   OAI21_X1 i_1_737_1332 (.A(n_1_737_1326), .B1(n_1_737_5597), .B2(n_1_737_2295), 
      .ZN(n_8));
   OAI21_X1 i_1_737_1333 (.A(n_1_737_2295), .B1(n_1_737_1328), .B2(n_1_737_1327), 
      .ZN(n_1_737_1326));
   NOR2_X1 i_1_737_1334 (.A1(n_1_737_5598), .A2(n_1_737_2293), .ZN(n_1_737_1327));
   AOI21_X1 i_1_737_1335 (.A(n_1_737_1329), .B1(n_1_737_2287), .B2(n_1_737_1330), 
      .ZN(n_1_737_1328));
   OAI21_X1 i_1_737_1336 (.A(n_1_737_2293), .B1(in_data[20]), .B2(n_1_737_2287), 
      .ZN(n_1_737_1329));
   AOI22_X1 i_1_737_1337 (.A1(in_data[24]), .A2(n_1_737_2290), .B1(in_data[28]), 
      .B2(n_1_737_2289), .ZN(n_1_737_1330));
   AOI21_X1 i_1_737_1338 (.A(n_1_737_1331), .B1(n_1_737_5597), .B2(n_1_737_2317), 
      .ZN(n_9));
   AOI211_X1 i_1_737_1339 (.A(n_1_737_1332), .B(n_1_737_2317), .C1(in_data[16]), 
      .C2(n_1_737_2300), .ZN(n_1_737_1331));
   AOI211_X1 i_1_737_1340 (.A(n_1_737_1333), .B(n_1_737_2300), .C1(n_1_737_5599), 
      .C2(n_1_737_2304), .ZN(n_1_737_1332));
   AOI221_X1 i_1_737_1341 (.A(n_1_737_2304), .B1(in_data[28]), .B2(n_1_737_2310), 
      .C1(in_data[24]), .C2(n_1_737_2309), .ZN(n_1_737_1333));
   AOI21_X1 i_1_737_1342 (.A(n_1_737_1334), .B1(n_1_737_5597), .B2(n_1_737_2349), 
      .ZN(n_10));
   AOI211_X1 i_1_737_1343 (.A(n_1_737_1335), .B(n_1_737_2349), .C1(in_data[16]), 
      .C2(n_1_737_2346), .ZN(n_1_737_1334));
   AOI221_X1 i_1_737_1344 (.A(n_1_737_2346), .B1(n_1_737_2339), .B2(n_1_737_1336), 
      .C1(n_1_737_5599), .C2(n_1_737_2338), .ZN(n_1_737_1335));
   OAI22_X1 i_1_737_1345 (.A1(in_data[24]), .A2(n_1_737_2344), .B1(in_data[28]), 
      .B2(n_1_737_2343), .ZN(n_1_737_1336));
   OAI21_X1 i_1_737_1346 (.A(n_1_737_1337), .B1(n_1_737_5596), .B2(n_1_737_2391), 
      .ZN(n_11));
   OAI221_X1 i_1_737_1347 (.A(n_1_737_2391), .B1(n_1_737_2386), .B2(n_1_737_1338), 
      .C1(in_data[12]), .C2(n_1_737_2385), .ZN(n_1_737_1337));
   AOI21_X1 i_1_737_1348 (.A(n_1_737_1339), .B1(n_1_737_5598), .B2(n_1_737_2394), 
      .ZN(n_1_737_1338));
   AOI211_X1 i_1_737_1349 (.A(n_1_737_1340), .B(n_1_737_2394), .C1(in_data[20]), 
      .C2(n_1_737_2396), .ZN(n_1_737_1339));
   AOI221_X1 i_1_737_1350 (.A(n_1_737_2396), .B1(n_1_737_5600), .B2(n_1_737_2389), 
      .C1(n_1_737_5601), .C2(n_1_737_2388), .ZN(n_1_737_1340));
   AOI21_X1 i_1_737_1351 (.A(n_1_737_1341), .B1(n_1_737_5597), .B2(n_1_737_2466), 
      .ZN(n_12));
   AOI221_X1 i_1_737_1352 (.A(n_1_737_2466), .B1(n_1_737_2464), .B2(n_1_737_1342), 
      .C1(in_data[16]), .C2(n_1_737_2463), .ZN(n_1_737_1341));
   AOI21_X1 i_1_737_1353 (.A(n_1_737_1343), .B1(n_1_737_5599), .B2(n_1_737_2455), 
      .ZN(n_1_737_1342));
   AOI221_X1 i_1_737_1354 (.A(n_1_737_2455), .B1(in_data[28]), .B2(n_1_737_2461), 
      .C1(in_data[24]), .C2(n_1_737_2460), .ZN(n_1_737_1343));
   AOI21_X1 i_1_737_1355 (.A(n_1_737_1344), .B1(n_1_737_5597), .B2(n_1_737_2498), 
      .ZN(n_13));
   AOI221_X1 i_1_737_1356 (.A(n_1_737_2498), .B1(n_1_737_2493), .B2(n_1_737_1345), 
      .C1(in_data[16]), .C2(n_1_737_2492), .ZN(n_1_737_1344));
   AOI21_X1 i_1_737_1357 (.A(n_1_737_1346), .B1(n_1_737_5599), .B2(n_1_737_2495), 
      .ZN(n_1_737_1345));
   AOI221_X1 i_1_737_1358 (.A(n_1_737_2495), .B1(in_data[28]), .B2(n_1_737_2490), 
      .C1(in_data[24]), .C2(n_1_737_2489), .ZN(n_1_737_1346));
   OAI21_X1 i_1_737_1359 (.A(n_1_737_1347), .B1(n_1_737_5596), .B2(n_1_737_2524), 
      .ZN(n_14));
   OAI221_X1 i_1_737_1360 (.A(n_1_737_2524), .B1(in_data[12]), .B2(n_1_737_2531), 
      .C1(n_1_737_2532), .C2(n_1_737_1348), .ZN(n_1_737_1347));
   OAI21_X1 i_1_737_1361 (.A(n_1_737_1349), .B1(n_1_737_5598), .B2(n_1_737_2522), 
      .ZN(n_1_737_1348));
   OAI21_X1 i_1_737_1362 (.A(n_1_737_2522), .B1(n_1_737_1351), .B2(n_1_737_1350), 
      .ZN(n_1_737_1349));
   NOR2_X1 i_1_737_1363 (.A1(n_1_737_5599), .A2(n_1_737_2528), .ZN(n_1_737_1350));
   AOI21_X1 i_1_737_1364 (.A(n_1_737_1352), .B1(n_1_737_5600), .B2(n_1_737_2526), 
      .ZN(n_1_737_1351));
   OAI21_X1 i_1_737_1365 (.A(n_1_737_2528), .B1(in_data[28]), .B2(n_1_737_2526), 
      .ZN(n_1_737_1352));
   AOI21_X1 i_1_737_1366 (.A(n_1_737_1353), .B1(n_1_737_5597), .B2(n_1_737_2550), 
      .ZN(n_15));
   AOI221_X1 i_1_737_1367 (.A(n_1_737_2550), .B1(n_1_737_2538), .B2(n_1_737_1354), 
      .C1(in_data[16]), .C2(n_1_737_2537), .ZN(n_1_737_1353));
   AOI21_X1 i_1_737_1368 (.A(n_1_737_1355), .B1(n_1_737_5599), .B2(n_1_737_2540), 
      .ZN(n_1_737_1354));
   AOI221_X1 i_1_737_1369 (.A(n_1_737_2540), .B1(in_data[28]), .B2(n_1_737_2545), 
      .C1(in_data[24]), .C2(n_1_737_2544), .ZN(n_1_737_1355));
   AOI21_X1 i_1_737_1370 (.A(n_1_737_1356), .B1(n_1_737_5597), .B2(n_1_737_2587), 
      .ZN(n_16));
   AOI211_X1 i_1_737_1371 (.A(n_1_737_1357), .B(n_1_737_2587), .C1(in_data[16]), 
      .C2(n_1_737_2574), .ZN(n_1_737_1356));
   AOI221_X1 i_1_737_1372 (.A(n_1_737_2574), .B1(n_1_737_2578), .B2(n_1_737_1358), 
      .C1(n_1_737_5599), .C2(n_1_737_2577), .ZN(n_1_737_1357));
   OAI22_X1 i_1_737_1373 (.A1(in_data[24]), .A2(n_1_737_2582), .B1(in_data[28]), 
      .B2(n_1_737_2581), .ZN(n_1_737_1358));
   AOI21_X1 i_1_737_1374 (.A(n_1_737_1359), .B1(n_1_737_5597), .B2(n_1_737_2615), 
      .ZN(n_17));
   AOI211_X1 i_1_737_1375 (.A(n_1_737_2615), .B(n_1_737_1360), .C1(in_data[16]), 
      .C2(n_1_737_2626), .ZN(n_1_737_1359));
   AOI211_X1 i_1_737_1376 (.A(n_1_737_2626), .B(n_1_737_1361), .C1(n_1_737_5599), 
      .C2(n_1_737_2623), .ZN(n_1_737_1360));
   AOI221_X1 i_1_737_1377 (.A(n_1_737_2623), .B1(in_data[24]), .B2(n_1_737_2620), 
      .C1(in_data[28]), .C2(n_1_737_2619), .ZN(n_1_737_1361));
   AOI21_X1 i_1_737_1378 (.A(n_1_737_1362), .B1(n_1_737_5597), .B2(n_1_737_2644), 
      .ZN(n_18));
   AOI221_X1 i_1_737_1379 (.A(n_1_737_2644), .B1(n_1_737_2641), .B2(n_1_737_1363), 
      .C1(in_data[16]), .C2(n_1_737_2640), .ZN(n_1_737_1362));
   AOI21_X1 i_1_737_1380 (.A(n_1_737_1364), .B1(n_1_737_5599), .B2(n_1_737_2632), 
      .ZN(n_1_737_1363));
   AOI221_X1 i_1_737_1381 (.A(n_1_737_2632), .B1(in_data[28]), .B2(n_1_737_2638), 
      .C1(in_data[24]), .C2(n_1_737_2637), .ZN(n_1_737_1364));
   OAI21_X1 i_1_737_1382 (.A(n_1_737_1365), .B1(n_1_737_5597), .B2(n_1_737_2896), 
      .ZN(n_19));
   OAI211_X1 i_1_737_1383 (.A(n_1_737_2896), .B(n_1_737_1366), .C1(in_data[16]), 
      .C2(n_1_737_2894), .ZN(n_1_737_1365));
   OAI221_X1 i_1_737_1384 (.A(n_1_737_2894), .B1(n_1_737_5599), .B2(n_1_737_2898), 
      .C1(n_1_737_1368), .C2(n_1_737_1367), .ZN(n_1_737_1366));
   OAI21_X1 i_1_737_1385 (.A(n_1_737_2898), .B1(in_data[24]), .B2(n_1_737_2892), 
      .ZN(n_1_737_1367));
   NOR2_X1 i_1_737_1386 (.A1(in_data[28]), .A2(n_1_737_2891), .ZN(n_1_737_1368));
   AOI21_X1 i_1_737_1387 (.A(n_1_737_1369), .B1(n_1_737_5597), .B2(n_1_737_3056), 
      .ZN(n_20));
   AOI211_X1 i_1_737_1388 (.A(n_1_737_1370), .B(n_1_737_3056), .C1(in_data[16]), 
      .C2(n_1_737_3053), .ZN(n_1_737_1369));
   AOI221_X1 i_1_737_1389 (.A(n_1_737_3053), .B1(n_1_737_3046), .B2(n_1_737_1371), 
      .C1(n_1_737_5599), .C2(n_1_737_3045), .ZN(n_1_737_1370));
   OAI22_X1 i_1_737_1390 (.A1(in_data[24]), .A2(n_1_737_3051), .B1(in_data[28]), 
      .B2(n_1_737_3050), .ZN(n_1_737_1371));
   AOI21_X1 i_1_737_1391 (.A(n_1_737_1372), .B1(n_1_737_5597), .B2(n_1_737_3133), 
      .ZN(n_21));
   AOI211_X1 i_1_737_1392 (.A(n_1_737_3133), .B(n_1_737_1373), .C1(in_data[16]), 
      .C2(n_1_737_3139), .ZN(n_1_737_1372));
   AOI211_X1 i_1_737_1393 (.A(n_1_737_1374), .B(n_1_737_3139), .C1(n_1_737_5599), 
      .C2(n_1_737_3141), .ZN(n_1_737_1373));
   AOI221_X1 i_1_737_1394 (.A(n_1_737_3141), .B1(in_data[28]), .B2(n_1_737_3136), 
      .C1(in_data[24]), .C2(n_1_737_3137), .ZN(n_1_737_1374));
   AOI22_X1 i_1_737_1395 (.A1(n_1_737_3165), .A2(n_1_737_1375), .B1(n_1_737_5597), 
      .B2(n_1_737_3164), .ZN(n_22));
   OAI21_X1 i_1_737_1396 (.A(n_1_737_1376), .B1(in_data[16]), .B2(n_1_737_3147), 
      .ZN(n_1_737_1375));
   OAI211_X1 i_1_737_1397 (.A(n_1_737_3147), .B(n_1_737_1377), .C1(n_1_737_5599), 
      .C2(n_1_737_3156), .ZN(n_1_737_1376));
   OAI221_X1 i_1_737_1398 (.A(n_1_737_3156), .B1(in_data[28]), .B2(n_1_737_3152), 
      .C1(in_data[24]), .C2(n_1_737_3151), .ZN(n_1_737_1377));
   AOI21_X1 i_1_737_1399 (.A(n_1_737_1378), .B1(n_1_737_5597), .B2(n_1_737_3576), 
      .ZN(n_23));
   NOR2_X1 i_1_737_1400 (.A1(n_1_737_3576), .A2(n_1_737_1379), .ZN(n_1_737_1378));
   OAI21_X1 i_1_737_1401 (.A(n_1_737_1380), .B1(n_1_737_5598), .B2(n_1_737_3583), 
      .ZN(n_1_737_1379));
   OAI211_X1 i_1_737_1402 (.A(n_1_737_1381), .B(n_1_737_3583), .C1(in_data[20]), 
      .C2(n_1_737_3580), .ZN(n_1_737_1380));
   OAI221_X1 i_1_737_1403 (.A(n_1_737_3580), .B1(n_1_737_5601), .B2(n_1_737_3586), 
      .C1(n_1_737_5600), .C2(n_1_737_3587), .ZN(n_1_737_1381));
   AOI22_X1 i_1_737_1404 (.A1(n_1_737_3612), .A2(n_1_737_1382), .B1(n_1_737_5597), 
      .B2(n_1_737_3611), .ZN(n_24));
   OAI21_X1 i_1_737_1405 (.A(n_1_737_1383), .B1(in_data[16]), .B2(n_1_737_3599), 
      .ZN(n_1_737_1382));
   OAI211_X1 i_1_737_1406 (.A(n_1_737_3599), .B(n_1_737_1384), .C1(n_1_737_5599), 
      .C2(n_1_737_3603), .ZN(n_1_737_1383));
   OAI221_X1 i_1_737_1407 (.A(n_1_737_3603), .B1(in_data[24]), .B2(n_1_737_3593), 
      .C1(in_data[28]), .C2(n_1_737_3594), .ZN(n_1_737_1384));
   AOI22_X1 i_1_737_1408 (.A1(n_1_737_3637), .A2(n_1_737_1385), .B1(n_1_737_5597), 
      .B2(n_1_737_3636), .ZN(n_25));
   OAI21_X1 i_1_737_1409 (.A(n_1_737_1386), .B1(in_data[16]), .B2(n_1_737_3624), 
      .ZN(n_1_737_1385));
   OAI211_X1 i_1_737_1410 (.A(n_1_737_3624), .B(n_1_737_1387), .C1(n_1_737_5599), 
      .C2(n_1_737_3632), .ZN(n_1_737_1386));
   OAI221_X1 i_1_737_1411 (.A(n_1_737_3632), .B1(in_data[24]), .B2(n_1_737_3618), 
      .C1(in_data[28]), .C2(n_1_737_3619), .ZN(n_1_737_1387));
   AOI22_X1 i_1_737_1412 (.A1(n_1_737_3662), .A2(n_1_737_1388), .B1(n_1_737_5597), 
      .B2(n_1_737_3663), .ZN(n_26));
   OAI21_X1 i_1_737_1413 (.A(n_1_737_1389), .B1(in_data[16]), .B2(n_1_737_3647), 
      .ZN(n_1_737_1388));
   OAI211_X1 i_1_737_1414 (.A(n_1_737_3647), .B(n_1_737_1390), .C1(n_1_737_5599), 
      .C2(n_1_737_3657), .ZN(n_1_737_1389));
   OAI221_X1 i_1_737_1415 (.A(n_1_737_3657), .B1(in_data[24]), .B2(n_1_737_3651), 
      .C1(in_data[28]), .C2(n_1_737_3652), .ZN(n_1_737_1390));
   AOI22_X1 i_1_737_1416 (.A1(n_1_737_3690), .A2(n_1_737_1391), .B1(n_1_737_5597), 
      .B2(n_1_737_3689), .ZN(n_27));
   OAI21_X1 i_1_737_1417 (.A(n_1_737_1392), .B1(in_data[16]), .B2(n_1_737_3677), 
      .ZN(n_1_737_1391));
   OAI211_X1 i_1_737_1418 (.A(n_1_737_3677), .B(n_1_737_1393), .C1(n_1_737_5599), 
      .C2(n_1_737_3681), .ZN(n_1_737_1392));
   OAI221_X1 i_1_737_1419 (.A(n_1_737_3681), .B1(in_data[24]), .B2(n_1_737_3671), 
      .C1(in_data[28]), .C2(n_1_737_3672), .ZN(n_1_737_1393));
   AOI22_X1 i_1_737_1420 (.A1(n_1_737_3817), .A2(n_1_737_1394), .B1(n_1_737_5597), 
      .B2(n_1_737_3816), .ZN(n_28));
   OAI21_X1 i_1_737_1421 (.A(n_1_737_1395), .B1(in_data[16]), .B2(n_1_737_3813), 
      .ZN(n_1_737_1394));
   OAI211_X1 i_1_737_1422 (.A(n_1_737_3813), .B(n_1_737_1396), .C1(n_1_737_5599), 
      .C2(n_1_737_3822), .ZN(n_1_737_1395));
   OAI221_X1 i_1_737_1423 (.A(n_1_737_3822), .B1(in_data[28]), .B2(n_1_737_3825), 
      .C1(in_data[24]), .C2(n_1_737_3826), .ZN(n_1_737_1396));
   AOI21_X1 i_1_737_1424 (.A(n_1_737_1397), .B1(n_1_737_5597), .B2(n_1_737_3910), 
      .ZN(n_29));
   AOI211_X1 i_1_737_1425 (.A(n_1_737_1398), .B(n_1_737_3910), .C1(in_data[16]), 
      .C2(n_1_737_3891), .ZN(n_1_737_1397));
   AOI211_X1 i_1_737_1426 (.A(n_1_737_1399), .B(n_1_737_3891), .C1(n_1_737_5599), 
      .C2(n_1_737_3904), .ZN(n_1_737_1398));
   AOI221_X1 i_1_737_1427 (.A(n_1_737_3904), .B1(in_data[28]), .B2(n_1_737_3897), 
      .C1(in_data[24]), .C2(n_1_737_3898), .ZN(n_1_737_1399));
   AOI22_X1 i_1_737_1428 (.A1(n_1_737_4179), .A2(n_1_737_1400), .B1(n_1_737_5597), 
      .B2(n_1_737_4180), .ZN(n_30));
   OAI21_X1 i_1_737_1429 (.A(n_1_737_1401), .B1(in_data[16]), .B2(n_1_737_4160), 
      .ZN(n_1_737_1400));
   OAI211_X1 i_1_737_1430 (.A(n_1_737_4160), .B(n_1_737_1402), .C1(n_1_737_5599), 
      .C2(n_1_737_4173), .ZN(n_1_737_1401));
   OAI221_X1 i_1_737_1431 (.A(n_1_737_4173), .B1(in_data[24]), .B2(n_1_737_4166), 
      .C1(in_data[28]), .C2(n_1_737_4167), .ZN(n_1_737_1402));
   OAI21_X1 i_1_737_1432 (.A(n_1_737_1403), .B1(n_1_737_5597), .B2(n_1_737_4202), 
      .ZN(n_31));
   NAND2_X1 i_1_737_1433 (.A1(n_1_737_4202), .A2(n_1_737_1404), .ZN(n_1_737_1403));
   AOI21_X1 i_1_737_1434 (.A(n_1_737_1405), .B1(n_1_737_5598), .B2(n_1_737_4191), 
      .ZN(n_1_737_1404));
   AOI221_X1 i_1_737_1435 (.A(n_1_737_4191), .B1(n_1_737_4196), .B2(n_1_737_1406), 
      .C1(in_data[20]), .C2(n_1_737_4195), .ZN(n_1_737_1405));
   AOI22_X1 i_1_737_1436 (.A1(n_1_737_5601), .A2(n_1_737_4187), .B1(n_1_737_5600), 
      .B2(n_1_737_4186), .ZN(n_1_737_1406));
   AOI22_X1 i_1_737_1437 (.A1(n_1_737_4281), .A2(n_1_737_1407), .B1(n_1_737_5597), 
      .B2(n_1_737_4280), .ZN(n_32));
   OAI21_X1 i_1_737_1438 (.A(n_1_737_1408), .B1(in_data[16]), .B2(n_1_737_4259), 
      .ZN(n_1_737_1407));
   OAI211_X1 i_1_737_1439 (.A(n_1_737_4259), .B(n_1_737_1409), .C1(n_1_737_5599), 
      .C2(n_1_737_4274), .ZN(n_1_737_1408));
   OAI221_X1 i_1_737_1440 (.A(n_1_737_4274), .B1(in_data[28]), .B2(n_1_737_4268), 
      .C1(in_data[24]), .C2(n_1_737_4267), .ZN(n_1_737_1409));
   AOI22_X1 i_1_737_1441 (.A1(n_1_737_4321), .A2(n_1_737_1410), .B1(n_1_737_5597), 
      .B2(n_1_737_4320), .ZN(n_33));
   OAI21_X1 i_1_737_1442 (.A(n_1_737_1411), .B1(in_data[16]), .B2(n_1_737_4327), 
      .ZN(n_1_737_1410));
   OAI221_X1 i_1_737_1443 (.A(n_1_737_4327), .B1(n_1_737_1413), .B2(n_1_737_1412), 
      .C1(n_1_737_5599), .C2(n_1_737_4324), .ZN(n_1_737_1411));
   OAI21_X1 i_1_737_1444 (.A(n_1_737_4324), .B1(in_data[28]), .B2(n_1_737_4330), 
      .ZN(n_1_737_1412));
   AND2_X1 i_1_737_1445 (.A1(n_1_737_5600), .A2(n_1_737_4330), .ZN(n_1_737_1413));
   AOI22_X1 i_1_737_1446 (.A1(n_1_737_4589), .A2(n_1_737_1414), .B1(n_1_737_5597), 
      .B2(n_1_737_4590), .ZN(n_34));
   OAI21_X1 i_1_737_1447 (.A(n_1_737_1415), .B1(in_data[16]), .B2(n_1_737_4572), 
      .ZN(n_1_737_1414));
   OAI211_X1 i_1_737_1448 (.A(n_1_737_4572), .B(n_1_737_1416), .C1(n_1_737_5599), 
      .C2(n_1_737_4584), .ZN(n_1_737_1415));
   OAI221_X1 i_1_737_1449 (.A(n_1_737_4584), .B1(in_data[24]), .B2(n_1_737_4578), 
      .C1(in_data[28]), .C2(n_1_737_4579), .ZN(n_1_737_1416));
   OAI21_X1 i_1_737_1450 (.A(n_1_737_1417), .B1(n_1_737_5597), .B2(n_1_737_4601), 
      .ZN(n_35));
   OAI21_X1 i_1_737_1451 (.A(n_1_737_4601), .B1(n_1_737_1419), .B2(n_1_737_1418), 
      .ZN(n_1_737_1417));
   NOR2_X1 i_1_737_1452 (.A1(n_1_737_5598), .A2(n_1_737_4598), .ZN(n_1_737_1418));
   AOI21_X1 i_1_737_1453 (.A(n_1_737_1420), .B1(n_1_737_5599), .B2(n_1_737_4605), 
      .ZN(n_1_737_1419));
   OAI21_X1 i_1_737_1454 (.A(n_1_737_4598), .B1(n_1_737_4605), .B2(n_1_737_1421), 
      .ZN(n_1_737_1420));
   OAI22_X1 i_1_737_1455 (.A1(n_1_737_5601), .A2(n_1_737_4609), .B1(n_1_737_5600), 
      .B2(n_1_737_4610), .ZN(n_1_737_1421));
   AOI22_X1 i_1_737_1456 (.A1(n_1_737_4672), .A2(n_1_737_1422), .B1(n_1_737_5597), 
      .B2(n_1_737_4671), .ZN(n_36));
   OAI21_X1 i_1_737_1457 (.A(n_1_737_1423), .B1(in_data[16]), .B2(n_1_737_4654), 
      .ZN(n_1_737_1422));
   OAI211_X1 i_1_737_1458 (.A(n_1_737_4654), .B(n_1_737_1424), .C1(n_1_737_5599), 
      .C2(n_1_737_4660), .ZN(n_1_737_1423));
   OAI221_X1 i_1_737_1459 (.A(n_1_737_4660), .B1(in_data[28]), .B2(n_1_737_4649), 
      .C1(in_data[24]), .C2(n_1_737_4648), .ZN(n_1_737_1424));
   OAI21_X1 i_1_737_1460 (.A(n_1_737_1425), .B1(n_1_737_5596), .B2(n_1_737_1431), 
      .ZN(n_37));
   NAND2_X1 i_1_737_1461 (.A1(n_1_737_1431), .A2(n_1_737_1426), .ZN(n_1_737_1425));
   AOI21_X1 i_1_737_1462 (.A(n_1_737_1427), .B1(n_1_737_5597), .B2(n_1_737_2037), 
      .ZN(n_1_737_1426));
   AOI211_X1 i_1_737_1463 (.A(n_1_737_1428), .B(n_1_737_2037), .C1(in_data[16]), 
      .C2(n_1_737_2031), .ZN(n_1_737_1427));
   NOR2_X1 i_1_737_1464 (.A1(n_1_737_2031), .A2(n_1_737_1429), .ZN(n_1_737_1428));
   AOI22_X1 i_1_737_1465 (.A1(n_1_737_2035), .A2(n_1_737_1430), .B1(in_data[20]), 
      .B2(n_1_737_2034), .ZN(n_1_737_1429));
   OAI22_X1 i_1_737_1466 (.A1(n_1_737_5600), .A2(n_1_737_2029), .B1(n_1_737_5601), 
      .B2(n_1_737_2028), .ZN(n_1_737_1430));
   OAI21_X1 i_1_737_1467 (.A(n_136), .B1(n_1_737_5602), .B2(n_135), .ZN(
      n_1_737_1431));
   OAI21_X1 i_1_737_1468 (.A(n_1_737_1432), .B1(n_1_737_5596), .B2(n_1_737_1437), 
      .ZN(n_38));
   OAI211_X1 i_1_737_1469 (.A(n_1_737_1433), .B(n_1_737_1437), .C1(in_data[12]), 
      .C2(n_1_737_2055), .ZN(n_1_737_1432));
   NAND2_X1 i_1_737_1470 (.A1(n_1_737_2055), .A2(n_1_737_1434), .ZN(n_1_737_1433));
   AOI21_X1 i_1_737_1471 (.A(n_1_737_1435), .B1(in_data[16]), .B2(n_1_737_2052), 
      .ZN(n_1_737_1434));
   AOI221_X1 i_1_737_1472 (.A(n_1_737_2052), .B1(n_1_737_5599), .B2(n_1_737_2044), 
      .C1(n_1_737_2045), .C2(n_1_737_1436), .ZN(n_1_737_1435));
   AOI22_X1 i_1_737_1473 (.A1(in_data[28]), .A2(n_1_737_2050), .B1(in_data[24]), 
      .B2(n_1_737_2049), .ZN(n_1_737_1436));
   OAI21_X1 i_1_737_1474 (.A(n_140), .B1(n_1_737_5602), .B2(n_139), .ZN(
      n_1_737_1437));
   INV_X1 i_1_737_1475 (.A(n_1_737_1438), .ZN(n_39));
   OAI21_X1 i_1_737_1476 (.A(n_1_737_1439), .B1(in_data[8]), .B2(n_1_737_1440), 
      .ZN(n_1_737_1438));
   OAI221_X1 i_1_737_1477 (.A(n_1_737_1440), .B1(n_1_737_5597), .B2(n_1_737_2070), 
      .C1(n_1_737_2069), .C2(n_1_737_1441), .ZN(n_1_737_1439));
   OAI21_X1 i_1_737_1478 (.A(n_145), .B1(n_1_737_5602), .B2(n_144), .ZN(
      n_1_737_1440));
   AOI21_X1 i_1_737_1479 (.A(n_1_737_1442), .B1(in_data[16]), .B2(n_1_737_2063), 
      .ZN(n_1_737_1441));
   AOI211_X1 i_1_737_1480 (.A(n_1_737_1443), .B(n_1_737_2063), .C1(n_1_737_5599), 
      .C2(n_1_737_2066), .ZN(n_1_737_1442));
   AOI221_X1 i_1_737_1481 (.A(n_1_737_2066), .B1(in_data[28]), .B2(n_1_737_2061), 
      .C1(in_data[24]), .C2(n_1_737_2060), .ZN(n_1_737_1443));
   OAI22_X1 i_1_737_1482 (.A1(n_1_737_5596), .A2(n_1_737_1447), .B1(n_1_737_1446), 
      .B2(n_1_737_1444), .ZN(n_40));
   OAI21_X1 i_1_737_1483 (.A(n_1_737_1447), .B1(n_1_737_1448), .B2(n_1_737_1445), 
      .ZN(n_1_737_1444));
   OAI21_X1 i_1_737_1484 (.A(n_1_737_2116), .B1(n_1_737_5598), .B2(n_1_737_2114), 
      .ZN(n_1_737_1445));
   NOR2_X1 i_1_737_1485 (.A1(in_data[12]), .A2(n_1_737_2116), .ZN(n_1_737_1446));
   OAI21_X1 i_1_737_1486 (.A(n_156), .B1(n_1_737_5602), .B2(n_155), .ZN(
      n_1_737_1447));
   AOI21_X1 i_1_737_1487 (.A(n_1_737_1449), .B1(n_1_737_2109), .B2(n_1_737_1450), 
      .ZN(n_1_737_1448));
   OAI21_X1 i_1_737_1488 (.A(n_1_737_2114), .B1(in_data[20]), .B2(n_1_737_2109), 
      .ZN(n_1_737_1449));
   AOI22_X1 i_1_737_1489 (.A1(in_data[28]), .A2(n_1_737_2112), .B1(in_data[24]), 
      .B2(n_1_737_2111), .ZN(n_1_737_1450));
   OAI21_X1 i_1_737_1490 (.A(n_1_737_1451), .B1(n_1_737_5596), .B2(n_1_737_2121), 
      .ZN(n_41));
   OAI221_X1 i_1_737_1491 (.A(n_1_737_2121), .B1(in_data[12]), .B2(n_1_737_2126), 
      .C1(n_1_737_2125), .C2(n_1_737_1452), .ZN(n_1_737_1451));
   AOI21_X1 i_1_737_1492 (.A(n_1_737_1453), .B1(n_1_737_5598), .B2(n_1_737_2130), 
      .ZN(n_1_737_1452));
   AOI211_X1 i_1_737_1493 (.A(n_1_737_1454), .B(n_1_737_2130), .C1(in_data[20]), 
      .C2(n_1_737_2123), .ZN(n_1_737_1453));
   AOI221_X1 i_1_737_1494 (.A(n_1_737_2123), .B1(n_1_737_5600), .B2(n_1_737_2132), 
      .C1(n_1_737_5601), .C2(n_1_737_2133), .ZN(n_1_737_1454));
   AOI22_X1 i_1_737_1495 (.A1(n_1_737_5596), .A2(n_1_737_1459), .B1(n_1_737_1460), 
      .B2(n_1_737_1455), .ZN(n_42));
   OAI21_X1 i_1_737_1496 (.A(n_1_737_1456), .B1(in_data[12]), .B2(n_1_737_2167), 
      .ZN(n_1_737_1455));
   OAI221_X1 i_1_737_1497 (.A(n_1_737_2167), .B1(n_1_737_2156), .B2(n_1_737_1457), 
      .C1(n_1_737_5598), .C2(n_1_737_2157), .ZN(n_1_737_1456));
   AOI21_X1 i_1_737_1498 (.A(n_1_737_1458), .B1(in_data[20]), .B2(n_1_737_2159), 
      .ZN(n_1_737_1457));
   AOI221_X1 i_1_737_1499 (.A(n_1_737_2159), .B1(n_1_737_5600), .B2(n_1_737_2164), 
      .C1(n_1_737_5601), .C2(n_1_737_2165), .ZN(n_1_737_1458));
   INV_X1 i_1_737_1500 (.A(n_1_737_1460), .ZN(n_1_737_1459));
   OAI21_X1 i_1_737_1501 (.A(n_167), .B1(n_1_737_5602), .B2(n_166), .ZN(
      n_1_737_1460));
   INV_X1 i_1_737_1502 (.A(n_1_737_1461), .ZN(n_43));
   OAI21_X1 i_1_737_1503 (.A(n_1_737_1462), .B1(in_data[8]), .B2(n_1_737_1466), 
      .ZN(n_1_737_1461));
   OAI211_X1 i_1_737_1504 (.A(n_1_737_1463), .B(n_1_737_1466), .C1(n_1_737_5597), 
      .C2(n_1_737_2186), .ZN(n_1_737_1462));
   OAI221_X1 i_1_737_1505 (.A(n_1_737_2186), .B1(n_1_737_2178), .B2(n_1_737_1464), 
      .C1(in_data[16]), .C2(n_1_737_2179), .ZN(n_1_737_1463));
   OAI21_X1 i_1_737_1506 (.A(n_1_737_1465), .B1(n_1_737_5599), .B2(n_1_737_2182), 
      .ZN(n_1_737_1464));
   OAI221_X1 i_1_737_1507 (.A(n_1_737_2182), .B1(in_data[24]), .B2(n_1_737_2174), 
      .C1(in_data[28]), .C2(n_1_737_2173), .ZN(n_1_737_1465));
   OAI21_X1 i_1_737_1508 (.A(n_172), .B1(n_1_737_5602), .B2(n_171), .ZN(
      n_1_737_1466));
   OAI21_X1 i_1_737_1509 (.A(n_1_737_1467), .B1(n_1_737_5596), .B2(n_1_737_1472), 
      .ZN(n_44));
   OAI211_X1 i_1_737_1510 (.A(n_1_737_1468), .B(n_1_737_1472), .C1(in_data[12]), 
      .C2(n_1_737_2201), .ZN(n_1_737_1467));
   OAI211_X1 i_1_737_1511 (.A(n_1_737_1469), .B(n_1_737_2201), .C1(n_1_737_5598), 
      .C2(n_1_737_2196), .ZN(n_1_737_1468));
   NAND2_X1 i_1_737_1512 (.A1(n_1_737_2196), .A2(n_1_737_1470), .ZN(n_1_737_1469));
   OAI21_X1 i_1_737_1513 (.A(n_1_737_1471), .B1(n_1_737_5599), .B2(n_1_737_2199), 
      .ZN(n_1_737_1470));
   OAI221_X1 i_1_737_1514 (.A(n_1_737_2199), .B1(in_data[28]), .B2(n_1_737_2193), 
      .C1(in_data[24]), .C2(n_1_737_2194), .ZN(n_1_737_1471));
   OAI21_X1 i_1_737_1515 (.A(n_177), .B1(n_1_737_5602), .B2(n_176), .ZN(
      n_1_737_1472));
   AOI22_X1 i_1_737_1516 (.A1(n_1_737_5596), .A2(n_1_737_1477), .B1(n_1_737_1478), 
      .B2(n_1_737_1473), .ZN(n_45));
   OAI21_X1 i_1_737_1517 (.A(n_1_737_1474), .B1(in_data[12]), .B2(n_1_737_2216), 
      .ZN(n_1_737_1473));
   OAI221_X1 i_1_737_1518 (.A(n_1_737_2216), .B1(n_1_737_2211), .B2(n_1_737_1475), 
      .C1(n_1_737_5598), .C2(n_1_737_2212), .ZN(n_1_737_1474));
   AOI21_X1 i_1_737_1519 (.A(n_1_737_1476), .B1(in_data[20]), .B2(n_1_737_2214), 
      .ZN(n_1_737_1475));
   AOI221_X1 i_1_737_1520 (.A(n_1_737_2214), .B1(n_1_737_5601), .B2(n_1_737_2209), 
      .C1(n_1_737_5600), .C2(n_1_737_2208), .ZN(n_1_737_1476));
   INV_X1 i_1_737_1521 (.A(n_1_737_1478), .ZN(n_1_737_1477));
   OAI21_X1 i_1_737_1522 (.A(n_182), .B1(n_1_737_5602), .B2(n_181), .ZN(
      n_1_737_1478));
   OAI22_X1 i_1_737_1523 (.A1(n_1_737_1480), .A2(n_1_737_1479), .B1(n_1_737_5596), 
      .B2(n_1_737_1483), .ZN(n_46));
   OAI21_X1 i_1_737_1524 (.A(n_1_737_1483), .B1(in_data[12]), .B2(n_1_737_2235), 
      .ZN(n_1_737_1479));
   AOI221_X1 i_1_737_1525 (.A(n_1_737_2234), .B1(n_1_737_2225), .B2(n_1_737_1481), 
      .C1(in_data[16]), .C2(n_1_737_2224), .ZN(n_1_737_1480));
   AOI22_X1 i_1_737_1526 (.A1(n_1_737_2228), .A2(n_1_737_1482), .B1(n_1_737_5599), 
      .B2(n_1_737_2227), .ZN(n_1_737_1481));
   OAI22_X1 i_1_737_1527 (.A1(in_data[24]), .A2(n_1_737_2231), .B1(in_data[28]), 
      .B2(n_1_737_2230), .ZN(n_1_737_1482));
   OAI21_X1 i_1_737_1528 (.A(n_187), .B1(n_1_737_5602), .B2(n_186), .ZN(
      n_1_737_1483));
   INV_X1 i_1_737_1529 (.A(n_1_737_1484), .ZN(n_47));
   OAI21_X1 i_1_737_1530 (.A(n_1_737_1485), .B1(in_data[8]), .B2(n_1_737_1490), 
      .ZN(n_1_737_1484));
   OAI211_X1 i_1_737_1531 (.A(n_1_737_1486), .B(n_1_737_1490), .C1(n_1_737_5597), 
      .C2(n_1_737_2247), .ZN(n_1_737_1485));
   OAI221_X1 i_1_737_1532 (.A(n_1_737_2247), .B1(n_1_737_1488), .B2(n_1_737_1487), 
      .C1(in_data[16]), .C2(n_1_737_2241), .ZN(n_1_737_1486));
   OAI21_X1 i_1_737_1533 (.A(n_1_737_2241), .B1(n_1_737_5599), .B2(n_1_737_2244), 
      .ZN(n_1_737_1487));
   AOI21_X1 i_1_737_1534 (.A(n_1_737_1489), .B1(n_1_737_5601), .B2(n_1_737_2239), 
      .ZN(n_1_737_1488));
   OAI21_X1 i_1_737_1535 (.A(n_1_737_2244), .B1(in_data[24]), .B2(n_1_737_2239), 
      .ZN(n_1_737_1489));
   OAI21_X1 i_1_737_1536 (.A(n_192), .B1(n_1_737_5602), .B2(n_191), .ZN(
      n_1_737_1490));
   OAI21_X1 i_1_737_1537 (.A(n_1_737_1491), .B1(n_1_737_5596), .B2(n_1_737_1492), 
      .ZN(n_48));
   OAI221_X1 i_1_737_1538 (.A(n_1_737_1492), .B1(in_data[12]), .B2(n_1_737_2262), 
      .C1(n_1_737_2263), .C2(n_1_737_1493), .ZN(n_1_737_1491));
   OAI21_X1 i_1_737_1539 (.A(n_197), .B1(n_1_737_5602), .B2(n_196), .ZN(
      n_1_737_1492));
   AOI21_X1 i_1_737_1540 (.A(n_1_737_1494), .B1(n_1_737_5598), .B2(n_1_737_2258), 
      .ZN(n_1_737_1493));
   AOI211_X1 i_1_737_1541 (.A(n_1_737_2258), .B(n_1_737_1495), .C1(in_data[20]), 
      .C2(n_1_737_2260), .ZN(n_1_737_1494));
   AOI221_X1 i_1_737_1542 (.A(n_1_737_2260), .B1(n_1_737_5601), .B2(n_1_737_2256), 
      .C1(n_1_737_5600), .C2(n_1_737_2255), .ZN(n_1_737_1495));
   OAI21_X1 i_1_737_1543 (.A(n_1_737_1496), .B1(n_1_737_5596), .B2(n_1_737_1501), 
      .ZN(n_49));
   NAND2_X1 i_1_737_1544 (.A1(n_1_737_1501), .A2(n_1_737_1497), .ZN(n_1_737_1496));
   AOI21_X1 i_1_737_1545 (.A(n_1_737_1498), .B1(n_1_737_5597), .B2(n_1_737_2331), 
      .ZN(n_1_737_1497));
   AOI221_X1 i_1_737_1546 (.A(n_1_737_2331), .B1(n_1_737_2326), .B2(n_1_737_1499), 
      .C1(in_data[16]), .C2(n_1_737_2325), .ZN(n_1_737_1498));
   AOI21_X1 i_1_737_1547 (.A(n_1_737_1500), .B1(n_1_737_5599), .B2(n_1_737_2328), 
      .ZN(n_1_737_1499));
   AOI221_X1 i_1_737_1548 (.A(n_1_737_2328), .B1(in_data[28]), .B2(n_1_737_2323), 
      .C1(in_data[24]), .C2(n_1_737_2322), .ZN(n_1_737_1500));
   OAI21_X1 i_1_737_1549 (.A(n_211), .B1(n_1_737_5602), .B2(n_210), .ZN(
      n_1_737_1501));
   INV_X1 i_1_737_1550 (.A(n_1_737_1502), .ZN(n_50));
   OAI21_X1 i_1_737_1551 (.A(n_1_737_1503), .B1(in_data[8]), .B2(n_1_737_1504), 
      .ZN(n_1_737_1502));
   OAI211_X1 i_1_737_1552 (.A(n_1_737_1504), .B(n_1_737_1505), .C1(n_1_737_5597), 
      .C2(n_1_737_2365), .ZN(n_1_737_1503));
   OAI21_X1 i_1_737_1553 (.A(n_219), .B1(n_1_737_5602), .B2(n_218), .ZN(
      n_1_737_1504));
   OAI221_X1 i_1_737_1554 (.A(n_1_737_2365), .B1(n_1_737_1507), .B2(n_1_737_1506), 
      .C1(in_data[16]), .C2(n_1_737_2354), .ZN(n_1_737_1505));
   OAI21_X1 i_1_737_1555 (.A(n_1_737_2354), .B1(n_1_737_5599), .B2(n_1_737_2356), 
      .ZN(n_1_737_1506));
   AOI21_X1 i_1_737_1556 (.A(n_1_737_1508), .B1(n_1_737_5600), .B2(n_1_737_2359), 
      .ZN(n_1_737_1507));
   OAI21_X1 i_1_737_1557 (.A(n_1_737_2356), .B1(in_data[28]), .B2(n_1_737_2359), 
      .ZN(n_1_737_1508));
   INV_X1 i_1_737_1558 (.A(n_1_737_1509), .ZN(n_51));
   OAI21_X1 i_1_737_1559 (.A(n_1_737_1510), .B1(in_data[8]), .B2(n_1_737_1511), 
      .ZN(n_1_737_1509));
   OAI211_X1 i_1_737_1560 (.A(n_1_737_1511), .B(n_1_737_1512), .C1(n_1_737_5597), 
      .C2(n_1_737_2380), .ZN(n_1_737_1510));
   OAI21_X1 i_1_737_1561 (.A(n_224), .B1(n_1_737_5602), .B2(n_223), .ZN(
      n_1_737_1511));
   OAI221_X1 i_1_737_1562 (.A(n_1_737_2380), .B1(n_1_737_1514), .B2(n_1_737_1513), 
      .C1(in_data[16]), .C2(n_1_737_2369), .ZN(n_1_737_1512));
   OAI21_X1 i_1_737_1563 (.A(n_1_737_2369), .B1(n_1_737_5599), .B2(n_1_737_2371), 
      .ZN(n_1_737_1513));
   AOI21_X1 i_1_737_1564 (.A(n_1_737_1515), .B1(n_1_737_5600), .B2(n_1_737_2374), 
      .ZN(n_1_737_1514));
   OAI21_X1 i_1_737_1565 (.A(n_1_737_2371), .B1(in_data[28]), .B2(n_1_737_2374), 
      .ZN(n_1_737_1515));
   OAI21_X1 i_1_737_1566 (.A(n_1_737_1516), .B1(n_1_737_5596), .B2(n_1_737_1520), 
      .ZN(n_52));
   OAI221_X1 i_1_737_1567 (.A(n_1_737_1520), .B1(in_data[12]), .B2(n_1_737_2415), 
      .C1(n_1_737_2414), .C2(n_1_737_1517), .ZN(n_1_737_1516));
   AOI21_X1 i_1_737_1568 (.A(n_1_737_1518), .B1(n_1_737_5598), .B2(n_1_737_2406), 
      .ZN(n_1_737_1517));
   AOI211_X1 i_1_737_1569 (.A(n_1_737_2406), .B(n_1_737_1519), .C1(in_data[20]), 
      .C2(n_1_737_2410), .ZN(n_1_737_1518));
   AOI221_X1 i_1_737_1570 (.A(n_1_737_2410), .B1(n_1_737_5600), .B2(n_1_737_2402), 
      .C1(n_1_737_5601), .C2(n_1_737_2401), .ZN(n_1_737_1519));
   OAI21_X1 i_1_737_1571 (.A(n_230), .B1(n_1_737_5602), .B2(n_229), .ZN(
      n_1_737_1520));
   OAI21_X1 i_1_737_1572 (.A(n_1_737_1521), .B1(n_1_737_5596), .B2(n_1_737_1525), 
      .ZN(n_53));
   OAI221_X1 i_1_737_1573 (.A(n_1_737_1525), .B1(in_data[12]), .B2(n_1_737_2431), 
      .C1(n_1_737_2430), .C2(n_1_737_1522), .ZN(n_1_737_1521));
   AOI21_X1 i_1_737_1574 (.A(n_1_737_1523), .B1(n_1_737_5598), .B2(n_1_737_2424), 
      .ZN(n_1_737_1522));
   AOI211_X1 i_1_737_1575 (.A(n_1_737_2424), .B(n_1_737_1524), .C1(in_data[20]), 
      .C2(n_1_737_2427), .ZN(n_1_737_1523));
   AOI221_X1 i_1_737_1576 (.A(n_1_737_2427), .B1(n_1_737_5601), .B2(n_1_737_2422), 
      .C1(n_1_737_5600), .C2(n_1_737_2421), .ZN(n_1_737_1524));
   OAI21_X1 i_1_737_1577 (.A(n_235), .B1(n_1_737_5602), .B2(n_234), .ZN(
      n_1_737_1525));
   AOI22_X1 i_1_737_1578 (.A1(n_1_737_5596), .A2(n_1_737_1530), .B1(n_1_737_1531), 
      .B2(n_1_737_1526), .ZN(n_54));
   OAI21_X1 i_1_737_1579 (.A(n_1_737_1527), .B1(in_data[12]), .B2(n_1_737_2450), 
      .ZN(n_1_737_1526));
   OAI221_X1 i_1_737_1580 (.A(n_1_737_2450), .B1(n_1_737_2439), .B2(n_1_737_1528), 
      .C1(n_1_737_5598), .C2(n_1_737_2440), .ZN(n_1_737_1527));
   AOI21_X1 i_1_737_1581 (.A(n_1_737_1529), .B1(in_data[20]), .B2(n_1_737_2443), 
      .ZN(n_1_737_1528));
   AOI221_X1 i_1_737_1582 (.A(n_1_737_2443), .B1(n_1_737_5601), .B2(n_1_737_2448), 
      .C1(n_1_737_5600), .C2(n_1_737_2447), .ZN(n_1_737_1529));
   INV_X1 i_1_737_1583 (.A(n_1_737_1531), .ZN(n_1_737_1530));
   OAI21_X1 i_1_737_1584 (.A(n_240), .B1(n_1_737_5602), .B2(n_239), .ZN(
      n_1_737_1531));
   OAI22_X1 i_1_737_1585 (.A1(n_1_737_1533), .A2(n_1_737_1532), .B1(n_1_737_5596), 
      .B2(n_1_737_1536), .ZN(n_55));
   OAI21_X1 i_1_737_1586 (.A(n_1_737_1536), .B1(in_data[12]), .B2(n_1_737_2486), 
      .ZN(n_1_737_1532));
   AOI211_X1 i_1_737_1587 (.A(n_1_737_1534), .B(n_1_737_2485), .C1(in_data[16]), 
      .C2(n_1_737_2472), .ZN(n_1_737_1533));
   AOI211_X1 i_1_737_1588 (.A(n_1_737_1535), .B(n_1_737_2472), .C1(n_1_737_5599), 
      .C2(n_1_737_2475), .ZN(n_1_737_1534));
   AOI221_X1 i_1_737_1589 (.A(n_1_737_2475), .B1(in_data[28]), .B2(n_1_737_2480), 
      .C1(in_data[24]), .C2(n_1_737_2479), .ZN(n_1_737_1535));
   OAI21_X1 i_1_737_1590 (.A(n_250), .B1(n_1_737_5602), .B2(n_249), .ZN(
      n_1_737_1536));
   OAI21_X1 i_1_737_1591 (.A(n_1_737_1537), .B1(n_1_737_5596), .B2(n_1_737_1542), 
      .ZN(n_56));
   OAI211_X1 i_1_737_1592 (.A(n_1_737_1538), .B(n_1_737_1542), .C1(in_data[12]), 
      .C2(n_1_737_2517), .ZN(n_1_737_1537));
   OAI211_X1 i_1_737_1593 (.A(n_1_737_1539), .B(n_1_737_2517), .C1(n_1_737_5598), 
      .C2(n_1_737_2506), .ZN(n_1_737_1538));
   NAND2_X1 i_1_737_1594 (.A1(n_1_737_2506), .A2(n_1_737_1540), .ZN(n_1_737_1539));
   OAI21_X1 i_1_737_1595 (.A(n_1_737_1541), .B1(n_1_737_5599), .B2(n_1_737_2508), 
      .ZN(n_1_737_1540));
   OAI221_X1 i_1_737_1596 (.A(n_1_737_2508), .B1(in_data[28]), .B2(n_1_737_2511), 
      .C1(in_data[24]), .C2(n_1_737_2512), .ZN(n_1_737_1541));
   OAI21_X1 i_1_737_1597 (.A(n_258), .B1(n_1_737_5602), .B2(n_257), .ZN(
      n_1_737_1542));
   OAI21_X1 i_1_737_1598 (.A(n_1_737_1543), .B1(n_1_737_5596), .B2(n_1_737_1545), 
      .ZN(n_57));
   OAI211_X1 i_1_737_1599 (.A(n_1_737_1545), .B(n_1_737_1544), .C1(in_data[12]), 
      .C2(n_1_737_2570), .ZN(n_1_737_1543));
   OAI221_X1 i_1_737_1600 (.A(n_1_737_2570), .B1(n_1_737_2565), .B2(n_1_737_1546), 
      .C1(n_1_737_5598), .C2(n_1_737_2566), .ZN(n_1_737_1544));
   OAI21_X1 i_1_737_1601 (.A(n_269), .B1(n_1_737_5602), .B2(n_268), .ZN(
      n_1_737_1545));
   AOI21_X1 i_1_737_1602 (.A(n_1_737_1547), .B1(in_data[20]), .B2(n_1_737_2556), 
      .ZN(n_1_737_1546));
   AOI221_X1 i_1_737_1603 (.A(n_1_737_2556), .B1(n_1_737_5601), .B2(n_1_737_2562), 
      .C1(n_1_737_5600), .C2(n_1_737_2561), .ZN(n_1_737_1547));
   OAI22_X1 i_1_737_1604 (.A1(n_1_737_2600), .A2(n_1_737_1548), .B1(n_1_737_5596), 
      .B2(n_1_737_2599), .ZN(n_58));
   OAI21_X1 i_1_737_1605 (.A(n_1_737_1549), .B1(in_data[12]), .B2(n_1_737_2606), 
      .ZN(n_1_737_1548));
   OAI211_X1 i_1_737_1606 (.A(n_1_737_1550), .B(n_1_737_2606), .C1(n_1_737_5598), 
      .C2(n_1_737_2602), .ZN(n_1_737_1549));
   OAI211_X1 i_1_737_1607 (.A(n_1_737_1551), .B(n_1_737_2602), .C1(in_data[20]), 
      .C2(n_1_737_2604), .ZN(n_1_737_1550));
   OAI221_X1 i_1_737_1608 (.A(n_1_737_2604), .B1(n_1_737_5601), .B2(n_1_737_2594), 
      .C1(n_1_737_5600), .C2(n_1_737_2595), .ZN(n_1_737_1551));
   INV_X1 i_1_737_1609 (.A(n_1_737_1552), .ZN(n_59));
   OAI21_X1 i_1_737_1610 (.A(n_1_737_1553), .B1(in_data[8]), .B2(n_1_737_1558), 
      .ZN(n_1_737_1552));
   OAI211_X1 i_1_737_1611 (.A(n_1_737_1554), .B(n_1_737_1558), .C1(n_1_737_5597), 
      .C2(n_1_737_2663), .ZN(n_1_737_1553));
   OAI221_X1 i_1_737_1612 (.A(n_1_737_2663), .B1(n_1_737_1556), .B2(n_1_737_1555), 
      .C1(in_data[16]), .C2(n_1_737_2649), .ZN(n_1_737_1554));
   OAI21_X1 i_1_737_1613 (.A(n_1_737_2649), .B1(n_1_737_5599), .B2(n_1_737_2652), 
      .ZN(n_1_737_1555));
   AOI21_X1 i_1_737_1614 (.A(n_1_737_1557), .B1(n_1_737_5600), .B2(n_1_737_2656), 
      .ZN(n_1_737_1556));
   OAI21_X1 i_1_737_1615 (.A(n_1_737_2652), .B1(in_data[28]), .B2(n_1_737_2656), 
      .ZN(n_1_737_1557));
   OAI21_X1 i_1_737_1616 (.A(n_288), .B1(n_1_737_5602), .B2(n_287), .ZN(
      n_1_737_1558));
   OAI21_X1 i_1_737_1617 (.A(n_1_737_1559), .B1(n_1_737_5596), .B2(n_1_737_1560), 
      .ZN(n_60));
   OAI221_X1 i_1_737_1618 (.A(n_1_737_1560), .B1(in_data[12]), .B2(n_1_737_2681), 
      .C1(n_1_737_2680), .C2(n_1_737_1561), .ZN(n_1_737_1559));
   OAI21_X1 i_1_737_1619 (.A(n_293), .B1(n_1_737_5602), .B2(n_292), .ZN(
      n_1_737_1560));
   AOI21_X1 i_1_737_1620 (.A(n_1_737_1562), .B1(n_1_737_5598), .B2(n_1_737_2674), 
      .ZN(n_1_737_1561));
   AOI221_X1 i_1_737_1621 (.A(n_1_737_2674), .B1(n_1_737_2678), .B2(n_1_737_1563), 
      .C1(in_data[20]), .C2(n_1_737_2677), .ZN(n_1_737_1562));
   AOI22_X1 i_1_737_1622 (.A1(n_1_737_5601), .A2(n_1_737_2670), .B1(n_1_737_5600), 
      .B2(n_1_737_2669), .ZN(n_1_737_1563));
   INV_X1 i_1_737_1623 (.A(n_1_737_1564), .ZN(n_61));
   OAI21_X1 i_1_737_1624 (.A(n_1_737_1565), .B1(in_data[8]), .B2(n_1_737_1569), 
      .ZN(n_1_737_1564));
   OAI211_X1 i_1_737_1625 (.A(n_1_737_1566), .B(n_1_737_1569), .C1(n_1_737_5597), 
      .C2(n_1_737_2702), .ZN(n_1_737_1565));
   OAI221_X1 i_1_737_1626 (.A(n_1_737_2702), .B1(n_1_737_2691), .B2(n_1_737_1567), 
      .C1(in_data[16]), .C2(n_1_737_2692), .ZN(n_1_737_1566));
   AOI22_X1 i_1_737_1627 (.A1(n_1_737_2694), .A2(n_1_737_1568), .B1(n_1_737_5599), 
      .B2(n_1_737_2695), .ZN(n_1_737_1567));
   OAI22_X1 i_1_737_1628 (.A1(in_data[28]), .A2(n_1_737_2698), .B1(in_data[24]), 
      .B2(n_1_737_2699), .ZN(n_1_737_1568));
   OAI21_X1 i_1_737_1629 (.A(n_296), .B1(n_1_737_5602), .B2(n_295), .ZN(
      n_1_737_1569));
   OAI21_X1 i_1_737_1630 (.A(n_1_737_1570), .B1(n_1_737_5596), .B2(n_1_737_1575), 
      .ZN(n_62));
   OAI211_X1 i_1_737_1631 (.A(n_1_737_1571), .B(n_1_737_1575), .C1(in_data[12]), 
      .C2(n_1_737_2722), .ZN(n_1_737_1570));
   NAND2_X1 i_1_737_1632 (.A1(n_1_737_2722), .A2(n_1_737_1572), .ZN(n_1_737_1571));
   AOI21_X1 i_1_737_1633 (.A(n_1_737_1573), .B1(in_data[16]), .B2(n_1_737_2719), 
      .ZN(n_1_737_1572));
   AOI211_X1 i_1_737_1634 (.A(n_1_737_1574), .B(n_1_737_2719), .C1(n_1_737_5599), 
      .C2(n_1_737_2709), .ZN(n_1_737_1573));
   AOI221_X1 i_1_737_1635 (.A(n_1_737_2709), .B1(in_data[28]), .B2(n_1_737_2715), 
      .C1(in_data[24]), .C2(n_1_737_2714), .ZN(n_1_737_1574));
   OAI21_X1 i_1_737_1636 (.A(n_299), .B1(n_1_737_5602), .B2(n_298), .ZN(
      n_1_737_1575));
   OAI22_X1 i_1_737_1637 (.A1(n_1_737_5596), .A2(n_1_737_1581), .B1(n_1_737_1580), 
      .B2(n_1_737_1576), .ZN(n_63));
   AOI21_X1 i_1_737_1638 (.A(n_1_737_1577), .B1(in_data[12]), .B2(n_1_737_2741), 
      .ZN(n_1_737_1576));
   AOI221_X1 i_1_737_1639 (.A(n_1_737_2741), .B1(n_1_737_2731), .B2(n_1_737_1578), 
      .C1(n_1_737_5598), .C2(n_1_737_2730), .ZN(n_1_737_1577));
   AOI22_X1 i_1_737_1640 (.A1(n_1_737_2739), .A2(n_1_737_1579), .B1(in_data[20]), 
      .B2(n_1_737_2738), .ZN(n_1_737_1578));
   OAI22_X1 i_1_737_1641 (.A1(n_1_737_5601), .A2(n_1_737_2735), .B1(n_1_737_5600), 
      .B2(n_1_737_2736), .ZN(n_1_737_1579));
   INV_X1 i_1_737_1642 (.A(n_1_737_1581), .ZN(n_1_737_1580));
   OAI21_X1 i_1_737_1643 (.A(n_302), .B1(n_1_737_5602), .B2(n_301), .ZN(
      n_1_737_1581));
   OAI21_X1 i_1_737_1644 (.A(n_1_737_1582), .B1(n_1_737_5596), .B2(n_1_737_1586), 
      .ZN(n_64));
   OAI211_X1 i_1_737_1645 (.A(n_1_737_1583), .B(n_1_737_1586), .C1(in_data[12]), 
      .C2(n_1_737_2756), .ZN(n_1_737_1582));
   OAI211_X1 i_1_737_1646 (.A(n_1_737_1584), .B(n_1_737_2756), .C1(n_1_737_5598), 
      .C2(n_1_737_2747), .ZN(n_1_737_1583));
   OAI211_X1 i_1_737_1647 (.A(n_1_737_1585), .B(n_1_737_2747), .C1(in_data[20]), 
      .C2(n_1_737_2745), .ZN(n_1_737_1584));
   OAI221_X1 i_1_737_1648 (.A(n_1_737_2745), .B1(n_1_737_5601), .B2(n_1_737_2751), 
      .C1(n_1_737_5600), .C2(n_1_737_2752), .ZN(n_1_737_1585));
   OAI21_X1 i_1_737_1649 (.A(n_307), .B1(n_1_737_5602), .B2(n_306), .ZN(
      n_1_737_1586));
   AOI22_X1 i_1_737_1650 (.A1(n_1_737_5596), .A2(n_1_737_1591), .B1(n_1_737_1592), 
      .B2(n_1_737_1587), .ZN(n_65));
   OAI21_X1 i_1_737_1651 (.A(n_1_737_1588), .B1(in_data[12]), .B2(n_1_737_2775), 
      .ZN(n_1_737_1587));
   OAI221_X1 i_1_737_1652 (.A(n_1_737_2775), .B1(n_1_737_2760), .B2(n_1_737_1589), 
      .C1(n_1_737_5598), .C2(n_1_737_2761), .ZN(n_1_737_1588));
   AOI21_X1 i_1_737_1653 (.A(n_1_737_1590), .B1(in_data[20]), .B2(n_1_737_2764), 
      .ZN(n_1_737_1589));
   AOI221_X1 i_1_737_1654 (.A(n_1_737_2764), .B1(n_1_737_5601), .B2(n_1_737_2770), 
      .C1(n_1_737_5600), .C2(n_1_737_2769), .ZN(n_1_737_1590));
   INV_X1 i_1_737_1655 (.A(n_1_737_1592), .ZN(n_1_737_1591));
   OAI21_X1 i_1_737_1656 (.A(n_310), .B1(n_1_737_5602), .B2(n_309), .ZN(
      n_1_737_1592));
   OAI21_X1 i_1_737_1657 (.A(n_1_737_1593), .B1(n_1_737_5596), .B2(n_1_737_1598), 
      .ZN(n_66));
   NAND2_X1 i_1_737_1658 (.A1(n_1_737_1598), .A2(n_1_737_1594), .ZN(n_1_737_1593));
   AOI21_X1 i_1_737_1659 (.A(n_1_737_1595), .B1(n_1_737_5597), .B2(n_1_737_2794), 
      .ZN(n_1_737_1594));
   AOI211_X1 i_1_737_1660 (.A(n_1_737_1596), .B(n_1_737_2794), .C1(in_data[16]), 
      .C2(n_1_737_2790), .ZN(n_1_737_1595));
   AOI211_X1 i_1_737_1661 (.A(n_1_737_1597), .B(n_1_737_2790), .C1(n_1_737_5599), 
      .C2(n_1_737_2784), .ZN(n_1_737_1596));
   AOI221_X1 i_1_737_1662 (.A(n_1_737_2784), .B1(in_data[28]), .B2(n_1_737_2786), 
      .C1(in_data[24]), .C2(n_1_737_2787), .ZN(n_1_737_1597));
   OAI21_X1 i_1_737_1663 (.A(n_315), .B1(n_1_737_5602), .B2(n_314), .ZN(
      n_1_737_1598));
   AOI22_X1 i_1_737_1664 (.A1(n_1_737_5596), .A2(n_1_737_1603), .B1(n_1_737_1604), 
      .B2(n_1_737_1599), .ZN(n_67));
   OAI21_X1 i_1_737_1665 (.A(n_1_737_1600), .B1(in_data[12]), .B2(n_1_737_2814), 
      .ZN(n_1_737_1599));
   OAI221_X1 i_1_737_1666 (.A(n_1_737_2814), .B1(n_1_737_2799), .B2(n_1_737_1601), 
      .C1(n_1_737_5598), .C2(n_1_737_2800), .ZN(n_1_737_1600));
   AOI21_X1 i_1_737_1667 (.A(n_1_737_1602), .B1(in_data[20]), .B2(n_1_737_2803), 
      .ZN(n_1_737_1601));
   AOI221_X1 i_1_737_1668 (.A(n_1_737_2803), .B1(n_1_737_5601), .B2(n_1_737_2809), 
      .C1(n_1_737_5600), .C2(n_1_737_2808), .ZN(n_1_737_1602));
   INV_X1 i_1_737_1669 (.A(n_1_737_1604), .ZN(n_1_737_1603));
   OAI21_X1 i_1_737_1670 (.A(n_318), .B1(n_1_737_5602), .B2(n_317), .ZN(
      n_1_737_1604));
   OAI21_X1 i_1_737_1671 (.A(n_1_737_1605), .B1(n_1_737_5596), .B2(n_1_737_1609), 
      .ZN(n_68));
   OAI221_X1 i_1_737_1672 (.A(n_1_737_1609), .B1(n_1_737_2827), .B2(n_1_737_1606), 
      .C1(in_data[12]), .C2(n_1_737_2828), .ZN(n_1_737_1605));
   AOI21_X1 i_1_737_1673 (.A(n_1_737_1607), .B1(n_1_737_5598), .B2(n_1_737_2821), 
      .ZN(n_1_737_1606));
   AOI211_X1 i_1_737_1674 (.A(n_1_737_1608), .B(n_1_737_2821), .C1(in_data[20]), 
      .C2(n_1_737_2824), .ZN(n_1_737_1607));
   AOI221_X1 i_1_737_1675 (.A(n_1_737_2824), .B1(n_1_737_5600), .B2(n_1_737_2818), 
      .C1(n_1_737_5601), .C2(n_1_737_2819), .ZN(n_1_737_1608));
   OAI21_X1 i_1_737_1676 (.A(n_323), .B1(n_1_737_5602), .B2(n_322), .ZN(
      n_1_737_1609));
   OAI21_X1 i_1_737_1677 (.A(n_1_737_1610), .B1(n_1_737_5596), .B2(n_1_737_1614), 
      .ZN(n_69));
   OAI221_X1 i_1_737_1678 (.A(n_1_737_1614), .B1(n_1_737_2848), .B2(n_1_737_1611), 
      .C1(in_data[12]), .C2(n_1_737_2849), .ZN(n_1_737_1610));
   OAI22_X1 i_1_737_1679 (.A1(n_1_737_1613), .A2(n_1_737_1612), .B1(n_1_737_5598), 
      .B2(n_1_737_2845), .ZN(n_1_737_1611));
   OAI21_X1 i_1_737_1680 (.A(n_1_737_2845), .B1(in_data[20]), .B2(n_1_737_2836), 
      .ZN(n_1_737_1612));
   AOI221_X1 i_1_737_1681 (.A(n_1_737_2835), .B1(in_data[28]), .B2(n_1_737_2842), 
      .C1(in_data[24]), .C2(n_1_737_2841), .ZN(n_1_737_1613));
   OAI21_X1 i_1_737_1682 (.A(n_326), .B1(n_1_737_5602), .B2(n_325), .ZN(
      n_1_737_1614));
   OAI21_X1 i_1_737_1683 (.A(n_1_737_1615), .B1(n_1_737_5596), .B2(n_1_737_1620), 
      .ZN(n_70));
   OAI211_X1 i_1_737_1684 (.A(n_1_737_1616), .B(n_1_737_1620), .C1(in_data[12]), 
      .C2(n_1_737_2867), .ZN(n_1_737_1615));
   OAI211_X1 i_1_737_1685 (.A(n_1_737_1617), .B(n_1_737_2867), .C1(n_1_737_5598), 
      .C2(n_1_737_2864), .ZN(n_1_737_1616));
   NAND2_X1 i_1_737_1686 (.A1(n_1_737_2864), .A2(n_1_737_1618), .ZN(n_1_737_1617));
   OAI21_X1 i_1_737_1687 (.A(n_1_737_1619), .B1(n_1_737_5599), .B2(n_1_737_2856), 
      .ZN(n_1_737_1618));
   OAI221_X1 i_1_737_1688 (.A(n_1_737_2856), .B1(in_data[24]), .B2(n_1_737_2861), 
      .C1(in_data[28]), .C2(n_1_737_2860), .ZN(n_1_737_1619));
   OAI21_X1 i_1_737_1689 (.A(n_329), .B1(n_1_737_5602), .B2(n_328), .ZN(
      n_1_737_1620));
   AOI22_X1 i_1_737_1690 (.A1(n_1_737_5596), .A2(n_1_737_1625), .B1(n_1_737_1626), 
      .B2(n_1_737_1621), .ZN(n_71));
   OAI21_X1 i_1_737_1691 (.A(n_1_737_1622), .B1(in_data[12]), .B2(n_1_737_2887), 
      .ZN(n_1_737_1621));
   OAI221_X1 i_1_737_1692 (.A(n_1_737_2887), .B1(n_1_737_2872), .B2(n_1_737_1623), 
      .C1(n_1_737_5598), .C2(n_1_737_2873), .ZN(n_1_737_1622));
   AOI21_X1 i_1_737_1693 (.A(n_1_737_1624), .B1(in_data[20]), .B2(n_1_737_2876), 
      .ZN(n_1_737_1623));
   AOI221_X1 i_1_737_1694 (.A(n_1_737_2876), .B1(n_1_737_5601), .B2(n_1_737_2882), 
      .C1(n_1_737_5600), .C2(n_1_737_2881), .ZN(n_1_737_1624));
   INV_X1 i_1_737_1695 (.A(n_1_737_1626), .ZN(n_1_737_1625));
   OAI21_X1 i_1_737_1696 (.A(n_332), .B1(n_1_737_5602), .B2(n_331), .ZN(
      n_1_737_1626));
   OAI22_X1 i_1_737_1697 (.A1(n_1_737_5596), .A2(n_1_737_1632), .B1(n_1_737_1631), 
      .B2(n_1_737_1627), .ZN(n_72));
   AOI22_X1 i_1_737_1698 (.A1(in_data[12]), .A2(n_1_737_2918), .B1(n_1_737_2917), 
      .B2(n_1_737_1628), .ZN(n_1_737_1627));
   OAI21_X1 i_1_737_1699 (.A(n_1_737_1629), .B1(n_1_737_5598), .B2(n_1_737_2915), 
      .ZN(n_1_737_1628));
   OAI221_X1 i_1_737_1700 (.A(n_1_737_2915), .B1(n_1_737_2912), .B2(n_1_737_1630), 
      .C1(in_data[20]), .C2(n_1_737_2911), .ZN(n_1_737_1629));
   AOI22_X1 i_1_737_1701 (.A1(n_1_737_5601), .A2(n_1_737_2907), .B1(n_1_737_5600), 
      .B2(n_1_737_2908), .ZN(n_1_737_1630));
   INV_X1 i_1_737_1702 (.A(n_1_737_1632), .ZN(n_1_737_1631));
   OAI21_X1 i_1_737_1703 (.A(n_342), .B1(n_1_737_5602), .B2(n_341), .ZN(
      n_1_737_1632));
   OAI22_X1 i_1_737_1704 (.A1(n_1_737_5596), .A2(n_1_737_1640), .B1(n_1_737_1639), 
      .B2(n_1_737_1633), .ZN(n_73));
   OAI21_X1 i_1_737_1705 (.A(n_1_737_1634), .B1(in_data[12]), .B2(n_1_737_2936), 
      .ZN(n_1_737_1633));
   OAI211_X1 i_1_737_1706 (.A(n_1_737_1635), .B(n_1_737_2936), .C1(n_1_737_5598), 
      .C2(n_1_737_2929), .ZN(n_1_737_1634));
   OAI21_X1 i_1_737_1707 (.A(n_1_737_2929), .B1(n_1_737_1637), .B2(n_1_737_1636), 
      .ZN(n_1_737_1635));
   NOR2_X1 i_1_737_1708 (.A1(n_1_737_5599), .A2(n_1_737_2931), .ZN(n_1_737_1636));
   AOI21_X1 i_1_737_1709 (.A(n_1_737_1638), .B1(n_1_737_5600), .B2(n_1_737_2933), 
      .ZN(n_1_737_1637));
   OAI21_X1 i_1_737_1710 (.A(n_1_737_2931), .B1(in_data[28]), .B2(n_1_737_2933), 
      .ZN(n_1_737_1638));
   INV_X1 i_1_737_1711 (.A(n_1_737_1640), .ZN(n_1_737_1639));
   OAI21_X1 i_1_737_1712 (.A(n_347), .B1(n_1_737_5602), .B2(n_346), .ZN(
      n_1_737_1640));
   OAI21_X1 i_1_737_1713 (.A(n_1_737_1641), .B1(n_1_737_5596), .B2(n_1_737_1646), 
      .ZN(n_74));
   NAND2_X1 i_1_737_1714 (.A1(n_1_737_1646), .A2(n_1_737_1642), .ZN(n_1_737_1641));
   AOI21_X1 i_1_737_1715 (.A(n_1_737_1643), .B1(n_1_737_5597), .B2(n_1_737_2957), 
      .ZN(n_1_737_1642));
   AOI211_X1 i_1_737_1716 (.A(n_1_737_1644), .B(n_1_737_2957), .C1(in_data[16]), 
      .C2(n_1_737_2942), .ZN(n_1_737_1643));
   AOI211_X1 i_1_737_1717 (.A(n_1_737_1645), .B(n_1_737_2942), .C1(n_1_737_5599), 
      .C2(n_1_737_2946), .ZN(n_1_737_1644));
   AOI221_X1 i_1_737_1718 (.A(n_1_737_2946), .B1(in_data[28]), .B2(n_1_737_2951), 
      .C1(in_data[24]), .C2(n_1_737_2950), .ZN(n_1_737_1645));
   OAI21_X1 i_1_737_1719 (.A(n_350), .B1(n_1_737_5602), .B2(n_349), .ZN(
      n_1_737_1646));
   OAI21_X1 i_1_737_1720 (.A(n_1_737_1647), .B1(n_1_737_5596), .B2(n_1_737_1651), 
      .ZN(n_75));
   OAI221_X1 i_1_737_1721 (.A(n_1_737_1651), .B1(in_data[12]), .B2(n_1_737_2969), 
      .C1(n_1_737_2970), .C2(n_1_737_1648), .ZN(n_1_737_1647));
   AOI21_X1 i_1_737_1722 (.A(n_1_737_1649), .B1(n_1_737_5598), .B2(n_1_737_2965), 
      .ZN(n_1_737_1648));
   AOI211_X1 i_1_737_1723 (.A(n_1_737_1650), .B(n_1_737_2965), .C1(in_data[20]), 
      .C2(n_1_737_2967), .ZN(n_1_737_1649));
   AOI221_X1 i_1_737_1724 (.A(n_1_737_2967), .B1(n_1_737_5601), .B2(n_1_737_2963), 
      .C1(n_1_737_5600), .C2(n_1_737_2962), .ZN(n_1_737_1650));
   OAI21_X1 i_1_737_1725 (.A(n_355), .B1(n_1_737_5602), .B2(n_354), .ZN(
      n_1_737_1651));
   AOI22_X1 i_1_737_1726 (.A1(n_1_737_5596), .A2(n_1_737_1656), .B1(n_1_737_1657), 
      .B2(n_1_737_1652), .ZN(n_76));
   OAI21_X1 i_1_737_1727 (.A(n_1_737_1653), .B1(in_data[12]), .B2(n_1_737_2994), 
      .ZN(n_1_737_1652));
   OAI221_X1 i_1_737_1728 (.A(n_1_737_2994), .B1(n_1_737_2990), .B2(n_1_737_1654), 
      .C1(n_1_737_5598), .C2(n_1_737_2991), .ZN(n_1_737_1653));
   AOI21_X1 i_1_737_1729 (.A(n_1_737_1655), .B1(in_data[20]), .B2(n_1_737_2980), 
      .ZN(n_1_737_1654));
   AOI221_X1 i_1_737_1730 (.A(n_1_737_2980), .B1(n_1_737_5601), .B2(n_1_737_2987), 
      .C1(n_1_737_5600), .C2(n_1_737_2986), .ZN(n_1_737_1655));
   INV_X1 i_1_737_1731 (.A(n_1_737_1657), .ZN(n_1_737_1656));
   OAI21_X1 i_1_737_1732 (.A(n_360), .B1(n_1_737_5602), .B2(n_359), .ZN(
      n_1_737_1657));
   OAI22_X1 i_1_737_1733 (.A1(n_1_737_5596), .A2(n_1_737_1661), .B1(n_1_737_1660), 
      .B2(n_1_737_1658), .ZN(n_77));
   NAND2_X1 i_1_737_1734 (.A1(n_1_737_1661), .A2(n_1_737_1659), .ZN(n_1_737_1658));
   OAI221_X1 i_1_737_1735 (.A(n_1_737_3020), .B1(n_1_737_3002), .B2(n_1_737_1662), 
      .C1(n_1_737_5598), .C2(n_1_737_3003), .ZN(n_1_737_1659));
   NOR2_X1 i_1_737_1736 (.A1(in_data[12]), .A2(n_1_737_3020), .ZN(n_1_737_1660));
   OAI21_X1 i_1_737_1737 (.A(n_365), .B1(n_1_737_5602), .B2(n_364), .ZN(
      n_1_737_1661));
   AOI21_X1 i_1_737_1738 (.A(n_1_737_1663), .B1(in_data[20]), .B2(n_1_737_3007), 
      .ZN(n_1_737_1662));
   AOI221_X1 i_1_737_1739 (.A(n_1_737_3007), .B1(n_1_737_5601), .B2(n_1_737_3012), 
      .C1(n_1_737_5600), .C2(n_1_737_3013), .ZN(n_1_737_1663));
   OAI21_X1 i_1_737_1740 (.A(n_1_737_1664), .B1(n_1_737_5596), .B2(n_1_737_1669), 
      .ZN(n_78));
   OAI211_X1 i_1_737_1741 (.A(n_1_737_1665), .B(n_1_737_1669), .C1(in_data[12]), 
      .C2(n_1_737_3040), .ZN(n_1_737_1664));
   OAI211_X1 i_1_737_1742 (.A(n_1_737_1666), .B(n_1_737_3040), .C1(n_1_737_5598), 
      .C2(n_1_737_3037), .ZN(n_1_737_1665));
   NAND2_X1 i_1_737_1743 (.A1(n_1_737_3037), .A2(n_1_737_1667), .ZN(n_1_737_1666));
   OAI21_X1 i_1_737_1744 (.A(n_1_737_1668), .B1(n_1_737_5599), .B2(n_1_737_3029), 
      .ZN(n_1_737_1667));
   OAI221_X1 i_1_737_1745 (.A(n_1_737_3029), .B1(in_data[28]), .B2(n_1_737_3033), 
      .C1(in_data[24]), .C2(n_1_737_3034), .ZN(n_1_737_1668));
   OAI21_X1 i_1_737_1746 (.A(n_370), .B1(n_1_737_5602), .B2(n_369), .ZN(
      n_1_737_1669));
   OAI21_X1 i_1_737_1747 (.A(n_1_737_1670), .B1(n_1_737_5596), .B2(n_1_737_1675), 
      .ZN(n_79));
   NAND2_X1 i_1_737_1748 (.A1(n_1_737_1675), .A2(n_1_737_1671), .ZN(n_1_737_1670));
   AOI21_X1 i_1_737_1749 (.A(n_1_737_1672), .B1(n_1_737_5597), .B2(n_1_737_3076), 
      .ZN(n_1_737_1671));
   AOI221_X1 i_1_737_1750 (.A(n_1_737_3076), .B1(n_1_737_3064), .B2(n_1_737_1673), 
      .C1(in_data[16]), .C2(n_1_737_3063), .ZN(n_1_737_1672));
   AOI22_X1 i_1_737_1751 (.A1(n_1_737_3068), .A2(n_1_737_1674), .B1(n_1_737_5599), 
      .B2(n_1_737_3067), .ZN(n_1_737_1673));
   OAI22_X1 i_1_737_1752 (.A1(in_data[28]), .A2(n_1_737_3071), .B1(in_data[24]), 
      .B2(n_1_737_3072), .ZN(n_1_737_1674));
   OAI21_X1 i_1_737_1753 (.A(n_376), .B1(n_1_737_5602), .B2(n_375), .ZN(
      n_1_737_1675));
   OAI21_X1 i_1_737_1754 (.A(n_1_737_1676), .B1(n_1_737_5596), .B2(n_1_737_1681), 
      .ZN(n_80));
   OAI211_X1 i_1_737_1755 (.A(n_1_737_1677), .B(n_1_737_1681), .C1(in_data[12]), 
      .C2(n_1_737_3102), .ZN(n_1_737_1676));
   NAND2_X1 i_1_737_1756 (.A1(n_1_737_3102), .A2(n_1_737_1678), .ZN(n_1_737_1677));
   AOI21_X1 i_1_737_1757 (.A(n_1_737_1679), .B1(in_data[16]), .B2(n_1_737_3099), 
      .ZN(n_1_737_1678));
   AOI221_X1 i_1_737_1758 (.A(n_1_737_3099), .B1(n_1_737_5599), .B2(n_1_737_3088), 
      .C1(n_1_737_3089), .C2(n_1_737_1680), .ZN(n_1_737_1679));
   AOI22_X1 i_1_737_1759 (.A1(in_data[28]), .A2(n_1_737_3095), .B1(in_data[24]), 
      .B2(n_1_737_3096), .ZN(n_1_737_1680));
   OAI21_X1 i_1_737_1760 (.A(n_381), .B1(n_1_737_5602), .B2(n_380), .ZN(
      n_1_737_1681));
   AOI22_X1 i_1_737_1761 (.A1(n_1_737_5596), .A2(n_1_737_1686), .B1(n_1_737_1687), 
      .B2(n_1_737_1682), .ZN(n_81));
   OAI21_X1 i_1_737_1762 (.A(n_1_737_1683), .B1(in_data[12]), .B2(n_1_737_3127), 
      .ZN(n_1_737_1682));
   OAI221_X1 i_1_737_1763 (.A(n_1_737_3127), .B1(n_1_737_3112), .B2(n_1_737_1684), 
      .C1(n_1_737_5598), .C2(n_1_737_3113), .ZN(n_1_737_1683));
   AOI21_X1 i_1_737_1764 (.A(n_1_737_1685), .B1(in_data[20]), .B2(n_1_737_3116), 
      .ZN(n_1_737_1684));
   AOI221_X1 i_1_737_1765 (.A(n_1_737_3116), .B1(n_1_737_5601), .B2(n_1_737_3122), 
      .C1(n_1_737_5600), .C2(n_1_737_3121), .ZN(n_1_737_1685));
   INV_X1 i_1_737_1766 (.A(n_1_737_1687), .ZN(n_1_737_1686));
   OAI21_X1 i_1_737_1767 (.A(n_384), .B1(n_1_737_5602), .B2(n_383), .ZN(
      n_1_737_1687));
   OAI21_X1 i_1_737_1768 (.A(n_1_737_1688), .B1(n_1_737_5596), .B2(n_1_737_1689), 
      .ZN(n_82));
   OAI211_X1 i_1_737_1769 (.A(n_1_737_1689), .B(n_1_737_1690), .C1(in_data[12]), 
      .C2(n_1_737_3190), .ZN(n_1_737_1688));
   AOI21_X1 i_1_737_1770 (.A(n_398), .B1(n_1_737_5602), .B2(n_399), .ZN(
      n_1_737_1689));
   OAI211_X1 i_1_737_1771 (.A(n_1_737_1691), .B(n_1_737_3190), .C1(n_1_737_5598), 
      .C2(n_1_737_3178), .ZN(n_1_737_1690));
   OAI211_X1 i_1_737_1772 (.A(n_1_737_1692), .B(n_1_737_3178), .C1(in_data[20]), 
      .C2(n_1_737_3186), .ZN(n_1_737_1691));
   OAI221_X1 i_1_737_1773 (.A(n_1_737_3186), .B1(n_1_737_5601), .B2(n_1_737_3173), 
      .C1(n_1_737_5600), .C2(n_1_737_3174), .ZN(n_1_737_1692));
   INV_X1 i_1_737_1774 (.A(n_1_737_1693), .ZN(n_83));
   OAI21_X1 i_1_737_1775 (.A(n_1_737_1694), .B1(in_data[8]), .B2(n_1_737_1699), 
      .ZN(n_1_737_1693));
   OAI211_X1 i_1_737_1776 (.A(n_1_737_1699), .B(n_1_737_1695), .C1(n_1_737_5597), 
      .C2(n_1_737_3215), .ZN(n_1_737_1694));
   OAI211_X1 i_1_737_1777 (.A(n_1_737_3215), .B(n_1_737_1696), .C1(in_data[16]), 
      .C2(n_1_737_3211), .ZN(n_1_737_1695));
   OAI221_X1 i_1_737_1778 (.A(n_1_737_3211), .B1(n_1_737_5599), .B2(n_1_737_3202), 
      .C1(n_1_737_1698), .C2(n_1_737_1697), .ZN(n_1_737_1696));
   OAI21_X1 i_1_737_1779 (.A(n_1_737_3202), .B1(in_data[24]), .B2(n_1_737_3207), 
      .ZN(n_1_737_1697));
   NOR2_X1 i_1_737_1780 (.A1(in_data[28]), .A2(n_1_737_3206), .ZN(n_1_737_1698));
   AOI21_X1 i_1_737_1781 (.A(n_403), .B1(n_1_737_5602), .B2(n_404), .ZN(
      n_1_737_1699));
   INV_X1 i_1_737_1782 (.A(n_1_737_1700), .ZN(n_84));
   OAI21_X1 i_1_737_1783 (.A(n_1_737_1701), .B1(in_data[8]), .B2(n_1_737_1706), 
      .ZN(n_1_737_1700));
   OAI211_X1 i_1_737_1784 (.A(n_1_737_1706), .B(n_1_737_1702), .C1(n_1_737_5597), 
      .C2(n_1_737_3232), .ZN(n_1_737_1701));
   OAI211_X1 i_1_737_1785 (.A(n_1_737_3232), .B(n_1_737_1703), .C1(in_data[16]), 
      .C2(n_1_737_3243), .ZN(n_1_737_1702));
   OAI221_X1 i_1_737_1786 (.A(n_1_737_3243), .B1(n_1_737_5599), .B2(n_1_737_3239), 
      .C1(n_1_737_1705), .C2(n_1_737_1704), .ZN(n_1_737_1703));
   OAI21_X1 i_1_737_1787 (.A(n_1_737_3239), .B1(in_data[28]), .B2(n_1_737_3227), 
      .ZN(n_1_737_1704));
   NOR2_X1 i_1_737_1788 (.A1(in_data[24]), .A2(n_1_737_3228), .ZN(n_1_737_1705));
   AOI21_X1 i_1_737_1789 (.A(n_408), .B1(n_1_737_5602), .B2(n_409), .ZN(
      n_1_737_1706));
   OAI21_X1 i_1_737_1790 (.A(n_1_737_1707), .B1(n_1_737_5596), .B2(n_1_737_1712), 
      .ZN(n_85));
   OAI21_X1 i_1_737_1791 (.A(n_1_737_1712), .B1(n_1_737_1709), .B2(n_1_737_1708), 
      .ZN(n_1_737_1707));
   NOR2_X1 i_1_737_1792 (.A1(n_1_737_5597), .A2(n_1_737_3269), .ZN(n_1_737_1708));
   AOI211_X1 i_1_737_1793 (.A(n_1_737_3270), .B(n_1_737_1710), .C1(n_1_737_5598), 
      .C2(n_1_737_3254), .ZN(n_1_737_1709));
   AOI211_X1 i_1_737_1794 (.A(n_1_737_3254), .B(n_1_737_1711), .C1(in_data[20]), 
      .C2(n_1_737_3264), .ZN(n_1_737_1710));
   AOI221_X1 i_1_737_1795 (.A(n_1_737_3264), .B1(n_1_737_5600), .B2(n_1_737_3259), 
      .C1(n_1_737_5601), .C2(n_1_737_3258), .ZN(n_1_737_1711));
   AOI21_X1 i_1_737_1796 (.A(n_413), .B1(n_1_737_5602), .B2(n_414), .ZN(
      n_1_737_1712));
   OAI21_X1 i_1_737_1797 (.A(n_1_737_1713), .B1(n_1_737_5596), .B2(n_1_737_1714), 
      .ZN(n_86));
   OAI211_X1 i_1_737_1798 (.A(n_1_737_1714), .B(n_1_737_1715), .C1(in_data[12]), 
      .C2(n_1_737_3296), .ZN(n_1_737_1713));
   AOI21_X1 i_1_737_1799 (.A(n_418), .B1(n_1_737_5602), .B2(n_419), .ZN(
      n_1_737_1714));
   OAI211_X1 i_1_737_1800 (.A(n_1_737_1716), .B(n_1_737_3296), .C1(n_1_737_5598), 
      .C2(n_1_737_3283), .ZN(n_1_737_1715));
   OAI211_X1 i_1_737_1801 (.A(n_1_737_1717), .B(n_1_737_3283), .C1(in_data[20]), 
      .C2(n_1_737_3292), .ZN(n_1_737_1716));
   OAI221_X1 i_1_737_1802 (.A(n_1_737_3292), .B1(n_1_737_5601), .B2(n_1_737_3278), 
      .C1(n_1_737_5600), .C2(n_1_737_3279), .ZN(n_1_737_1717));
   OAI21_X1 i_1_737_1803 (.A(n_1_737_1718), .B1(n_1_737_5596), .B2(n_1_737_1722), 
      .ZN(n_87));
   OAI211_X1 i_1_737_1804 (.A(n_1_737_1719), .B(n_1_737_1722), .C1(in_data[12]), 
      .C2(n_1_737_3323), .ZN(n_1_737_1718));
   OAI221_X1 i_1_737_1805 (.A(n_1_737_3323), .B1(n_1_737_3307), .B2(n_1_737_1720), 
      .C1(n_1_737_5598), .C2(n_1_737_3308), .ZN(n_1_737_1719));
   AOI21_X1 i_1_737_1806 (.A(n_1_737_1721), .B1(in_data[20]), .B2(n_1_737_3318), 
      .ZN(n_1_737_1720));
   AOI221_X1 i_1_737_1807 (.A(n_1_737_3318), .B1(n_1_737_5600), .B2(n_1_737_3312), 
      .C1(n_1_737_5601), .C2(n_1_737_3313), .ZN(n_1_737_1721));
   AOI21_X1 i_1_737_1808 (.A(n_423), .B1(n_1_737_5602), .B2(n_424), .ZN(
      n_1_737_1722));
   OAI21_X1 i_1_737_1809 (.A(n_1_737_1723), .B1(n_1_737_5596), .B2(n_1_737_1724), 
      .ZN(n_88));
   OAI211_X1 i_1_737_1810 (.A(n_1_737_1724), .B(n_1_737_1725), .C1(in_data[12]), 
      .C2(n_1_737_3338), .ZN(n_1_737_1723));
   AOI21_X1 i_1_737_1811 (.A(n_428), .B1(n_1_737_5602), .B2(n_429), .ZN(
      n_1_737_1724));
   OAI211_X1 i_1_737_1812 (.A(n_1_737_1726), .B(n_1_737_3338), .C1(n_1_737_5598), 
      .C2(n_1_737_3335), .ZN(n_1_737_1725));
   OAI211_X1 i_1_737_1813 (.A(n_1_737_1727), .B(n_1_737_3335), .C1(in_data[20]), 
      .C2(n_1_737_3343), .ZN(n_1_737_1726));
   OAI221_X1 i_1_737_1814 (.A(n_1_737_3343), .B1(n_1_737_5601), .B2(n_1_737_3346), 
      .C1(n_1_737_5600), .C2(n_1_737_3347), .ZN(n_1_737_1727));
   INV_X1 i_1_737_1815 (.A(n_1_737_1728), .ZN(n_89));
   OAI21_X1 i_1_737_1816 (.A(n_1_737_1729), .B1(in_data[8]), .B2(n_1_737_1734), 
      .ZN(n_1_737_1728));
   OAI211_X1 i_1_737_1817 (.A(n_1_737_1734), .B(n_1_737_1730), .C1(n_1_737_5597), 
      .C2(n_1_737_3376), .ZN(n_1_737_1729));
   OAI21_X1 i_1_737_1818 (.A(n_1_737_1731), .B1(in_data[16]), .B2(n_1_737_3359), 
      .ZN(n_1_737_1730));
   NOR2_X1 i_1_737_1819 (.A1(n_1_737_3377), .A2(n_1_737_1732), .ZN(n_1_737_1731));
   AOI211_X1 i_1_737_1820 (.A(n_1_737_3358), .B(n_1_737_1733), .C1(in_data[20]), 
      .C2(n_1_737_3370), .ZN(n_1_737_1732));
   AOI221_X1 i_1_737_1821 (.A(n_1_737_3370), .B1(n_1_737_5601), .B2(n_1_737_3364), 
      .C1(n_1_737_5600), .C2(n_1_737_3365), .ZN(n_1_737_1733));
   AOI21_X1 i_1_737_1822 (.A(n_432), .B1(n_1_737_5602), .B2(n_433), .ZN(
      n_1_737_1734));
   INV_X1 i_1_737_1823 (.A(n_1_737_1735), .ZN(n_90));
   OAI21_X1 i_1_737_1824 (.A(n_1_737_1736), .B1(in_data[8]), .B2(n_1_737_1740), 
      .ZN(n_1_737_1735));
   OAI221_X1 i_1_737_1825 (.A(n_1_737_1740), .B1(n_1_737_5597), .B2(n_1_737_3411), 
      .C1(n_1_737_3412), .C2(n_1_737_1737), .ZN(n_1_737_1736));
   AOI22_X1 i_1_737_1826 (.A1(n_1_737_3394), .A2(n_1_737_1738), .B1(in_data[16]), 
      .B2(n_1_737_3393), .ZN(n_1_737_1737));
   OAI22_X1 i_1_737_1827 (.A1(n_1_737_3388), .A2(n_1_737_1739), .B1(n_1_737_5599), 
      .B2(n_1_737_3387), .ZN(n_1_737_1738));
   AOI22_X1 i_1_737_1828 (.A1(in_data[28]), .A2(n_1_737_3404), .B1(in_data[24]), 
      .B2(n_1_737_3405), .ZN(n_1_737_1739));
   AOI21_X1 i_1_737_1829 (.A(n_437), .B1(n_1_737_5602), .B2(n_438), .ZN(
      n_1_737_1740));
   OAI21_X1 i_1_737_1830 (.A(n_1_737_1741), .B1(n_1_737_5596), .B2(n_1_737_1746), 
      .ZN(n_91));
   OAI21_X1 i_1_737_1831 (.A(n_1_737_1746), .B1(n_1_737_1743), .B2(n_1_737_1742), 
      .ZN(n_1_737_1741));
   NOR2_X1 i_1_737_1832 (.A1(n_1_737_5597), .A2(n_1_737_3447), .ZN(n_1_737_1742));
   AOI211_X1 i_1_737_1833 (.A(n_1_737_3448), .B(n_1_737_1744), .C1(n_1_737_5598), 
      .C2(n_1_737_3428), .ZN(n_1_737_1743));
   AOI211_X1 i_1_737_1834 (.A(n_1_737_3428), .B(n_1_737_1745), .C1(in_data[20]), 
      .C2(n_1_737_3441), .ZN(n_1_737_1744));
   AOI221_X1 i_1_737_1835 (.A(n_1_737_3441), .B1(n_1_737_5600), .B2(n_1_737_3433), 
      .C1(n_1_737_5601), .C2(n_1_737_3434), .ZN(n_1_737_1745));
   AOI21_X1 i_1_737_1836 (.A(n_442), .B1(n_1_737_5602), .B2(n_443), .ZN(
      n_1_737_1746));
   OAI21_X1 i_1_737_1837 (.A(n_1_737_1747), .B1(n_1_737_5596), .B2(n_1_737_1748), 
      .ZN(n_92));
   OAI211_X1 i_1_737_1838 (.A(n_1_737_1748), .B(n_1_737_1749), .C1(in_data[12]), 
      .C2(n_1_737_3476), .ZN(n_1_737_1747));
   AOI21_X1 i_1_737_1839 (.A(n_447), .B1(n_1_737_5602), .B2(n_448), .ZN(
      n_1_737_1748));
   OAI211_X1 i_1_737_1840 (.A(n_1_737_1750), .B(n_1_737_3476), .C1(n_1_737_5598), 
      .C2(n_1_737_3466), .ZN(n_1_737_1749));
   OAI211_X1 i_1_737_1841 (.A(n_1_737_1751), .B(n_1_737_3466), .C1(in_data[20]), 
      .C2(n_1_737_3469), .ZN(n_1_737_1750));
   OAI221_X1 i_1_737_1842 (.A(n_1_737_3469), .B1(n_1_737_5601), .B2(n_1_737_3462), 
      .C1(n_1_737_5600), .C2(n_1_737_3463), .ZN(n_1_737_1751));
   INV_X1 i_1_737_1843 (.A(n_1_737_1752), .ZN(n_93));
   OAI21_X1 i_1_737_1844 (.A(n_1_737_1753), .B1(in_data[8]), .B2(n_1_737_1758), 
      .ZN(n_1_737_1752));
   OAI211_X1 i_1_737_1845 (.A(n_1_737_1758), .B(n_1_737_1754), .C1(n_1_737_5597), 
      .C2(n_1_737_3499), .ZN(n_1_737_1753));
   OAI211_X1 i_1_737_1846 (.A(n_1_737_3499), .B(n_1_737_1755), .C1(in_data[16]), 
      .C2(n_1_737_3490), .ZN(n_1_737_1754));
   OAI221_X1 i_1_737_1847 (.A(n_1_737_3490), .B1(n_1_737_5599), .B2(n_1_737_3495), 
      .C1(n_1_737_1757), .C2(n_1_737_1756), .ZN(n_1_737_1755));
   OAI21_X1 i_1_737_1848 (.A(n_1_737_3495), .B1(in_data[28]), .B2(n_1_737_3484), 
      .ZN(n_1_737_1756));
   NOR2_X1 i_1_737_1849 (.A1(in_data[24]), .A2(n_1_737_3485), .ZN(n_1_737_1757));
   AOI21_X1 i_1_737_1850 (.A(n_452), .B1(n_1_737_5602), .B2(n_453), .ZN(
      n_1_737_1758));
   INV_X1 i_1_737_1851 (.A(n_1_737_1759), .ZN(n_94));
   OAI21_X1 i_1_737_1852 (.A(n_1_737_1760), .B1(in_data[8]), .B2(n_1_737_1766), 
      .ZN(n_1_737_1759));
   OAI221_X1 i_1_737_1853 (.A(n_1_737_1766), .B1(n_1_737_5597), .B2(n_1_737_3537), 
      .C1(n_1_737_3538), .C2(n_1_737_1761), .ZN(n_1_737_1760));
   INV_X1 i_1_737_1854 (.A(n_1_737_1762), .ZN(n_1_737_1761));
   OAI21_X1 i_1_737_1855 (.A(n_1_737_1763), .B1(n_1_737_5598), .B2(n_1_737_3515), 
      .ZN(n_1_737_1762));
   OAI21_X1 i_1_737_1856 (.A(n_1_737_3515), .B1(n_1_737_1765), .B2(n_1_737_1764), 
      .ZN(n_1_737_1763));
   AND2_X1 i_1_737_1857 (.A1(in_data[20]), .A2(n_1_737_3531), .ZN(n_1_737_1764));
   AOI221_X1 i_1_737_1858 (.A(n_1_737_3531), .B1(n_1_737_5601), .B2(n_1_737_3523), 
      .C1(n_1_737_5600), .C2(n_1_737_3524), .ZN(n_1_737_1765));
   AOI21_X1 i_1_737_1859 (.A(n_457), .B1(n_1_737_5602), .B2(n_458), .ZN(
      n_1_737_1766));
   INV_X1 i_1_737_1860 (.A(n_1_737_1767), .ZN(n_95));
   OAI21_X1 i_1_737_1861 (.A(n_1_737_1768), .B1(in_data[8]), .B2(n_1_737_1773), 
      .ZN(n_1_737_1767));
   OAI211_X1 i_1_737_1862 (.A(n_1_737_1773), .B(n_1_737_1769), .C1(n_1_737_5597), 
      .C2(n_1_737_3567), .ZN(n_1_737_1768));
   OAI211_X1 i_1_737_1863 (.A(n_1_737_3567), .B(n_1_737_1770), .C1(in_data[16]), 
      .C2(n_1_737_3554), .ZN(n_1_737_1769));
   OAI221_X1 i_1_737_1864 (.A(n_1_737_3554), .B1(n_1_737_5599), .B2(n_1_737_3559), 
      .C1(n_1_737_1772), .C2(n_1_737_1771), .ZN(n_1_737_1770));
   OAI21_X1 i_1_737_1865 (.A(n_1_737_3559), .B1(in_data[24]), .B2(n_1_737_3549), 
      .ZN(n_1_737_1771));
   AND2_X1 i_1_737_1866 (.A1(n_1_737_5601), .A2(n_1_737_3549), .ZN(n_1_737_1772));
   AOI21_X1 i_1_737_1867 (.A(n_462), .B1(n_1_737_5602), .B2(n_463), .ZN(
      n_1_737_1773));
   OAI21_X1 i_1_737_1868 (.A(n_1_737_1774), .B1(n_1_737_5596), .B2(n_1_737_1778), 
      .ZN(n_96));
   OAI221_X1 i_1_737_1869 (.A(n_1_737_1778), .B1(n_1_737_3721), .B2(n_1_737_1775), 
      .C1(in_data[12]), .C2(n_1_737_3720), .ZN(n_1_737_1774));
   AOI22_X1 i_1_737_1870 (.A1(n_1_737_3705), .A2(n_1_737_1776), .B1(n_1_737_5598), 
      .B2(n_1_737_3704), .ZN(n_1_737_1775));
   AOI21_X1 i_1_737_1871 (.A(n_1_737_1777), .B1(in_data[20]), .B2(n_1_737_3715), 
      .ZN(n_1_737_1776));
   AOI221_X1 i_1_737_1872 (.A(n_1_737_3715), .B1(n_1_737_5600), .B2(n_1_737_3710), 
      .C1(n_1_737_5601), .C2(n_1_737_3709), .ZN(n_1_737_1777));
   AOI21_X1 i_1_737_1873 (.A(n_489), .B1(n_1_737_5602), .B2(n_490), .ZN(
      n_1_737_1778));
   OAI21_X1 i_1_737_1874 (.A(n_1_737_1779), .B1(n_1_737_5596), .B2(n_1_737_1780), 
      .ZN(n_97));
   OAI211_X1 i_1_737_1875 (.A(n_1_737_1780), .B(n_1_737_1781), .C1(in_data[12]), 
      .C2(n_1_737_3742), .ZN(n_1_737_1779));
   AOI21_X1 i_1_737_1876 (.A(n_494), .B1(n_1_737_5602), .B2(n_495), .ZN(
      n_1_737_1780));
   OAI211_X1 i_1_737_1877 (.A(n_1_737_1782), .B(n_1_737_3742), .C1(n_1_737_5598), 
      .C2(n_1_737_3730), .ZN(n_1_737_1781));
   OAI211_X1 i_1_737_1878 (.A(n_1_737_1783), .B(n_1_737_3730), .C1(in_data[20]), 
      .C2(n_1_737_3738), .ZN(n_1_737_1782));
   OAI221_X1 i_1_737_1879 (.A(n_1_737_3738), .B1(n_1_737_5601), .B2(n_1_737_3734), 
      .C1(n_1_737_5600), .C2(n_1_737_3733), .ZN(n_1_737_1783));
   INV_X1 i_1_737_1880 (.A(n_1_737_1784), .ZN(n_98));
   OAI21_X1 i_1_737_1881 (.A(n_1_737_1785), .B1(in_data[8]), .B2(n_1_737_1786), 
      .ZN(n_1_737_1784));
   OAI221_X1 i_1_737_1882 (.A(n_1_737_1786), .B1(n_1_737_5597), .B2(n_1_737_3800), 
      .C1(n_1_737_1789), .C2(n_1_737_1787), .ZN(n_1_737_1785));
   AOI21_X1 i_1_737_1883 (.A(n_499), .B1(n_1_737_5602), .B2(n_500), .ZN(
      n_1_737_1786));
   OAI21_X1 i_1_737_1884 (.A(n_1_737_3800), .B1(n_1_737_1790), .B2(n_1_737_1788), 
      .ZN(n_1_737_1787));
   OAI21_X1 i_1_737_1885 (.A(n_1_737_3790), .B1(n_1_737_5599), .B2(n_1_737_3770), 
      .ZN(n_1_737_1788));
   NOR2_X1 i_1_737_1886 (.A1(in_data[16]), .A2(n_1_737_3790), .ZN(n_1_737_1789));
   AOI21_X1 i_1_737_1887 (.A(n_1_737_1791), .B1(n_1_737_5600), .B2(n_1_737_3779), 
      .ZN(n_1_737_1790));
   OAI21_X1 i_1_737_1888 (.A(n_1_737_3770), .B1(in_data[28]), .B2(n_1_737_3779), 
      .ZN(n_1_737_1791));
   INV_X1 i_1_737_1889 (.A(n_1_737_1792), .ZN(n_99));
   OAI21_X1 i_1_737_1890 (.A(n_1_737_1793), .B1(in_data[8]), .B2(n_1_737_1797), 
      .ZN(n_1_737_1792));
   OAI211_X1 i_1_737_1891 (.A(n_1_737_1797), .B(n_1_737_1794), .C1(n_1_737_5597), 
      .C2(n_1_737_3852), .ZN(n_1_737_1793));
   OAI211_X1 i_1_737_1892 (.A(n_1_737_3852), .B(n_1_737_1795), .C1(in_data[16]), 
      .C2(n_1_737_3836), .ZN(n_1_737_1794));
   OAI211_X1 i_1_737_1893 (.A(n_1_737_3836), .B(n_1_737_1796), .C1(n_1_737_5599), 
      .C2(n_1_737_3848), .ZN(n_1_737_1795));
   OAI221_X1 i_1_737_1894 (.A(n_1_737_3848), .B1(in_data[28]), .B2(n_1_737_3843), 
      .C1(in_data[24]), .C2(n_1_737_3842), .ZN(n_1_737_1796));
   AOI21_X1 i_1_737_1895 (.A(n_509), .B1(n_1_737_5602), .B2(n_510), .ZN(
      n_1_737_1797));
   INV_X1 i_1_737_1896 (.A(n_1_737_1798), .ZN(n_100));
   OAI21_X1 i_1_737_1897 (.A(n_1_737_1799), .B1(in_data[8]), .B2(n_1_737_1804), 
      .ZN(n_1_737_1798));
   OAI211_X1 i_1_737_1898 (.A(n_1_737_1804), .B(n_1_737_1800), .C1(n_1_737_5597), 
      .C2(n_1_737_3877), .ZN(n_1_737_1799));
   OAI211_X1 i_1_737_1899 (.A(n_1_737_3877), .B(n_1_737_1801), .C1(in_data[16]), 
      .C2(n_1_737_3865), .ZN(n_1_737_1800));
   OAI221_X1 i_1_737_1900 (.A(n_1_737_3865), .B1(n_1_737_5599), .B2(n_1_737_3869), 
      .C1(n_1_737_1803), .C2(n_1_737_1802), .ZN(n_1_737_1801));
   OAI21_X1 i_1_737_1901 (.A(n_1_737_3869), .B1(in_data[28]), .B2(n_1_737_3860), 
      .ZN(n_1_737_1802));
   NOR2_X1 i_1_737_1902 (.A1(in_data[24]), .A2(n_1_737_3859), .ZN(n_1_737_1803));
   AOI21_X1 i_1_737_1903 (.A(n_514), .B1(n_1_737_5602), .B2(n_515), .ZN(
      n_1_737_1804));
   INV_X1 i_1_737_1904 (.A(n_1_737_1805), .ZN(n_101));
   OAI21_X1 i_1_737_1905 (.A(n_1_737_1806), .B1(in_data[8]), .B2(n_1_737_1810), 
      .ZN(n_1_737_1805));
   OAI221_X1 i_1_737_1906 (.A(n_1_737_1810), .B1(n_1_737_5597), .B2(n_1_737_3935), 
      .C1(n_1_737_3934), .C2(n_1_737_1807), .ZN(n_1_737_1806));
   AOI22_X1 i_1_737_1907 (.A1(n_1_737_3923), .A2(n_1_737_1808), .B1(in_data[16]), 
      .B2(n_1_737_3922), .ZN(n_1_737_1807));
   OAI22_X1 i_1_737_1908 (.A1(n_1_737_3926), .A2(n_1_737_1809), .B1(n_1_737_5599), 
      .B2(n_1_737_3927), .ZN(n_1_737_1808));
   AOI22_X1 i_1_737_1909 (.A1(in_data[28]), .A2(n_1_737_3917), .B1(in_data[24]), 
      .B2(n_1_737_3918), .ZN(n_1_737_1809));
   AOI21_X1 i_1_737_1910 (.A(n_524), .B1(n_1_737_5602), .B2(n_525), .ZN(
      n_1_737_1810));
   OAI21_X1 i_1_737_1911 (.A(n_1_737_1811), .B1(n_1_737_5596), .B2(n_1_737_1815), 
      .ZN(n_102));
   OAI221_X1 i_1_737_1912 (.A(n_1_737_1815), .B1(n_1_737_3972), .B2(n_1_737_1812), 
      .C1(in_data[12]), .C2(n_1_737_3971), .ZN(n_1_737_1811));
   AOI22_X1 i_1_737_1913 (.A1(n_1_737_3953), .A2(n_1_737_1813), .B1(n_1_737_5598), 
      .B2(n_1_737_3952), .ZN(n_1_737_1812));
   AOI21_X1 i_1_737_1914 (.A(n_1_737_1814), .B1(in_data[20]), .B2(n_1_737_3946), 
      .ZN(n_1_737_1813));
   AOI221_X1 i_1_737_1915 (.A(n_1_737_3946), .B1(n_1_737_5600), .B2(n_1_737_3965), 
      .C1(n_1_737_5601), .C2(n_1_737_3964), .ZN(n_1_737_1814));
   AOI21_X1 i_1_737_1916 (.A(n_529), .B1(n_1_737_5602), .B2(n_530), .ZN(
      n_1_737_1815));
   OAI21_X1 i_1_737_1917 (.A(n_1_737_1816), .B1(n_1_737_5596), .B2(n_1_737_1820), 
      .ZN(n_103));
   OAI221_X1 i_1_737_1918 (.A(n_1_737_1820), .B1(n_1_737_3998), .B2(n_1_737_1817), 
      .C1(in_data[12]), .C2(n_1_737_3999), .ZN(n_1_737_1816));
   AOI22_X1 i_1_737_1919 (.A1(n_1_737_3989), .A2(n_1_737_1818), .B1(n_1_737_5598), 
      .B2(n_1_737_3988), .ZN(n_1_737_1817));
   OAI22_X1 i_1_737_1920 (.A1(n_1_737_3993), .A2(n_1_737_1819), .B1(in_data[20]), 
      .B2(n_1_737_3994), .ZN(n_1_737_1818));
   AOI22_X1 i_1_737_1921 (.A1(n_1_737_5600), .A2(n_1_737_3983), .B1(n_1_737_5601), 
      .B2(n_1_737_3982), .ZN(n_1_737_1819));
   AOI21_X1 i_1_737_1922 (.A(n_534), .B1(n_1_737_5602), .B2(n_535), .ZN(
      n_1_737_1820));
   OAI21_X1 i_1_737_1923 (.A(n_1_737_1821), .B1(n_1_737_5596), .B2(n_1_737_1825), 
      .ZN(n_104));
   OAI211_X1 i_1_737_1924 (.A(n_1_737_1822), .B(n_1_737_1825), .C1(in_data[12]), 
      .C2(n_1_737_4063), .ZN(n_1_737_1821));
   OAI211_X1 i_1_737_1925 (.A(n_1_737_4063), .B(n_1_737_1823), .C1(n_1_737_5598), 
      .C2(n_1_737_4030), .ZN(n_1_737_1822));
   OAI221_X1 i_1_737_1926 (.A(n_1_737_4030), .B1(n_1_737_4053), .B2(n_1_737_1824), 
      .C1(in_data[20]), .C2(n_1_737_4052), .ZN(n_1_737_1823));
   AOI22_X1 i_1_737_1927 (.A1(n_1_737_5600), .A2(n_1_737_4041), .B1(n_1_737_5601), 
      .B2(n_1_737_4040), .ZN(n_1_737_1824));
   AOI21_X1 i_1_737_1928 (.A(n_539), .B1(n_1_737_5602), .B2(n_540), .ZN(
      n_1_737_1825));
   OAI21_X1 i_1_737_1929 (.A(n_1_737_1826), .B1(n_1_737_5596), .B2(n_1_737_1832), 
      .ZN(n_105));
   NAND2_X1 i_1_737_1930 (.A1(n_1_737_1832), .A2(n_1_737_1827), .ZN(n_1_737_1826));
   OAI21_X1 i_1_737_1931 (.A(n_1_737_1828), .B1(n_1_737_5597), .B2(n_1_737_4078), 
      .ZN(n_1_737_1827));
   OAI211_X1 i_1_737_1932 (.A(n_1_737_4078), .B(n_1_737_1829), .C1(in_data[16]), 
      .C2(n_1_737_4085), .ZN(n_1_737_1828));
   OAI221_X1 i_1_737_1933 (.A(n_1_737_4085), .B1(n_1_737_5599), .B2(n_1_737_4088), 
      .C1(n_1_737_1831), .C2(n_1_737_1830), .ZN(n_1_737_1829));
   OAI21_X1 i_1_737_1934 (.A(n_1_737_4088), .B1(in_data[28]), .B2(n_1_737_4081), 
      .ZN(n_1_737_1830));
   NOR2_X1 i_1_737_1935 (.A1(in_data[24]), .A2(n_1_737_4082), .ZN(n_1_737_1831));
   AOI21_X1 i_1_737_1936 (.A(n_544), .B1(n_1_737_5602), .B2(n_545), .ZN(
      n_1_737_1832));
   INV_X1 i_1_737_1937 (.A(n_1_737_1833), .ZN(n_106));
   OAI21_X1 i_1_737_1938 (.A(n_1_737_1834), .B1(in_data[8]), .B2(n_1_737_1839), 
      .ZN(n_1_737_1833));
   OAI221_X1 i_1_737_1939 (.A(n_1_737_1839), .B1(n_1_737_5597), .B2(n_1_737_4097), 
      .C1(n_1_737_1837), .C2(n_1_737_1835), .ZN(n_1_737_1834));
   OAI21_X1 i_1_737_1940 (.A(n_1_737_4097), .B1(n_1_737_1838), .B2(n_1_737_1836), 
      .ZN(n_1_737_1835));
   OAI21_X1 i_1_737_1941 (.A(n_1_737_4109), .B1(n_1_737_5599), .B2(n_1_737_4102), 
      .ZN(n_1_737_1836));
   NOR2_X1 i_1_737_1942 (.A1(in_data[16]), .A2(n_1_737_4109), .ZN(n_1_737_1837));
   AOI221_X1 i_1_737_1943 (.A(n_1_737_4103), .B1(n_1_737_5601), .B2(n_1_737_4114), 
      .C1(n_1_737_5600), .C2(n_1_737_4115), .ZN(n_1_737_1838));
   AOI21_X1 i_1_737_1944 (.A(n_547), .B1(n_1_737_5602), .B2(n_548), .ZN(
      n_1_737_1839));
   OAI21_X1 i_1_737_1945 (.A(n_1_737_1840), .B1(n_1_737_5596), .B2(n_1_737_1841), 
      .ZN(n_107));
   OAI211_X1 i_1_737_1946 (.A(n_1_737_1841), .B(n_1_737_1842), .C1(in_data[12]), 
      .C2(n_1_737_4146), .ZN(n_1_737_1840));
   AOI21_X1 i_1_737_1947 (.A(n_551), .B1(n_1_737_5602), .B2(n_552), .ZN(
      n_1_737_1841));
   OAI211_X1 i_1_737_1948 (.A(n_1_737_1843), .B(n_1_737_4146), .C1(n_1_737_5598), 
      .C2(n_1_737_4128), .ZN(n_1_737_1842));
   OAI211_X1 i_1_737_1949 (.A(n_1_737_1844), .B(n_1_737_4128), .C1(in_data[20]), 
      .C2(n_1_737_4139), .ZN(n_1_737_1843));
   OAI221_X1 i_1_737_1950 (.A(n_1_737_4139), .B1(n_1_737_5601), .B2(n_1_737_4123), 
      .C1(n_1_737_5600), .C2(n_1_737_4122), .ZN(n_1_737_1844));
   INV_X1 i_1_737_1951 (.A(n_1_737_1845), .ZN(n_108));
   OAI21_X1 i_1_737_1952 (.A(n_1_737_1846), .B1(in_data[8]), .B2(n_1_737_1851), 
      .ZN(n_1_737_1845));
   OAI211_X1 i_1_737_1953 (.A(n_1_737_1847), .B(n_1_737_1851), .C1(n_1_737_5597), 
      .C2(n_1_737_4244), .ZN(n_1_737_1846));
   OAI211_X1 i_1_737_1954 (.A(n_1_737_4244), .B(n_1_737_1848), .C1(in_data[16]), 
      .C2(n_1_737_4219), .ZN(n_1_737_1847));
   OAI221_X1 i_1_737_1955 (.A(n_1_737_4219), .B1(n_1_737_5599), .B2(n_1_737_4227), 
      .C1(n_1_737_1850), .C2(n_1_737_1849), .ZN(n_1_737_1848));
   OAI21_X1 i_1_737_1956 (.A(n_1_737_4227), .B1(in_data[24]), .B2(n_1_737_4211), 
      .ZN(n_1_737_1849));
   NOR2_X1 i_1_737_1957 (.A1(in_data[28]), .A2(n_1_737_4212), .ZN(n_1_737_1850));
   AOI21_X1 i_1_737_1958 (.A(n_563), .B1(n_1_737_5602), .B2(n_564), .ZN(
      n_1_737_1851));
   OAI21_X1 i_1_737_1959 (.A(n_1_737_1852), .B1(n_1_737_5596), .B2(n_1_737_1853), 
      .ZN(n_109));
   OAI211_X1 i_1_737_1960 (.A(n_1_737_1853), .B(n_1_737_1854), .C1(in_data[12]), 
      .C2(n_1_737_4309), .ZN(n_1_737_1852));
   AOI21_X1 i_1_737_1961 (.A(n_571), .B1(n_1_737_5602), .B2(n_572), .ZN(
      n_1_737_1853));
   OAI211_X1 i_1_737_1962 (.A(n_1_737_1855), .B(n_1_737_4309), .C1(n_1_737_5598), 
      .C2(n_1_737_4304), .ZN(n_1_737_1854));
   OAI211_X1 i_1_737_1963 (.A(n_1_737_1856), .B(n_1_737_4304), .C1(in_data[20]), 
      .C2(n_1_737_4293), .ZN(n_1_737_1855));
   OAI221_X1 i_1_737_1964 (.A(n_1_737_4293), .B1(n_1_737_5601), .B2(n_1_737_4299), 
      .C1(n_1_737_5600), .C2(n_1_737_4298), .ZN(n_1_737_1856));
   OAI21_X1 i_1_737_1965 (.A(n_1_737_1857), .B1(n_1_737_5596), .B2(n_1_737_1862), 
      .ZN(n_110));
   OAI21_X1 i_1_737_1966 (.A(n_1_737_1862), .B1(n_1_737_1859), .B2(n_1_737_1858), 
      .ZN(n_1_737_1857));
   NOR2_X1 i_1_737_1967 (.A1(n_1_737_5597), .A2(n_1_737_4361), .ZN(n_1_737_1858));
   AOI211_X1 i_1_737_1968 (.A(n_1_737_4362), .B(n_1_737_1860), .C1(n_1_737_5598), 
      .C2(n_1_737_4342), .ZN(n_1_737_1859));
   AOI211_X1 i_1_737_1969 (.A(n_1_737_4342), .B(n_1_737_1861), .C1(in_data[20]), 
      .C2(n_1_737_4355), .ZN(n_1_737_1860));
   AOI221_X1 i_1_737_1970 (.A(n_1_737_4355), .B1(n_1_737_5601), .B2(n_1_737_4349), 
      .C1(n_1_737_5600), .C2(n_1_737_4350), .ZN(n_1_737_1861));
   AOI21_X1 i_1_737_1971 (.A(n_579), .B1(n_1_737_5602), .B2(n_580), .ZN(
      n_1_737_1862));
   OAI22_X1 i_1_737_1972 (.A1(n_1_737_1865), .A2(n_1_737_1863), .B1(n_1_737_5596), 
      .B2(n_1_737_1866), .ZN(n_111));
   AOI21_X1 i_1_737_1973 (.A(n_1_737_1864), .B1(in_data[12]), .B2(n_1_737_4393), 
      .ZN(n_1_737_1863));
   AOI211_X1 i_1_737_1974 (.A(n_1_737_1867), .B(n_1_737_4393), .C1(n_1_737_5598), 
      .C2(n_1_737_4376), .ZN(n_1_737_1864));
   INV_X1 i_1_737_1975 (.A(n_1_737_1866), .ZN(n_1_737_1865));
   AOI21_X1 i_1_737_1976 (.A(n_583), .B1(n_1_737_5602), .B2(n_584), .ZN(
      n_1_737_1866));
   INV_X1 i_1_737_1977 (.A(n_1_737_1868), .ZN(n_1_737_1867));
   OAI211_X1 i_1_737_1978 (.A(n_1_737_1869), .B(n_1_737_4377), .C1(n_1_737_5599), 
      .C2(n_1_737_4383), .ZN(n_1_737_1868));
   OAI221_X1 i_1_737_1979 (.A(n_1_737_4383), .B1(in_data[28]), .B2(n_1_737_4370), 
      .C1(in_data[24]), .C2(n_1_737_4369), .ZN(n_1_737_1869));
   AOI211_X1 i_1_737_1983 (.A(n_1_737_4417), .B(n_1_737_1873), .C1(in_data[20]), 
      .C2(n_1_737_4405), .ZN(n_1_737_1872));
   AOI221_X1 i_1_737_1984 (.A(n_1_737_4405), .B1(n_1_737_5601), .B2(n_1_737_4440), 
      .C1(n_1_737_5600), .C2(n_1_737_4441), .ZN(n_1_737_1873));
   OAI21_X1 i_1_737_1987 (.A(n_1_737_1876), .B1(n_1_737_5596), .B2(n_1_737_1877), 
      .ZN(n_112));
   OAI211_X1 i_1_737_1988 (.A(n_1_737_1877), .B(n_1_737_1878), .C1(in_data[12]), 
      .C2(n_1_737_4478), .ZN(n_1_737_1876));
   AOI21_X1 i_1_737_1989 (.A(n_589), .B1(n_1_737_5602), .B2(n_590), .ZN(
      n_1_737_1877));
   OAI211_X1 i_1_737_1990 (.A(n_1_737_1879), .B(n_1_737_4478), .C1(n_1_737_5598), 
      .C2(n_1_737_4469), .ZN(n_1_737_1878));
   OAI211_X1 i_1_737_1991 (.A(n_1_737_1880), .B(n_1_737_4469), .C1(in_data[20]), 
      .C2(n_1_737_4472), .ZN(n_1_737_1879));
   OAI221_X1 i_1_737_1992 (.A(n_1_737_4472), .B1(n_1_737_5601), .B2(n_1_737_4464), 
      .C1(n_1_737_5600), .C2(n_1_737_4465), .ZN(n_1_737_1880));
   OAI21_X1 i_1_737_1993 (.A(n_1_737_1881), .B1(n_1_737_5596), .B2(n_1_737_1885), 
      .ZN(n_113));
   OAI221_X1 i_1_737_1994 (.A(n_1_737_1885), .B1(n_1_737_4506), .B2(n_1_737_1882), 
      .C1(in_data[12]), .C2(n_1_737_4505), .ZN(n_1_737_1881));
   OAI22_X1 i_1_737_1995 (.A1(n_1_737_1884), .A2(n_1_737_1883), .B1(n_1_737_5598), 
      .B2(n_1_737_4487), .ZN(n_1_737_1882));
   OAI21_X1 i_1_737_1996 (.A(n_1_737_4487), .B1(in_data[20]), .B2(n_1_737_4499), 
      .ZN(n_1_737_1883));
   AOI221_X1 i_1_737_1997 (.A(n_1_737_4500), .B1(in_data[28]), .B2(n_1_737_4493), 
      .C1(in_data[24]), .C2(n_1_737_4494), .ZN(n_1_737_1884));
   AOI21_X1 i_1_737_1998 (.A(n_593), .B1(n_1_737_5602), .B2(n_594), .ZN(
      n_1_737_1885));
   INV_X1 i_1_737_1999 (.A(n_1_737_1886), .ZN(n_114));
   OAI21_X1 i_1_737_2000 (.A(n_1_737_1887), .B1(in_data[8]), .B2(n_1_737_1891), 
      .ZN(n_1_737_1886));
   OAI211_X1 i_1_737_2001 (.A(n_1_737_1888), .B(n_1_737_1891), .C1(n_1_737_5597), 
      .C2(n_1_737_4555), .ZN(n_1_737_1887));
   OAI211_X1 i_1_737_2002 (.A(n_1_737_4555), .B(n_1_737_1889), .C1(in_data[16]), 
      .C2(n_1_737_4529), .ZN(n_1_737_1888));
   OAI211_X1 i_1_737_2003 (.A(n_1_737_4529), .B(n_1_737_1890), .C1(n_1_737_5599), 
      .C2(n_1_737_4546), .ZN(n_1_737_1889));
   OAI221_X1 i_1_737_2004 (.A(n_1_737_4546), .B1(in_data[28]), .B2(n_1_737_4522), 
      .C1(in_data[24]), .C2(n_1_737_4521), .ZN(n_1_737_1890));
   AOI21_X1 i_1_737_2005 (.A(n_598), .B1(n_1_737_5602), .B2(n_599), .ZN(
      n_1_737_1891));
   OAI21_X1 i_1_737_2006 (.A(n_1_737_1892), .B1(n_1_737_5596), .B2(n_1_737_1893), 
      .ZN(n_115));
   OAI211_X1 i_1_737_2007 (.A(n_1_737_1893), .B(n_1_737_1894), .C1(in_data[12]), 
      .C2(n_1_737_4639), .ZN(n_1_737_1892));
   AOI21_X1 i_1_737_2008 (.A(n_609), .B1(n_1_737_5602), .B2(n_610), .ZN(
      n_1_737_1893));
   OAI211_X1 i_1_737_2009 (.A(n_1_737_1895), .B(n_1_737_4639), .C1(n_1_737_5598), 
      .C2(n_1_737_4618), .ZN(n_1_737_1894));
   OAI211_X1 i_1_737_2010 (.A(n_1_737_1896), .B(n_1_737_4618), .C1(in_data[20]), 
      .C2(n_1_737_4633), .ZN(n_1_737_1895));
   OAI221_X1 i_1_737_2011 (.A(n_1_737_4633), .B1(n_1_737_5601), .B2(n_1_737_4628), 
      .C1(n_1_737_5600), .C2(n_1_737_4627), .ZN(n_1_737_1896));
   OAI21_X1 i_1_737_2012 (.A(n_1_737_1897), .B1(n_1_737_5596), .B2(n_1_737_1901), 
      .ZN(n_116));
   OAI221_X1 i_1_737_2013 (.A(n_1_737_1901), .B1(n_1_737_4709), .B2(n_1_737_1898), 
      .C1(in_data[12]), .C2(n_1_737_4708), .ZN(n_1_737_1897));
   OAI21_X1 i_1_737_2014 (.A(n_1_737_1899), .B1(n_1_737_5598), .B2(n_1_737_4687), 
      .ZN(n_1_737_1898));
   OAI221_X1 i_1_737_2015 (.A(n_1_737_4687), .B1(n_1_737_4701), .B2(n_1_737_1900), 
      .C1(in_data[20]), .C2(n_1_737_4700), .ZN(n_1_737_1899));
   AOI22_X1 i_1_737_2016 (.A1(n_1_737_5600), .A2(n_1_737_4694), .B1(n_1_737_5601), 
      .B2(n_1_737_4693), .ZN(n_1_737_1900));
   AOI21_X1 i_1_737_2017 (.A(n_617), .B1(n_1_737_5602), .B2(n_618), .ZN(
      n_1_737_1901));
   OAI21_X1 i_1_737_2018 (.A(n_1_737_1902), .B1(n_1_737_5596), .B2(n_1_737_1906), 
      .ZN(n_117));
   OAI221_X1 i_1_737_2019 (.A(n_1_737_1906), .B1(n_1_737_1904), .B2(n_1_737_1903), 
      .C1(in_data[12]), .C2(n_1_737_4720), .ZN(n_1_737_1902));
   OAI21_X1 i_1_737_2020 (.A(n_1_737_4720), .B1(n_1_737_5598), .B2(n_1_737_4729), 
      .ZN(n_1_737_1903));
   AOI211_X1 i_1_737_2021 (.A(n_1_737_1905), .B(n_1_737_4728), .C1(n_1_737_5599), 
      .C2(n_1_737_4732), .ZN(n_1_737_1904));
   AOI221_X1 i_1_737_2022 (.A(n_1_737_4732), .B1(in_data[28]), .B2(n_1_737_4725), 
      .C1(in_data[24]), .C2(n_1_737_4724), .ZN(n_1_737_1905));
   AOI21_X1 i_1_737_2023 (.A(n_621), .B1(n_1_737_5602), .B2(n_622), .ZN(
      n_1_737_1906));
   OAI21_X1 i_1_737_2024 (.A(n_1_737_1907), .B1(n_1_737_5596), .B2(n_1_737_1911), 
      .ZN(n_118));
   OAI211_X1 i_1_737_2025 (.A(n_1_737_1908), .B(n_1_737_1911), .C1(in_data[12]), 
      .C2(n_1_737_4782), .ZN(n_1_737_1907));
   OAI211_X1 i_1_737_2026 (.A(n_1_737_4782), .B(n_1_737_1909), .C1(n_1_737_5598), 
      .C2(n_1_737_4754), .ZN(n_1_737_1908));
   OAI211_X1 i_1_737_2027 (.A(n_1_737_1910), .B(n_1_737_4754), .C1(in_data[20]), 
      .C2(n_1_737_4764), .ZN(n_1_737_1909));
   OAI221_X1 i_1_737_2028 (.A(n_1_737_4764), .B1(n_1_737_5601), .B2(n_1_737_4743), 
      .C1(n_1_737_5600), .C2(n_1_737_4744), .ZN(n_1_737_1910));
   AOI21_X1 i_1_737_2029 (.A(n_625), .B1(n_1_737_5602), .B2(n_626), .ZN(
      n_1_737_1911));
   OAI21_X1 i_1_737_2030 (.A(n_1_737_1912), .B1(n_1_737_5596), .B2(n_1_737_1913), 
      .ZN(n_119));
   OAI211_X1 i_1_737_2031 (.A(n_1_737_1913), .B(n_1_737_1914), .C1(in_data[12]), 
      .C2(n_1_737_4805), .ZN(n_1_737_1912));
   AOI21_X1 i_1_737_2032 (.A(n_629), .B1(n_1_737_5602), .B2(n_630), .ZN(
      n_1_737_1913));
   OAI211_X1 i_1_737_2033 (.A(n_1_737_1915), .B(n_1_737_4805), .C1(n_1_737_5598), 
      .C2(n_1_737_4795), .ZN(n_1_737_1914));
   OAI211_X1 i_1_737_2034 (.A(n_1_737_1916), .B(n_1_737_4795), .C1(in_data[20]), 
      .C2(n_1_737_4801), .ZN(n_1_737_1915));
   OAI221_X1 i_1_737_2035 (.A(n_1_737_4801), .B1(n_1_737_5601), .B2(n_1_737_4792), 
      .C1(n_1_737_5600), .C2(n_1_737_4793), .ZN(n_1_737_1916));
   INV_X1 i_1_737_2036 (.A(n_1_737_1917), .ZN(n_120));
   OAI21_X1 i_1_737_2037 (.A(n_1_737_1918), .B1(in_data[8]), .B2(n_1_737_1924), 
      .ZN(n_1_737_1917));
   OAI221_X1 i_1_737_2038 (.A(n_1_737_1924), .B1(n_1_737_5597), .B2(n_1_737_4855), 
      .C1(n_1_737_4856), .C2(n_1_737_1919), .ZN(n_1_737_1918));
   INV_X1 i_1_737_2039 (.A(n_1_737_1920), .ZN(n_1_737_1919));
   OAI21_X1 i_1_737_2040 (.A(n_1_737_1921), .B1(n_1_737_5598), .B2(n_1_737_4825), 
      .ZN(n_1_737_1920));
   OAI21_X1 i_1_737_2041 (.A(n_1_737_4825), .B1(n_1_737_1923), .B2(n_1_737_1922), 
      .ZN(n_1_737_1921));
   AND2_X1 i_1_737_2042 (.A1(in_data[20]), .A2(n_1_737_4846), .ZN(n_1_737_1922));
   AOI221_X1 i_1_737_2043 (.A(n_1_737_4846), .B1(n_1_737_5600), .B2(n_1_737_4837), 
      .C1(n_1_737_5601), .C2(n_1_737_4836), .ZN(n_1_737_1923));
   AOI21_X1 i_1_737_2044 (.A(n_633), .B1(n_1_737_5602), .B2(n_634), .ZN(
      n_1_737_1924));
   INV_X1 i_1_737_2045 (.A(n_1_737_1925), .ZN(n_121));
   OAI21_X1 i_1_737_2046 (.A(n_1_737_1926), .B1(in_data[8]), .B2(n_1_737_1930), 
      .ZN(n_1_737_1925));
   OAI211_X1 i_1_737_2047 (.A(n_1_737_1930), .B(n_1_737_1927), .C1(n_1_737_5597), 
      .C2(n_1_737_4870), .ZN(n_1_737_1926));
   OAI211_X1 i_1_737_2048 (.A(n_1_737_4870), .B(n_1_737_1928), .C1(in_data[16]), 
      .C2(n_1_737_4867), .ZN(n_1_737_1927));
   OAI211_X1 i_1_737_2049 (.A(n_1_737_4867), .B(n_1_737_1929), .C1(n_1_737_5599), 
      .C2(n_1_737_4877), .ZN(n_1_737_1928));
   OAI221_X1 i_1_737_2050 (.A(n_1_737_4877), .B1(in_data[24]), .B2(n_1_737_4874), 
      .C1(in_data[28]), .C2(n_1_737_4873), .ZN(n_1_737_1929));
   AOI21_X1 i_1_737_2051 (.A(n_637), .B1(n_1_737_5602), .B2(n_638), .ZN(
      n_1_737_1930));
   OAI21_X1 i_1_737_2052 (.A(n_1_737_1931), .B1(n_1_737_5596), .B2(n_1_737_1935), 
      .ZN(n_122));
   OAI211_X1 i_1_737_2053 (.A(n_1_737_1932), .B(n_1_737_1935), .C1(in_data[12]), 
      .C2(n_1_737_4907), .ZN(n_1_737_1931));
   OAI211_X1 i_1_737_2054 (.A(n_1_737_4907), .B(n_1_737_1933), .C1(n_1_737_5598), 
      .C2(n_1_737_4891), .ZN(n_1_737_1932));
   OAI211_X1 i_1_737_2055 (.A(n_1_737_1934), .B(n_1_737_4891), .C1(in_data[20]), 
      .C2(n_1_737_4897), .ZN(n_1_737_1933));
   OAI221_X1 i_1_737_2056 (.A(n_1_737_4897), .B1(n_1_737_5601), .B2(n_1_737_4886), 
      .C1(n_1_737_5600), .C2(n_1_737_4885), .ZN(n_1_737_1934));
   AOI21_X1 i_1_737_2057 (.A(n_640), .B1(n_1_737_5602), .B2(n_641), .ZN(
      n_1_737_1935));
   OAI21_X1 i_1_737_2058 (.A(n_1_737_1936), .B1(n_1_737_5596), .B2(n_1_737_1937), 
      .ZN(n_123));
   OAI211_X1 i_1_737_2059 (.A(n_1_737_1937), .B(n_1_737_1938), .C1(in_data[12]), 
      .C2(n_1_737_4956), .ZN(n_1_737_1936));
   AOI21_X1 i_1_737_2060 (.A(n_645), .B1(n_1_737_5602), .B2(n_646), .ZN(
      n_1_737_1937));
   OAI211_X1 i_1_737_2061 (.A(n_1_737_1939), .B(n_1_737_4956), .C1(n_1_737_5598), 
      .C2(n_1_737_4934), .ZN(n_1_737_1938));
   OAI211_X1 i_1_737_2062 (.A(n_1_737_1940), .B(n_1_737_4934), .C1(in_data[20]), 
      .C2(n_1_737_4949), .ZN(n_1_737_1939));
   OAI221_X1 i_1_737_2063 (.A(n_1_737_4949), .B1(n_1_737_5601), .B2(n_1_737_4928), 
      .C1(n_1_737_5600), .C2(n_1_737_4927), .ZN(n_1_737_1940));
   INV_X1 i_1_737_2064 (.A(n_1_737_1941), .ZN(n_124));
   OAI21_X1 i_1_737_2065 (.A(n_1_737_1942), .B1(in_data[8]), .B2(n_1_737_1946), 
      .ZN(n_1_737_1941));
   OAI221_X1 i_1_737_2066 (.A(n_1_737_1946), .B1(n_1_737_5597), .B2(n_1_737_4995), 
      .C1(n_1_737_4994), .C2(n_1_737_1943), .ZN(n_1_737_1942));
   AOI22_X1 i_1_737_2067 (.A1(n_1_737_4974), .A2(n_1_737_1944), .B1(in_data[16]), 
      .B2(n_1_737_4973), .ZN(n_1_737_1943));
   OAI21_X1 i_1_737_2068 (.A(n_1_737_1945), .B1(n_1_737_5599), .B2(n_1_737_4981), 
      .ZN(n_1_737_1944));
   OAI221_X1 i_1_737_2069 (.A(n_1_737_4981), .B1(in_data[28]), .B2(n_1_737_4968), 
      .C1(in_data[24]), .C2(n_1_737_4967), .ZN(n_1_737_1945));
   AOI21_X1 i_1_737_2070 (.A(n_649), .B1(n_1_737_5602), .B2(n_650), .ZN(
      n_1_737_1946));
   OAI22_X1 i_1_737_2071 (.A1(n_1_737_1949), .A2(n_1_737_1947), .B1(n_1_737_5596), 
      .B2(n_1_737_1948), .ZN(n_125));
   OAI21_X1 i_1_737_2072 (.A(n_1_737_1948), .B1(in_data[12]), .B2(n_1_737_5017), 
      .ZN(n_1_737_1947));
   AOI21_X1 i_1_737_2073 (.A(n_653), .B1(n_1_737_5602), .B2(n_654), .ZN(
      n_1_737_1948));
   AND2_X1 i_1_737_2074 (.A1(n_1_737_5017), .A2(n_1_737_1950), .ZN(n_1_737_1949));
   OAI21_X1 i_1_737_2075 (.A(n_1_737_1951), .B1(in_data[16]), .B2(n_1_737_5007), 
      .ZN(n_1_737_1950));
   OAI211_X1 i_1_737_2076 (.A(n_1_737_5007), .B(n_1_737_1952), .C1(n_1_737_5599), 
      .C2(n_1_737_5010), .ZN(n_1_737_1951));
   OAI221_X1 i_1_737_2077 (.A(n_1_737_5010), .B1(in_data[28]), .B2(n_1_737_5003), 
      .C1(in_data[24]), .C2(n_1_737_5004), .ZN(n_1_737_1952));
   OAI21_X1 i_1_737_2078 (.A(n_1_737_1953), .B1(n_1_737_5596), .B2(n_1_737_1954), 
      .ZN(n_126));
   OAI211_X1 i_1_737_2079 (.A(n_1_737_1954), .B(n_1_737_1955), .C1(in_data[12]), 
      .C2(n_1_737_5058), .ZN(n_1_737_1953));
   AOI21_X1 i_1_737_2080 (.A(n_656), .B1(n_1_737_5602), .B2(n_657), .ZN(
      n_1_737_1954));
   OAI211_X1 i_1_737_2081 (.A(n_1_737_1956), .B(n_1_737_5058), .C1(n_1_737_5598), 
      .C2(n_1_737_5031), .ZN(n_1_737_1955));
   OAI211_X1 i_1_737_2082 (.A(n_1_737_1957), .B(n_1_737_5031), .C1(in_data[20]), 
      .C2(n_1_737_5049), .ZN(n_1_737_1956));
   OAI221_X1 i_1_737_2083 (.A(n_1_737_5049), .B1(n_1_737_5601), .B2(n_1_737_5042), 
      .C1(n_1_737_5600), .C2(n_1_737_5041), .ZN(n_1_737_1957));
   OAI21_X1 i_1_737_2084 (.A(n_1_737_1958), .B1(n_1_737_5596), .B2(n_1_737_1959), 
      .ZN(n_127));
   OAI211_X1 i_1_737_2085 (.A(n_1_737_1959), .B(n_1_737_1960), .C1(in_data[12]), 
      .C2(n_1_737_5125), .ZN(n_1_737_1958));
   AOI21_X1 i_1_737_2086 (.A(n_661), .B1(n_1_737_5602), .B2(n_662), .ZN(
      n_1_737_1959));
   OAI211_X1 i_1_737_2087 (.A(n_1_737_1961), .B(n_1_737_5125), .C1(n_1_737_5598), 
      .C2(n_1_737_5114), .ZN(n_1_737_1960));
   OAI211_X1 i_1_737_2088 (.A(n_1_737_1962), .B(n_1_737_5114), .C1(in_data[20]), 
      .C2(n_1_737_5090), .ZN(n_1_737_1961));
   OAI221_X1 i_1_737_2089 (.A(n_1_737_5090), .B1(n_1_737_5601), .B2(n_1_737_5102), 
      .C1(n_1_737_5600), .C2(n_1_737_5103), .ZN(n_1_737_1962));
   OAI21_X1 i_1_737_2090 (.A(n_1_737_1963), .B1(n_1_737_5596), .B2(n_1_737_1968), 
      .ZN(n_128));
   NAND2_X1 i_1_737_2091 (.A1(n_1_737_1968), .A2(n_1_737_1964), .ZN(n_1_737_1963));
   OAI22_X1 i_1_737_2092 (.A1(n_1_737_5363), .A2(n_1_737_1965), .B1(n_1_737_5597), 
      .B2(n_1_737_5362), .ZN(n_1_737_1964));
   AOI22_X1 i_1_737_2093 (.A1(n_1_737_5186), .A2(n_1_737_1966), .B1(in_data[16]), 
      .B2(n_1_737_5187), .ZN(n_1_737_1965));
   OAI21_X1 i_1_737_2094 (.A(n_1_737_1967), .B1(n_1_737_5599), .B2(n_1_737_5233), 
      .ZN(n_1_737_1966));
   OAI221_X1 i_1_737_2095 (.A(n_1_737_5233), .B1(in_data[28]), .B2(n_1_737_5280), 
      .C1(in_data[24]), .C2(n_1_737_5279), .ZN(n_1_737_1967));
   AOI21_X1 i_1_737_2096 (.A(n_743), .B1(n_1_737_5602), .B2(n_744), .ZN(
      n_1_737_1968));
   NOR2_X1 i_1_737_2097 (.A1(n_1_737_3943), .A2(n_1_737_2057), .ZN(n_129));
   OAI21_X1 i_1_737_2102 (.A(n_1_737_5298), .B1(n_1_737_5299), .B2(n_1_737_3155), 
      .ZN(n_1_737_1972));
   OAI21_X1 i_1_737_2104 (.A(n_1_737_5366), .B1(n_1_737_5367), .B2(n_1_737_3169), 
      .ZN(n_1_737_1974));
   INV_X1 i_1_737_2105 (.A(n_1_737_1976), .ZN(n_1_737_1975));
   INV_X1 i_1_737_2107 (.A(n_1_737_1978), .ZN(n_1_737_1977));
   NOR2_X1 i_1_737_2110 (.A1(\out_as[6] [6]), .A2(n_1_737_1980), .ZN(n_130));
   OR2_X1 i_1_737_2111 (.A1(n_1_737_5067), .A2(n_1_737_1984), .ZN(n_1_737_1980));
   OR2_X1 i_1_737_2112 (.A1(n_1_737_5148), .A2(n_1_737_1984), .ZN(n_1_737_1981));
   OR2_X1 i_1_737_2113 (.A1(n_1_737_5150), .A2(n_1_737_1984), .ZN(n_1_737_1982));
   OR2_X1 i_1_737_2114 (.A1(\out_as[6] [2]), .A2(n_1_737_1984), .ZN(n_1_737_1983));
   OR2_X1 i_1_737_2115 (.A1(\out_as[6] [1]), .A2(\out_as[6] [0]), .ZN(
      n_1_737_1984));
   NAND3_X1 i_1_737_2116 (.A1(n_1_737_2014), .A2(n_1_737_2003), .A3(n_1_737_1985), 
      .ZN(n_131));
   NOR3_X1 i_1_737_2117 (.A1(n_1_737_1993), .A2(n_1_737_1987), .A3(n_1_737_1998), 
      .ZN(n_1_737_1985));
   INV_X1 i_1_737_2118 (.A(n_1_737_1987), .ZN(n_1_737_1986));
   OAI21_X1 i_1_737_2119 (.A(n_1_737_5236), .B1(n_1_737_5274), .B2(n_1_737_1988), 
      .ZN(n_1_737_1987));
   OR2_X1 i_1_737_2120 (.A1(\out_as[2] [4]), .A2(n_1_737_1989), .ZN(n_1_737_1988));
   OR2_X1 i_1_737_2121 (.A1(\out_as[2] [3]), .A2(n_1_737_1990), .ZN(n_1_737_1989));
   OR2_X1 i_1_737_2122 (.A1(\out_as[2] [2]), .A2(n_1_737_1991), .ZN(n_1_737_1990));
   OR2_X1 i_1_737_2123 (.A1(\out_as[2] [1]), .A2(\out_as[2] [0]), .ZN(
      n_1_737_1991));
   INV_X1 i_1_737_2124 (.A(n_1_737_1993), .ZN(n_1_737_1992));
   OAI21_X1 i_1_737_2125 (.A(n_1_737_5298), .B1(n_1_737_5320), .B2(n_1_737_1994), 
      .ZN(n_1_737_1993));
   OR2_X1 i_1_737_2126 (.A1(\out_as[1] [4]), .A2(n_1_737_1995), .ZN(n_1_737_1994));
   OR2_X1 i_1_737_2127 (.A1(\out_as[1] [3]), .A2(n_1_737_1996), .ZN(n_1_737_1995));
   OR2_X1 i_1_737_2128 (.A1(\out_as[1] [2]), .A2(n_1_737_1997), .ZN(n_1_737_1996));
   NAND2_X1 i_1_737_2129 (.A1(n_1_737_5653), .A2(n_1_737_5652), .ZN(n_1_737_1997));
   OAI21_X1 i_1_737_2130 (.A(n_1_737_5366), .B1(n_1_737_5386), .B2(n_1_737_1999), 
      .ZN(n_1_737_1998));
   OR2_X1 i_1_737_2131 (.A1(\out_as[4] [4]), .A2(n_1_737_2000), .ZN(n_1_737_1999));
   OR2_X1 i_1_737_2132 (.A1(\out_as[4] [3]), .A2(n_1_737_2001), .ZN(n_1_737_2000));
   OR2_X1 i_1_737_2133 (.A1(\out_as[4] [2]), .A2(n_1_737_2002), .ZN(n_1_737_2001));
   NAND2_X1 i_1_737_2134 (.A1(n_1_737_5614), .A2(n_1_737_5613), .ZN(n_1_737_2002));
   NOR3_X1 i_1_737_2135 (.A1(n_1_737_2009), .A2(n_1_737_2004), .A3(n_1_737_5336), 
      .ZN(n_1_737_2003));
   NOR2_X1 i_1_737_2136 (.A1(n_1_737_5358), .A2(n_1_737_2005), .ZN(n_1_737_2004));
   OR2_X1 i_1_737_2137 (.A1(\out_as[0] [4]), .A2(n_1_737_2006), .ZN(n_1_737_2005));
   OR2_X1 i_1_737_2138 (.A1(\out_as[0] [3]), .A2(n_1_737_2007), .ZN(n_1_737_2006));
   OR2_X1 i_1_737_2139 (.A1(\out_as[0] [2]), .A2(n_1_737_2008), .ZN(n_1_737_2007));
   NAND2_X1 i_1_737_2140 (.A1(n_1_737_5673), .A2(n_1_737_5672), .ZN(n_1_737_2008));
   OAI21_X1 i_1_737_2141 (.A(n_1089), .B1(n_1_737_5167), .B2(n_1_737_2010), 
      .ZN(n_1_737_2009));
   OR2_X1 i_1_737_2142 (.A1(n_1_737_5160), .A2(n_1_737_2013), .ZN(n_1_737_2010));
   OR2_X1 i_1_737_2143 (.A1(n_1_737_5162), .A2(n_1_737_2013), .ZN(n_1_737_2011));
   OR2_X1 i_1_737_2144 (.A1(\out_as[5] [2]), .A2(n_1_737_2013), .ZN(n_1_737_2012));
   OR2_X1 i_1_737_2145 (.A1(\out_as[5] [1]), .A2(\out_as[5] [0]), .ZN(
      n_1_737_2013));
   INV_X1 i_1_737_2146 (.A(n_1_737_2015), .ZN(n_1_737_2014));
   OAI21_X1 i_1_737_2147 (.A(n_1_737_5190), .B1(n_1_737_5215), .B2(n_1_737_2016), 
      .ZN(n_1_737_2015));
   OR2_X1 i_1_737_2148 (.A1(\out_as[3] [4]), .A2(n_1_737_2017), .ZN(n_1_737_2016));
   OR2_X1 i_1_737_2149 (.A1(\out_as[3] [3]), .A2(n_1_737_2018), .ZN(n_1_737_2017));
   OR2_X1 i_1_737_2150 (.A1(\out_as[3] [2]), .A2(n_1_737_2019), .ZN(n_1_737_2018));
   OR2_X1 i_1_737_2151 (.A1(\out_as[3] [1]), .A2(\out_as[3] [0]), .ZN(
      n_1_737_2019));
   NOR2_X1 i_1_737_2152 (.A1(n_1_737_5140), .A2(n_1_737_2020), .ZN(n_132));
   OR2_X1 i_1_737_2153 (.A1(n_1_737_5143), .A2(n_1_737_2023), .ZN(n_1_737_2020));
   OR2_X1 i_1_737_2154 (.A1(n_1_737_5145), .A2(n_1_737_2023), .ZN(n_1_737_2021));
   OR2_X1 i_1_737_2155 (.A1(\out_as[7] [2]), .A2(n_1_737_2023), .ZN(n_1_737_2022));
   OR2_X1 i_1_737_2156 (.A1(\out_as[7] [1]), .A2(\out_as[7] [0]), .ZN(
      n_1_737_2023));
   OR2_X1 i_1_737_2157 (.A1(\out_as[7] [3]), .A2(n_1_737_2025), .ZN(n_1_737_2024));
   OR2_X1 i_1_737_2158 (.A1(\out_as[7] [2]), .A2(\out_as[7] [1]), .ZN(
      n_1_737_2025));
   NOR2_X1 i_1_737_2159 (.A1(n_1_737_958), .A2(n_1_737_2026), .ZN(n_133));
   NAND2_X1 i_1_737_2160 (.A1(n_1_737_958), .A2(n_1_737_2026), .ZN(n_134));
   NAND3_X1 i_1_737_2161 (.A1(n_1311), .A2(n_1_737_3222), .A3(\out_bs[6] [6]), 
      .ZN(n_1_737_2026));
   NOR3_X1 i_1_737_2162 (.A1(n_1_737_4119), .A2(n_1_737_3109), .A3(n_1_737_957), 
      .ZN(n_135));
   OAI21_X1 i_1_737_2163 (.A(n_1_737_957), .B1(n_1_737_4119), .B2(n_1_737_3109), 
      .ZN(n_136));
   OAI211_X1 i_1_737_2164 (.A(n_1_737_2040), .B(n_1_737_2027), .C1(n_1_737_952), 
      .C2(n_1_737_2042), .ZN(n_137));
   NOR4_X1 i_1_737_2165 (.A1(n_1_737_2031), .A2(n_1_737_2028), .A3(n_1_737_2034), 
      .A4(n_1_737_2037), .ZN(n_1_737_2027));
   INV_X1 i_1_737_2166 (.A(n_1_737_2029), .ZN(n_1_737_2028));
   OAI21_X1 i_1_737_2167 (.A(n_1_737_2030), .B1(n_1_737_5407), .B2(n_1_737_5297), 
      .ZN(n_1_737_2029));
   OAI22_X1 i_1_737_2168 (.A1(n_1_737_4653), .A2(n_1_737_2312), .B1(n_1_737_953), 
      .B2(n_1_737_5298), .ZN(n_1_737_2030));
   AOI21_X1 i_1_737_2169 (.A(n_1_737_2032), .B1(n_1_737_955), .B2(n_1_737_5190), 
      .ZN(n_1_737_2031));
   INV_X1 i_1_737_2170 (.A(n_1_737_2033), .ZN(n_1_737_2032));
   OAI22_X1 i_1_737_2171 (.A1(n_1_737_4658), .A2(n_1_737_2303), .B1(n_1_737_955), 
      .B2(n_1_737_5190), .ZN(n_1_737_2033));
   INV_X1 i_1_737_2172 (.A(n_1_737_2035), .ZN(n_1_737_2034));
   OAI21_X1 i_1_737_2173 (.A(n_1_737_2036), .B1(n_1_737_5406), .B2(n_1_737_5235), 
      .ZN(n_1_737_2035));
   OAI22_X1 i_1_737_2174 (.A1(n_1_737_4664), .A2(n_1_737_2307), .B1(n_1_737_954), 
      .B2(n_1_737_5236), .ZN(n_1_737_2036));
   AOI21_X1 i_1_737_2175 (.A(n_1_737_2038), .B1(n_1_737_956), .B2(n_1_737_5366), 
      .ZN(n_1_737_2037));
   INV_X1 i_1_737_2176 (.A(n_1_737_2039), .ZN(n_1_737_2038));
   OAI22_X1 i_1_737_2177 (.A1(n_1_737_4676), .A2(n_1_737_2320), .B1(n_1_737_956), 
      .B2(n_1_737_5366), .ZN(n_1_737_2039));
   INV_X1 i_1_737_2178 (.A(n_1_737_2041), .ZN(n_1_737_2040));
   AOI21_X1 i_1_737_2179 (.A(n_1_737_5337), .B1(n_1_737_952), .B2(n_1_737_2042), 
      .ZN(n_1_737_2041));
   NAND3_X1 i_1_737_2180 (.A1(\out_bs[0] [5]), .A2(n_1_737_4138), .A3(
      \out_bs[0] [6]), .ZN(n_1_737_2042));
   AND2_X1 i_1_737_2181 (.A1(n_1272), .A2(n_746), .ZN(n_138));
   NOR3_X1 i_1_737_2182 (.A1(n_1_737_4964), .A2(n_1_737_2171), .A3(n_1_737_950), 
      .ZN(n_139));
   OAI21_X1 i_1_737_2183 (.A(n_1_737_950), .B1(n_1_737_4964), .B2(n_1_737_2171), 
      .ZN(n_140));
   NAND4_X1 i_1_737_2184 (.A1(n_1_737_2045), .A2(n_1_737_2043), .A3(n_1_737_2047), 
      .A4(n_1_737_2055), .ZN(n_141));
   OAI21_X1 i_1_737_2185 (.A(n_1_737_5411), .B1(n_1_737_5336), .B2(n_1_737_2048), 
      .ZN(n_1_737_2043));
   INV_X1 i_1_737_2186 (.A(n_1_737_2045), .ZN(n_1_737_2044));
   OAI21_X1 i_1_737_2187 (.A(n_1_737_2046), .B1(n_1_737_5409), .B2(n_1_737_5235), 
      .ZN(n_1_737_2045));
   OAI22_X1 i_1_737_2188 (.A1(n_1_737_4706), .A2(n_1_737_2307), .B1(n_1_737_947), 
      .B2(n_1_737_5236), .ZN(n_1_737_2046));
   AOI211_X1 i_1_737_2189 (.A(n_1_737_2049), .B(n_1_737_2052), .C1(n_1_737_5336), 
      .C2(n_1_737_2048), .ZN(n_1_737_2047));
   NOR2_X1 i_1_737_2190 (.A1(n_1_737_4685), .A2(n_1_737_2315), .ZN(n_1_737_2048));
   INV_X1 i_1_737_2191 (.A(n_1_737_2050), .ZN(n_1_737_2049));
   OAI21_X1 i_1_737_2192 (.A(n_1_737_2051), .B1(n_1_737_5410), .B2(n_1_737_5297), 
      .ZN(n_1_737_2050));
   OAI22_X1 i_1_737_2193 (.A1(n_1_737_4698), .A2(n_1_737_2312), .B1(n_1_737_946), 
      .B2(n_1_737_5298), .ZN(n_1_737_2051));
   AOI21_X1 i_1_737_2194 (.A(n_1_737_2053), .B1(n_1_737_948), .B2(n_1_737_5190), 
      .ZN(n_1_737_2052));
   INV_X1 i_1_737_2195 (.A(n_1_737_2054), .ZN(n_1_737_2053));
   OAI22_X1 i_1_737_2196 (.A1(n_1_737_4691), .A2(n_1_737_2303), .B1(n_1_737_948), 
      .B2(n_1_737_5190), .ZN(n_1_737_2054));
   OAI21_X1 i_1_737_2197 (.A(n_1_737_2056), .B1(n_1_737_5408), .B2(n_1_737_5365), 
      .ZN(n_1_737_2055));
   OAI22_X1 i_1_737_2198 (.A1(n_1_737_4714), .A2(n_1_737_2320), .B1(n_1_737_949), 
      .B2(n_1_737_5366), .ZN(n_1_737_2056));
   NOR2_X1 i_1_737_2199 (.A1(n_1_737_944), .A2(n_1_737_2057), .ZN(n_142));
   NAND2_X1 i_1_737_2200 (.A1(n_1_737_944), .A2(n_1_737_2057), .ZN(n_143));
   NAND2_X1 i_1_737_2201 (.A1(\out_bs[6] [6]), .A2(n_1_737_3222), .ZN(
      n_1_737_2057));
   NOR2_X1 i_1_737_2202 (.A1(n_1_737_943), .A2(n_1_737_2058), .ZN(n_144));
   NAND2_X1 i_1_737_2203 (.A1(n_1_737_943), .A2(n_1_737_2058), .ZN(n_145));
   NAND3_X1 i_1_737_2204 (.A1(n_845), .A2(n_1_737_4209), .A3(n_844), .ZN(
      n_1_737_2058));
   OAI211_X1 i_1_737_2205 (.A(n_1_737_2073), .B(n_1_737_2059), .C1(n_1_737_938), 
      .C2(n_1_737_2075), .ZN(n_146));
   NOR4_X1 i_1_737_2206 (.A1(n_1_737_2063), .A2(n_1_737_2060), .A3(n_1_737_2066), 
      .A4(n_1_737_2069), .ZN(n_1_737_2059));
   INV_X1 i_1_737_2207 (.A(n_1_737_2061), .ZN(n_1_737_2060));
   OAI21_X1 i_1_737_2208 (.A(n_1_737_2062), .B1(n_1_737_5413), .B2(n_1_737_5297), 
      .ZN(n_1_737_2061));
   OAI22_X1 i_1_737_2209 (.A1(n_1_737_4218), .A2(n_1_737_3015), .B1(n_1_737_939), 
      .B2(n_1_737_5298), .ZN(n_1_737_2062));
   AOI21_X1 i_1_737_2210 (.A(n_1_737_2064), .B1(n_1_737_941), .B2(n_1_737_5190), 
      .ZN(n_1_737_2063));
   INV_X1 i_1_737_2211 (.A(n_1_737_2065), .ZN(n_1_737_2064));
   OAI22_X1 i_1_737_2212 (.A1(n_1_737_4225), .A2(n_1_737_3005), .B1(n_1_737_941), 
      .B2(n_1_737_5190), .ZN(n_1_737_2065));
   AOI21_X1 i_1_737_2213 (.A(n_1_737_2067), .B1(n_1_737_940), .B2(n_1_737_5236), 
      .ZN(n_1_737_2066));
   INV_X1 i_1_737_2214 (.A(n_1_737_2068), .ZN(n_1_737_2067));
   OAI22_X1 i_1_737_2215 (.A1(n_1_737_4234), .A2(n_1_737_3010), .B1(n_1_737_940), 
      .B2(n_1_737_5236), .ZN(n_1_737_2068));
   INV_X1 i_1_737_2216 (.A(n_1_737_2070), .ZN(n_1_737_2069));
   OAI21_X1 i_1_737_2217 (.A(n_1_737_2071), .B1(n_1_737_5412), .B2(n_1_737_5365), 
      .ZN(n_1_737_2070));
   OAI21_X1 i_1_737_2218 (.A(n_1_737_2072), .B1(n_1_737_942), .B2(n_1_737_5366), 
      .ZN(n_1_737_2071));
   NAND2_X1 i_1_737_2219 (.A1(n_1_737_4253), .A2(n_1_737_3023), .ZN(n_1_737_2072));
   INV_X1 i_1_737_2220 (.A(n_1_737_2074), .ZN(n_1_737_2073));
   AOI21_X1 i_1_737_2221 (.A(n_1_737_5337), .B1(n_1_737_938), .B2(n_1_737_2075), 
      .ZN(n_1_737_2074));
   NAND3_X1 i_1_737_2222 (.A1(\out_bs[0] [5]), .A2(n_1_737_4243), .A3(
      \out_bs[0] [6]), .ZN(n_1_737_2075));
   NOR3_X1 i_1_737_2223 (.A1(n_1_737_4207), .A2(n_1_737_3109), .A3(n_1_737_936), 
      .ZN(n_147));
   OAI21_X1 i_1_737_2224 (.A(n_1_737_936), .B1(n_1_737_4207), .B2(n_1_737_3109), 
      .ZN(n_148));
   NAND4_X1 i_1_737_2225 (.A1(n_1_737_2078), .A2(n_1_737_2076), .A3(n_1_737_2080), 
      .A4(n_1_737_2088), .ZN(n_149));
   OAI21_X1 i_1_737_2226 (.A(n_1_737_5418), .B1(n_1_737_5336), .B2(n_1_737_2081), 
      .ZN(n_1_737_2076));
   INV_X1 i_1_737_2227 (.A(n_1_737_2078), .ZN(n_1_737_2077));
   OAI21_X1 i_1_737_2228 (.A(n_1_737_2079), .B1(n_1_737_5416), .B2(n_1_737_5235), 
      .ZN(n_1_737_2078));
   OAI22_X1 i_1_737_2229 (.A1(n_1_737_4231), .A2(n_1_737_3010), .B1(n_1_737_933), 
      .B2(n_1_737_5236), .ZN(n_1_737_2079));
   AOI211_X1 i_1_737_2230 (.A(n_1_737_2082), .B(n_1_737_2085), .C1(n_1_737_5336), 
      .C2(n_1_737_2081), .ZN(n_1_737_2080));
   NOR2_X1 i_1_737_2231 (.A1(n_1_737_4242), .A2(n_1_737_3018), .ZN(n_1_737_2081));
   INV_X1 i_1_737_2232 (.A(n_1_737_2083), .ZN(n_1_737_2082));
   OAI21_X1 i_1_737_2233 (.A(n_1_737_2084), .B1(n_1_737_5417), .B2(n_1_737_5297), 
      .ZN(n_1_737_2083));
   OAI22_X1 i_1_737_2234 (.A1(n_1_737_4216), .A2(n_1_737_3015), .B1(n_1_737_932), 
      .B2(n_1_737_5298), .ZN(n_1_737_2084));
   AOI21_X1 i_1_737_2235 (.A(n_1_737_2086), .B1(n_1_737_934), .B2(n_1_737_5190), 
      .ZN(n_1_737_2085));
   AOI22_X1 i_1_737_2236 (.A1(n_1_737_4223), .A2(n_1_737_3006), .B1(n_1_737_5415), 
      .B2(n_1_737_5189), .ZN(n_1_737_2086));
   INV_X1 i_1_737_2237 (.A(n_1_737_2088), .ZN(n_1_737_2087));
   OAI21_X1 i_1_737_2238 (.A(n_1_737_2089), .B1(n_1_737_5414), .B2(n_1_737_5365), 
      .ZN(n_1_737_2088));
   OAI22_X1 i_1_737_2239 (.A1(n_1_737_4250), .A2(n_1_737_3022), .B1(n_1_737_935), 
      .B2(n_1_737_5366), .ZN(n_1_737_2089));
   NOR3_X1 i_1_737_2240 (.A1(n_1_737_4813), .A2(n_1_737_2298), .A3(n_1_737_929), 
      .ZN(n_150));
   OAI21_X1 i_1_737_2241 (.A(n_1_737_929), .B1(n_1_737_4813), .B2(n_1_737_2298), 
      .ZN(n_151));
   OAI211_X1 i_1_737_2242 (.A(n_1_737_2102), .B(n_1_737_2090), .C1(n_1_737_924), 
      .C2(n_1_737_2104), .ZN(n_152));
   NOR4_X1 i_1_737_2243 (.A1(n_1_737_2094), .A2(n_1_737_2091), .A3(n_1_737_2097), 
      .A4(n_1_737_2100), .ZN(n_1_737_2090));
   INV_X1 i_1_737_2244 (.A(n_1_737_2092), .ZN(n_1_737_2091));
   OAI21_X1 i_1_737_2245 (.A(n_1_737_2093), .B1(n_1_737_5421), .B2(n_1_737_5297), 
      .ZN(n_1_737_2092));
   OAI22_X1 i_1_737_2246 (.A1(n_1_737_4844), .A2(n_1_737_2312), .B1(n_1_737_925), 
      .B2(n_1_737_5298), .ZN(n_1_737_2093));
   INV_X1 i_1_737_2247 (.A(n_1_737_2095), .ZN(n_1_737_2094));
   OAI21_X1 i_1_737_2248 (.A(n_1_737_2096), .B1(n_1_737_5420), .B2(n_1_737_5189), 
      .ZN(n_1_737_2095));
   OAI22_X1 i_1_737_2249 (.A1(n_1_737_4834), .A2(n_1_737_2303), .B1(n_1_737_927), 
      .B2(n_1_737_5190), .ZN(n_1_737_2096));
   AOI21_X1 i_1_737_2250 (.A(n_1_737_2098), .B1(n_1_737_926), .B2(n_1_737_5236), 
      .ZN(n_1_737_2097));
   INV_X1 i_1_737_2251 (.A(n_1_737_2099), .ZN(n_1_737_2098));
   OAI22_X1 i_1_737_2252 (.A1(n_1_737_4853), .A2(n_1_737_2307), .B1(n_1_737_926), 
      .B2(n_1_737_5236), .ZN(n_1_737_2099));
   AOI21_X1 i_1_737_2253 (.A(n_1_737_2101), .B1(n_1_737_928), .B2(n_1_737_5366), 
      .ZN(n_1_737_2100));
   AOI22_X1 i_1_737_2254 (.A1(n_1_737_4285), .A2(n_1_737_3023), .B1(n_1_737_5419), 
      .B2(n_1_737_5365), .ZN(n_1_737_2101));
   INV_X1 i_1_737_2255 (.A(n_1_737_2103), .ZN(n_1_737_2102));
   AOI21_X1 i_1_737_2256 (.A(n_1_737_5337), .B1(n_1_737_924), .B2(n_1_737_2104), 
      .ZN(n_1_737_2103));
   NAND3_X1 i_1_737_2257 (.A1(\out_bs[0] [5]), .A2(n_1_737_4266), .A3(
      \out_bs[0] [6]), .ZN(n_1_737_2104));
   NOR2_X1 i_1_737_2258 (.A1(n_1_737_923), .A2(n_1_737_2105), .ZN(n_153));
   NAND2_X1 i_1_737_2259 (.A1(n_1_737_923), .A2(n_1_737_2105), .ZN(n_154));
   NAND3_X1 i_1_737_2260 (.A1(n_1_737_4015), .A2(n_1_737_3330), .A3(
      \out_bs[6] [6]), .ZN(n_1_737_2105));
   NOR3_X1 i_1_737_2261 (.A1(n_1_737_4809), .A2(n_1_737_2298), .A3(n_1_737_922), 
      .ZN(n_155));
   OAI21_X1 i_1_737_2262 (.A(n_1_737_922), .B1(n_1_737_4809), .B2(n_1_737_2298), 
      .ZN(n_156));
   NAND4_X1 i_1_737_2263 (.A1(n_1_737_2109), .A2(n_1_737_2106), .A3(n_1_737_2114), 
      .A4(n_1_737_2116), .ZN(n_157));
   AOI21_X1 i_1_737_2264 (.A(n_1_737_2111), .B1(n_1_737_2108), .B2(n_1_737_2107), 
      .ZN(n_1_737_2106));
   NAND2_X1 i_1_737_2265 (.A1(n_1_737_917), .A2(n_1_737_5337), .ZN(n_1_737_2107));
   OAI22_X1 i_1_737_2266 (.A1(n_1_737_4820), .A2(n_1_737_2315), .B1(n_1_737_917), 
      .B2(n_1_737_5337), .ZN(n_1_737_2108));
   OAI21_X1 i_1_737_2267 (.A(n_1_737_2110), .B1(n_1_737_5424), .B2(n_1_737_5235), 
      .ZN(n_1_737_2109));
   OAI22_X1 i_1_737_2268 (.A1(n_1_737_4851), .A2(n_1_737_2307), .B1(n_1_737_919), 
      .B2(n_1_737_5236), .ZN(n_1_737_2110));
   INV_X1 i_1_737_2269 (.A(n_1_737_2112), .ZN(n_1_737_2111));
   OAI21_X1 i_1_737_2270 (.A(n_1_737_2113), .B1(n_1_737_5425), .B2(n_1_737_5297), 
      .ZN(n_1_737_2112));
   OAI22_X1 i_1_737_2271 (.A1(n_1_737_4840), .A2(n_1_737_2312), .B1(n_1_737_918), 
      .B2(n_1_737_5298), .ZN(n_1_737_2113));
   OAI21_X1 i_1_737_2272 (.A(n_1_737_2115), .B1(n_1_737_5423), .B2(n_1_737_5189), 
      .ZN(n_1_737_2114));
   OAI22_X1 i_1_737_2273 (.A1(n_1_737_4830), .A2(n_1_737_2303), .B1(n_1_737_920), 
      .B2(n_1_737_5190), .ZN(n_1_737_2115));
   OAI21_X1 i_1_737_2274 (.A(n_1_737_2117), .B1(n_1_737_5422), .B2(n_1_737_5365), 
      .ZN(n_1_737_2116));
   OAI22_X1 i_1_737_2275 (.A1(n_1_737_4861), .A2(n_1_737_2320), .B1(n_1_737_921), 
      .B2(n_1_737_5366), .ZN(n_1_737_2117));
   NOR2_X1 i_1_737_2276 (.A1(n_1_737_916), .A2(n_1_737_2118), .ZN(n_158));
   NAND2_X1 i_1_737_2277 (.A1(n_1_737_916), .A2(n_1_737_2118), .ZN(n_159));
   NAND2_X1 i_1_737_2278 (.A1(\out_bs[6] [6]), .A2(n_1_737_3330), .ZN(
      n_1_737_2118));
   NAND3_X1 i_1_737_2279 (.A1(n_1_737_2133), .A2(n_1_737_2128), .A3(n_1_737_2119), 
      .ZN(n_160));
   NOR3_X1 i_1_737_2280 (.A1(n_1_737_2123), .A2(n_1_737_2120), .A3(n_1_737_2125), 
      .ZN(n_1_737_2119));
   OAI21_X1 i_1_737_2281 (.A(n_1_737_2121), .B1(n_1_737_910), .B2(n_1_737_2190), 
      .ZN(n_1_737_2120));
   OAI21_X1 i_1_737_2282 (.A(n_1_737_2122), .B1(n_1_737_5602), .B2(n_1_737_5426), 
      .ZN(n_1_737_2121));
   OAI21_X1 i_1_737_2283 (.A(n_1_737_2171), .B1(n_1089), .B2(n_1_737_915), 
      .ZN(n_1_737_2122));
   OAI22_X1 i_1_737_2284 (.A1(n_1_737_912), .A2(n_1_737_2185), .B1(n_1_737_5236), 
      .B2(n_1_737_2124), .ZN(n_1_737_2123));
   AND2_X1 i_1_737_2285 (.A1(n_1_737_912), .A2(n_1_737_2185), .ZN(n_1_737_2124));
   INV_X1 i_1_737_2286 (.A(n_1_737_2126), .ZN(n_1_737_2125));
   OAI21_X1 i_1_737_2287 (.A(n_1_737_2127), .B1(n_1_737_5427), .B2(n_1_737_5365), 
      .ZN(n_1_737_2126));
   OAI22_X1 i_1_737_2288 (.A1(n_1_737_5625), .A2(n_1_737_3457), .B1(n_1_737_914), 
      .B2(n_1_737_5366), .ZN(n_1_737_2127));
   AOI21_X1 i_1_737_2289 (.A(n_1_737_2130), .B1(n_1_737_5336), .B2(n_1_737_2129), 
      .ZN(n_1_737_2128));
   NAND2_X1 i_1_737_2290 (.A1(n_1_737_910), .A2(n_1_737_2190), .ZN(n_1_737_2129));
   OAI22_X1 i_1_737_2291 (.A1(n_1_737_913), .A2(n_1_737_2181), .B1(n_1_737_5190), 
      .B2(n_1_737_2131), .ZN(n_1_737_2130));
   AND2_X1 i_1_737_2292 (.A1(n_1_737_913), .A2(n_1_737_2181), .ZN(n_1_737_2131));
   INV_X1 i_1_737_2293 (.A(n_1_737_2133), .ZN(n_1_737_2132));
   OAI21_X1 i_1_737_2294 (.A(n_1_737_2134), .B1(n_1_737_5297), .B2(n_1_737_2176), 
      .ZN(n_1_737_2133));
   OAI21_X1 i_1_737_2295 (.A(n_1_737_911), .B1(n_1_737_5298), .B2(n_1_737_2177), 
      .ZN(n_1_737_2134));
   NOR2_X1 i_1_737_2296 (.A1(n_1_737_908), .A2(n_1_737_2135), .ZN(n_161));
   NAND2_X1 i_1_737_2297 (.A1(n_1_737_908), .A2(n_1_737_2135), .ZN(n_162));
   OAI21_X1 i_1_737_2298 (.A(n_1_737_2299), .B1(n_846), .B2(n_1_737_4883), 
      .ZN(n_1_737_2135));
   OR3_X1 i_1_737_2299 (.A1(n_1_737_2150), .A2(n_1_737_2136), .A3(n_1_737_2142), 
      .ZN(n_163));
   NAND2_X1 i_1_737_2300 (.A1(n_1_737_2140), .A2(n_1_737_2137), .ZN(n_1_737_2136));
   OAI21_X1 i_1_737_2301 (.A(n_1_737_2138), .B1(n_1_737_5429), .B2(n_1_737_5189), 
      .ZN(n_1_737_2137));
   OAI22_X1 i_1_737_2302 (.A1(n_1_737_5638), .A2(n_1_737_3363), .B1(n_1_737_906), 
      .B2(n_1_737_5190), .ZN(n_1_737_2138));
   INV_X1 i_1_737_2303 (.A(n_1_737_2140), .ZN(n_1_737_2139));
   OAI21_X1 i_1_737_2304 (.A(n_1_737_2141), .B1(n_1_737_5428), .B2(n_1_737_5365), 
      .ZN(n_1_737_2140));
   OAI22_X1 i_1_737_2305 (.A1(n_1_737_5625), .A2(n_1_737_3382), .B1(n_1_737_907), 
      .B2(n_1_737_5366), .ZN(n_1_737_2141));
   OAI221_X1 i_1_737_2306 (.A(n_1_737_2143), .B1(n_1_737_5337), .B2(n_1_737_2148), 
      .C1(n_1_737_903), .C2(n_1_737_2147), .ZN(n_1_737_2142));
   INV_X1 i_1_737_2307 (.A(n_1_737_2144), .ZN(n_1_737_2143));
   OAI22_X1 i_1_737_2308 (.A1(n_1_737_904), .A2(n_1_737_5298), .B1(n_1_737_2146), 
      .B2(n_1_737_2145), .ZN(n_1_737_2144));
   AOI21_X1 i_1_737_2309 (.A(n_1_737_2176), .B1(n_1_737_4890), .B2(n_1_737_2313), 
      .ZN(n_1_737_2145));
   AND2_X1 i_1_737_2310 (.A1(n_1_737_904), .A2(n_1_737_5298), .ZN(n_1_737_2146));
   NOR2_X1 i_1_737_2311 (.A1(n_1_737_5336), .A2(n_1_737_2149), .ZN(n_1_737_2147));
   INV_X1 i_1_737_2312 (.A(n_1_737_2149), .ZN(n_1_737_2148));
   NOR2_X1 i_1_737_2313 (.A1(n_1_737_5671), .A2(n_1_737_3357), .ZN(n_1_737_2149));
   INV_X1 i_1_737_2314 (.A(n_1_737_2151), .ZN(n_1_737_2150));
   OAI21_X1 i_1_737_2315 (.A(n_1_737_2152), .B1(n_1_737_5430), .B2(n_1_737_5235), 
      .ZN(n_1_737_2151));
   OAI22_X1 i_1_737_2316 (.A1(n_1_737_5651), .A2(n_1_737_3374), .B1(n_1_737_905), 
      .B2(n_1_737_5236), .ZN(n_1_737_2152));
   NOR2_X1 i_1_737_2317 (.A1(n_1_737_902), .A2(n_1_737_2153), .ZN(n_164));
   NAND2_X1 i_1_737_2318 (.A1(n_1_737_902), .A2(n_1_737_2153), .ZN(n_165));
   OAI21_X1 i_1_737_2319 (.A(n_1_737_2253), .B1(n_847), .B2(n_1_737_4921), 
      .ZN(n_1_737_2153));
   NOR2_X1 i_1_737_2320 (.A1(n_1_737_901), .A2(n_1_737_2154), .ZN(n_166));
   NAND2_X1 i_1_737_2321 (.A1(n_1_737_901), .A2(n_1_737_2154), .ZN(n_167));
   AOI22_X1 i_1_737_2322 (.A1(n_1_737_4404), .A2(n_1_737_3110), .B1(n_844), 
      .B2(n_1_737_3386), .ZN(n_1_737_2154));
   NAND3_X1 i_1_737_2323 (.A1(n_1_737_2157), .A2(n_1_737_2155), .A3(n_1_737_2167), 
      .ZN(n_168));
   AOI211_X1 i_1_737_2324 (.A(n_1_737_2164), .B(n_1_737_2159), .C1(n_1_737_2163), 
      .C2(n_1_737_2162), .ZN(n_1_737_2155));
   INV_X1 i_1_737_2325 (.A(n_1_737_2157), .ZN(n_1_737_2156));
   OAI21_X1 i_1_737_2326 (.A(n_1_737_2158), .B1(n_1_737_5432), .B2(n_1_737_5189), 
      .ZN(n_1_737_2157));
   OAI22_X1 i_1_737_2327 (.A1(n_1_737_5638), .A2(n_1_737_5679), .B1(n_1_737_899), 
      .B2(n_1_737_5190), .ZN(n_1_737_2158));
   AOI21_X1 i_1_737_2328 (.A(n_1_737_2160), .B1(n_1_737_898), .B2(n_1_737_5236), 
      .ZN(n_1_737_2159));
   INV_X1 i_1_737_2329 (.A(n_1_737_2161), .ZN(n_1_737_2160));
   OAI22_X1 i_1_737_2330 (.A1(n_1_737_5651), .A2(n_1_737_5680), .B1(n_1_737_898), 
      .B2(n_1_737_5236), .ZN(n_1_737_2161));
   NAND2_X1 i_1_737_2331 (.A1(n_1_737_896), .A2(n_1_737_5337), .ZN(n_1_737_2162));
   OAI22_X1 i_1_737_2332 (.A1(n_1_737_5671), .A2(n_1_737_3403), .B1(n_1_737_896), 
      .B2(n_1_737_5337), .ZN(n_1_737_2163));
   INV_X1 i_1_737_2333 (.A(n_1_737_2165), .ZN(n_1_737_2164));
   OAI21_X1 i_1_737_2334 (.A(n_1_737_2166), .B1(n_1_737_5433), .B2(n_1_737_5297), 
      .ZN(n_1_737_2165));
   OAI22_X1 i_1_737_2335 (.A1(n_1_737_897), .A2(n_1_737_5298), .B1(n_1_737_5664), 
      .B2(n_1_737_3410), .ZN(n_1_737_2166));
   OAI21_X1 i_1_737_2336 (.A(n_1_737_2168), .B1(n_1_737_5431), .B2(n_1_737_5365), 
      .ZN(n_1_737_2167));
   OAI22_X1 i_1_737_2337 (.A1(n_1_737_5625), .A2(n_1_737_3417), .B1(n_1_737_900), 
      .B2(n_1_737_5366), .ZN(n_1_737_2168));
   NOR2_X1 i_1_737_2338 (.A1(n_1_737_895), .A2(n_1_737_2169), .ZN(n_169));
   NAND2_X1 i_1_737_2339 (.A1(n_1_737_895), .A2(n_1_737_2169), .ZN(n_170));
   OAI21_X1 i_1_737_2340 (.A(n_1_737_2253), .B1(n_847), .B2(n_1_737_3883), 
      .ZN(n_1_737_2169));
   NOR2_X1 i_1_737_2341 (.A1(n_1_737_894), .A2(n_1_737_2170), .ZN(n_171));
   NAND2_X1 i_1_737_2342 (.A1(n_1_737_894), .A2(n_1_737_2170), .ZN(n_172));
   OAI21_X1 i_1_737_2343 (.A(n_1_737_2299), .B1(n_846), .B2(n_1_737_4965), 
      .ZN(n_1_737_2170));
   NAND2_X1 i_1_737_2344 (.A1(n_1_737_4404), .A2(n_1_737_3110), .ZN(n_1_737_2171));
   NAND3_X1 i_1_737_2345 (.A1(n_1_737_2186), .A2(n_1_737_2172), .A3(n_1_737_2188), 
      .ZN(n_173));
   NOR3_X1 i_1_737_2346 (.A1(n_1_737_2178), .A2(n_1_737_2173), .A3(n_1_737_2183), 
      .ZN(n_1_737_2172));
   INV_X1 i_1_737_2347 (.A(n_1_737_2174), .ZN(n_1_737_2173));
   OAI21_X1 i_1_737_2348 (.A(n_1_737_2175), .B1(n_1_737_5437), .B2(n_1_737_5297), 
      .ZN(n_1_737_2174));
   OAI221_X1 i_1_737_2349 (.A(n_1_737_2177), .B1(n_1_737_5664), .B2(n_1_737_3438), 
      .C1(n_1_737_890), .C2(n_1_737_5298), .ZN(n_1_737_2175));
   INV_X1 i_1_737_2350 (.A(n_1_737_2177), .ZN(n_1_737_2176));
   NAND2_X1 i_1_737_2351 (.A1(\out_bs[1] [6]), .A2(n_1_737_3440), .ZN(
      n_1_737_2177));
   INV_X1 i_1_737_2352 (.A(n_1_737_2179), .ZN(n_1_737_2178));
   OAI21_X1 i_1_737_2353 (.A(n_1_737_2180), .B1(n_1_737_5435), .B2(n_1_737_5189), 
      .ZN(n_1_737_2179));
   OAI221_X1 i_1_737_2354 (.A(n_1_737_2181), .B1(n_1_737_4979), .B2(n_1_737_2303), 
      .C1(n_1_737_892), .C2(n_1_737_5190), .ZN(n_1_737_2180));
   NAND2_X1 i_1_737_2355 (.A1(n_1_737_4427), .A2(n_1_737_3006), .ZN(n_1_737_2181));
   INV_X1 i_1_737_2356 (.A(n_1_737_2183), .ZN(n_1_737_2182));
   AOI21_X1 i_1_737_2357 (.A(n_1_737_2184), .B1(n_1_737_891), .B2(n_1_737_5236), 
      .ZN(n_1_737_2183));
   AOI22_X1 i_1_737_2358 (.A1(\out_bs[2] [6]), .A2(n_1_737_3445), .B1(
      n_1_737_5436), .B2(n_1_737_5235), .ZN(n_1_737_2184));
   NAND2_X1 i_1_737_2359 (.A1(n_1_737_4416), .A2(n_1_737_3011), .ZN(n_1_737_2185));
   OAI21_X1 i_1_737_2360 (.A(n_1_737_2187), .B1(n_1_737_5434), .B2(n_1_737_5365), 
      .ZN(n_1_737_2186));
   OAI22_X1 i_1_737_2361 (.A1(n_1_737_5625), .A2(n_1_737_3454), .B1(n_1_737_893), 
      .B2(n_1_737_5366), .ZN(n_1_737_2187));
   OAI21_X1 i_1_737_2362 (.A(n_1_737_2189), .B1(n_1_737_5438), .B2(n_1_737_5336), 
      .ZN(n_1_737_2188));
   OAI221_X1 i_1_737_2363 (.A(n_1_737_2190), .B1(n_1_737_4992), .B2(n_1_737_2315), 
      .C1(n_1_737_889), .C2(n_1_737_5337), .ZN(n_1_737_2189));
   NAND2_X1 i_1_737_2364 (.A1(\out_bs[0] [6]), .A2(n_1_737_3427), .ZN(
      n_1_737_2190));
   NOR3_X1 i_1_737_2365 (.A1(n_1_737_4513), .A2(n_1_737_2252), .A3(n_1_737_888), 
      .ZN(n_174));
   OAI21_X1 i_1_737_2366 (.A(n_1_737_888), .B1(n_1_737_4513), .B2(n_1_737_2252), 
      .ZN(n_175));
   NOR2_X1 i_1_737_2367 (.A1(n_1_737_887), .A2(n_1_737_2191), .ZN(n_176));
   NAND2_X1 i_1_737_2368 (.A1(n_1_737_887), .A2(n_1_737_2191), .ZN(n_177));
   NAND3_X1 i_1_737_2369 (.A1(n_845), .A2(n_1_737_4519), .A3(n_844), .ZN(
      n_1_737_2191));
   NAND4_X1 i_1_737_2370 (.A1(n_1_737_2199), .A2(n_1_737_2192), .A3(n_1_737_2196), 
      .A4(n_1_737_2201), .ZN(n_178));
   AOI21_X1 i_1_737_2371 (.A(n_1_737_2193), .B1(n_1_737_2204), .B2(n_1_737_2203), 
      .ZN(n_1_737_2192));
   INV_X1 i_1_737_2372 (.A(n_1_737_2194), .ZN(n_1_737_2193));
   OAI21_X1 i_1_737_2373 (.A(n_1_737_2195), .B1(n_1_737_5442), .B2(n_1_737_5297), 
      .ZN(n_1_737_2194));
   OAI22_X1 i_1_737_2374 (.A1(n_1_737_4528), .A2(n_1_737_3015), .B1(n_1_737_883), 
      .B2(n_1_737_5298), .ZN(n_1_737_2195));
   OAI21_X1 i_1_737_2375 (.A(n_1_737_2197), .B1(n_1_737_5440), .B2(n_1_737_5189), 
      .ZN(n_1_737_2196));
   OAI21_X1 i_1_737_2376 (.A(n_1_737_2198), .B1(n_1_737_885), .B2(n_1_737_5190), 
      .ZN(n_1_737_2197));
   NAND2_X1 i_1_737_2377 (.A1(n_1_737_4535), .A2(n_1_737_3006), .ZN(n_1_737_2198));
   OAI21_X1 i_1_737_2378 (.A(n_1_737_2200), .B1(n_1_737_5441), .B2(n_1_737_5235), 
      .ZN(n_1_737_2199));
   OAI22_X1 i_1_737_2379 (.A1(n_1_737_5257), .A2(n_1_737_2307), .B1(n_1_737_884), 
      .B2(n_1_737_5236), .ZN(n_1_737_2200));
   OAI21_X1 i_1_737_2380 (.A(n_1_737_2202), .B1(n_1_737_5439), .B2(n_1_737_5365), 
      .ZN(n_1_737_2201));
   OAI22_X1 i_1_737_2381 (.A1(n_1_737_5398), .A2(n_1_737_2320), .B1(n_1_737_886), 
      .B2(n_1_737_5366), .ZN(n_1_737_2202));
   OAI21_X1 i_1_737_2382 (.A(n_1_737_882), .B1(n_1_737_5337), .B2(n_1_737_2205), 
      .ZN(n_1_737_2203));
   NAND2_X1 i_1_737_2383 (.A1(n_1_737_5337), .A2(n_1_737_2205), .ZN(n_1_737_2204));
   NAND2_X1 i_1_737_2384 (.A1(n_1_737_4544), .A2(n_1_737_3019), .ZN(n_1_737_2205));
   NOR2_X1 i_1_737_2385 (.A1(n_1_737_881), .A2(n_1_737_2206), .ZN(n_179));
   NAND2_X1 i_1_737_2386 (.A1(n_1_737_881), .A2(n_1_737_2206), .ZN(n_180));
   OAI21_X1 i_1_737_2387 (.A(n_1_737_2253), .B1(n_847), .B2(n_1_737_3942), 
      .ZN(n_1_737_2206));
   NOR3_X1 i_1_737_2388 (.A1(n_1_737_5021), .A2(n_1_737_2298), .A3(n_1_737_880), 
      .ZN(n_181));
   OAI21_X1 i_1_737_2389 (.A(n_1_737_880), .B1(n_1_737_5021), .B2(n_1_737_2298), 
      .ZN(n_182));
   NAND3_X1 i_1_737_2390 (.A1(n_1_737_2212), .A2(n_1_737_2207), .A3(n_1_737_2216), 
      .ZN(n_183));
   AOI211_X1 i_1_737_2391 (.A(n_1_737_2208), .B(n_1_737_2214), .C1(n_1_737_2219), 
      .C2(n_1_737_2218), .ZN(n_1_737_2207));
   INV_X1 i_1_737_2392 (.A(n_1_737_2209), .ZN(n_1_737_2208));
   OAI21_X1 i_1_737_2393 (.A(n_1_737_2210), .B1(n_1_737_5446), .B2(n_1_737_5297), 
      .ZN(n_1_737_2209));
   OAI22_X1 i_1_737_2394 (.A1(n_1_737_5045), .A2(n_1_737_2312), .B1(n_1_737_876), 
      .B2(n_1_737_5298), .ZN(n_1_737_2210));
   INV_X1 i_1_737_2395 (.A(n_1_737_2212), .ZN(n_1_737_2211));
   OAI21_X1 i_1_737_2396 (.A(n_1_737_2213), .B1(n_1_737_5444), .B2(n_1_737_5189), 
      .ZN(n_1_737_2212));
   OAI22_X1 i_1_737_2397 (.A1(n_1_737_5036), .A2(n_1_737_2303), .B1(n_1_737_878), 
      .B2(n_1_737_5190), .ZN(n_1_737_2213));
   AOI21_X1 i_1_737_2398 (.A(n_1_737_2215), .B1(n_1_737_877), .B2(n_1_737_5236), 
      .ZN(n_1_737_2214));
   AOI22_X1 i_1_737_2399 (.A1(n_1_737_4504), .A2(n_1_737_3011), .B1(n_1_737_5445), 
      .B2(n_1_737_5235), .ZN(n_1_737_2215));
   OAI21_X1 i_1_737_2400 (.A(n_1_737_2217), .B1(n_1_737_5443), .B2(n_1_737_5365), 
      .ZN(n_1_737_2216));
   OAI22_X1 i_1_737_2401 (.A1(n_1_737_5063), .A2(n_1_737_2320), .B1(n_1_737_879), 
      .B2(n_1_737_5366), .ZN(n_1_737_2217));
   NAND2_X1 i_1_737_2402 (.A1(n_1_737_875), .A2(n_1_737_5337), .ZN(n_1_737_2218));
   OAI22_X1 i_1_737_2403 (.A1(n_1_737_5028), .A2(n_1_737_2315), .B1(n_1_737_875), 
      .B2(n_1_737_5337), .ZN(n_1_737_2219));
   NOR2_X1 i_1_737_2404 (.A1(n_1_737_874), .A2(n_1_737_2220), .ZN(n_184));
   NAND2_X1 i_1_737_2405 (.A1(n_1_737_874), .A2(n_1_737_2220), .ZN(n_185));
   NAND2_X1 i_1_737_2406 (.A1(n_1_737_4512), .A2(n_1_737_3084), .ZN(n_1_737_2220));
   NOR3_X1 i_1_737_2407 (.A1(n_1_737_4517), .A2(n_1_737_3109), .A3(n_1_737_873), 
      .ZN(n_186));
   OAI21_X1 i_1_737_2408 (.A(n_1_737_873), .B1(n_1_737_4517), .B2(n_1_737_3109), 
      .ZN(n_187));
   OR4_X1 i_1_737_2409 (.A1(n_1_737_2227), .A2(n_1_737_2221), .A3(n_1_737_2224), 
      .A4(n_1_737_2234), .ZN(n_188));
   OAI211_X1 i_1_737_2410 (.A(n_1_737_2222), .B(n_1_737_2231), .C1(n_1_737_868), 
      .C2(n_1_737_2233), .ZN(n_1_737_2221));
   INV_X1 i_1_737_2411 (.A(n_1_737_2223), .ZN(n_1_737_2222));
   AOI21_X1 i_1_737_2412 (.A(n_1_737_5337), .B1(n_1_737_868), .B2(n_1_737_2233), 
      .ZN(n_1_737_2223));
   INV_X1 i_1_737_2413 (.A(n_1_737_2225), .ZN(n_1_737_2224));
   OAI21_X1 i_1_737_2414 (.A(n_1_737_2226), .B1(n_1_737_5448), .B2(n_1_737_5189), 
      .ZN(n_1_737_2225));
   OAI22_X1 i_1_737_2415 (.A1(n_1_737_5638), .A2(n_1_737_3519), .B1(n_1_737_871), 
      .B2(n_1_737_5190), .ZN(n_1_737_2226));
   INV_X1 i_1_737_2416 (.A(n_1_737_2228), .ZN(n_1_737_2227));
   OAI21_X1 i_1_737_2417 (.A(n_1_737_2229), .B1(n_1_737_5449), .B2(n_1_737_5235), 
      .ZN(n_1_737_2228));
   OAI22_X1 i_1_737_2418 (.A1(n_1_737_5651), .A2(n_1_737_3535), .B1(n_1_737_870), 
      .B2(n_1_737_5236), .ZN(n_1_737_2229));
   INV_X1 i_1_737_2419 (.A(n_1_737_2231), .ZN(n_1_737_2230));
   OAI21_X1 i_1_737_2420 (.A(n_1_737_2232), .B1(n_1_737_5450), .B2(n_1_737_5297), 
      .ZN(n_1_737_2231));
   OAI22_X1 i_1_737_2421 (.A1(n_1_737_5664), .A2(n_1_737_3528), .B1(n_1_737_869), 
      .B2(n_1_737_5298), .ZN(n_1_737_2232));
   NAND2_X1 i_1_737_2422 (.A1(\out_bs[0] [6]), .A2(n_1_737_3513), .ZN(
      n_1_737_2233));
   INV_X1 i_1_737_2423 (.A(n_1_737_2235), .ZN(n_1_737_2234));
   OAI21_X1 i_1_737_2424 (.A(n_1_737_2236), .B1(n_1_737_5447), .B2(n_1_737_5365), 
      .ZN(n_1_737_2235));
   OAI22_X1 i_1_737_2425 (.A1(n_1_737_5625), .A2(n_1_737_3542), .B1(n_1_737_872), 
      .B2(n_1_737_5366), .ZN(n_1_737_2236));
   NOR2_X1 i_1_737_2426 (.A1(n_1_737_867), .A2(n_1_737_2237), .ZN(n_189));
   NAND2_X1 i_1_737_2427 (.A1(n_1_737_867), .A2(n_1_737_2237), .ZN(n_190));
   OAI21_X1 i_1_737_2428 (.A(n_1_737_2253), .B1(n_847), .B2(n_1_737_4015), 
      .ZN(n_1_737_2237));
   NOR3_X1 i_1_737_2429 (.A1(n_1_737_5171), .A2(n_1_737_2298), .A3(n_1_737_866), 
      .ZN(n_191));
   OAI21_X1 i_1_737_2430 (.A(n_1_737_866), .B1(n_1_737_5171), .B2(n_1_737_2298), 
      .ZN(n_192));
   OR3_X1 i_1_737_2431 (.A1(n_1_737_2250), .A2(n_1_737_2249), .A3(n_1_737_2238), 
      .ZN(n_193));
   NAND4_X1 i_1_737_2432 (.A1(n_1_737_2241), .A2(n_1_737_2239), .A3(n_1_737_2244), 
      .A4(n_1_737_2247), .ZN(n_1_737_2238));
   OAI21_X1 i_1_737_2433 (.A(n_1_737_2240), .B1(n_1_737_5454), .B2(n_1_737_5297), 
      .ZN(n_1_737_2239));
   OAI22_X1 i_1_737_2434 (.A1(n_1_737_5286), .A2(n_1_737_2312), .B1(n_1_737_862), 
      .B2(n_1_737_5298), .ZN(n_1_737_2240));
   OAI21_X1 i_1_737_2435 (.A(n_1_737_2242), .B1(n_1_737_5452), .B2(n_1_737_5189), 
      .ZN(n_1_737_2241));
   OAI21_X1 i_1_737_2436 (.A(n_1_737_2243), .B1(n_1_737_864), .B2(n_1_737_5190), 
      .ZN(n_1_737_2242));
   NAND2_X1 i_1_737_2437 (.A1(n_1_737_4576), .A2(n_1_737_3006), .ZN(n_1_737_2243));
   OAI21_X1 i_1_737_2438 (.A(n_1_737_2245), .B1(n_1_737_5453), .B2(n_1_737_5235), 
      .ZN(n_1_737_2244));
   OAI21_X1 i_1_737_2439 (.A(n_1_737_2246), .B1(n_1_737_863), .B2(n_1_737_5236), 
      .ZN(n_1_737_2245));
   NAND2_X1 i_1_737_2440 (.A1(n_1_737_4588), .A2(n_1_737_3011), .ZN(n_1_737_2246));
   OAI21_X1 i_1_737_2441 (.A(n_1_737_2248), .B1(n_1_737_5451), .B2(n_1_737_5365), 
      .ZN(n_1_737_2247));
   OAI22_X1 i_1_737_2442 (.A1(n_1_737_5395), .A2(n_1_737_2320), .B1(n_1_737_865), 
      .B2(n_1_737_5366), .ZN(n_1_737_2248));
   AOI21_X1 i_1_737_2443 (.A(n_1_737_5337), .B1(n_1_737_861), .B2(n_1_737_2251), 
      .ZN(n_1_737_2249));
   NOR2_X1 i_1_737_2444 (.A1(n_1_737_861), .A2(n_1_737_2251), .ZN(n_1_737_2250));
   NAND2_X1 i_1_737_2445 (.A1(n_1_737_4571), .A2(n_1_737_3019), .ZN(n_1_737_2251));
   NOR2_X1 i_1_737_2446 (.A1(n_1_737_860), .A2(n_1_737_2252), .ZN(n_194));
   NAND2_X1 i_1_737_2447 (.A1(n_1_737_860), .A2(n_1_737_2252), .ZN(n_195));
   INV_X1 i_1_737_2448 (.A(n_1_737_2253), .ZN(n_1_737_2252));
   NOR2_X1 i_1_737_2449 (.A1(n_1_737_5607), .A2(n_1_737_3546), .ZN(n_1_737_2253));
   NOR2_X1 i_1_737_2450 (.A1(n_1_737_859), .A2(n_1_737_2298), .ZN(n_196));
   NAND2_X1 i_1_737_2451 (.A1(n_1_737_859), .A2(n_1_737_2298), .ZN(n_197));
   OAI211_X1 i_1_737_2452 (.A(n_1_737_2265), .B(n_1_737_2254), .C1(n_1_737_854), 
      .C2(n_1_737_2315), .ZN(n_198));
   NOR4_X1 i_1_737_2453 (.A1(n_1_737_2258), .A2(n_1_737_2255), .A3(n_1_737_2260), 
      .A4(n_1_737_2263), .ZN(n_1_737_2254));
   INV_X1 i_1_737_2454 (.A(n_1_737_2256), .ZN(n_1_737_2255));
   OAI21_X1 i_1_737_2455 (.A(n_1_737_2257), .B1(n_1_737_5297), .B2(n_1_737_2313), 
      .ZN(n_1_737_2256));
   OAI21_X1 i_1_737_2456 (.A(n_1_737_855), .B1(n_1_737_5298), .B2(n_1_737_2312), 
      .ZN(n_1_737_2257));
   OAI22_X1 i_1_737_2457 (.A1(n_1_737_857), .A2(n_1_737_2303), .B1(n_1_737_5190), 
      .B2(n_1_737_2259), .ZN(n_1_737_2258));
   AND2_X1 i_1_737_2458 (.A1(n_1_737_857), .A2(n_1_737_2303), .ZN(n_1_737_2259));
   OAI22_X1 i_1_737_2459 (.A1(n_1_737_856), .A2(n_1_737_2307), .B1(n_1_737_5236), 
      .B2(n_1_737_2261), .ZN(n_1_737_2260));
   AND2_X1 i_1_737_2460 (.A1(n_1_737_856), .A2(n_1_737_2307), .ZN(n_1_737_2261));
   INV_X1 i_1_737_2461 (.A(n_1_737_2263), .ZN(n_1_737_2262));
   OAI22_X1 i_1_737_2462 (.A1(n_1_737_858), .A2(n_1_737_2320), .B1(n_1_737_5366), 
      .B2(n_1_737_2264), .ZN(n_1_737_2263));
   AND2_X1 i_1_737_2463 (.A1(n_1_737_858), .A2(n_1_737_2320), .ZN(n_1_737_2264));
   INV_X1 i_1_737_2464 (.A(n_1_737_2266), .ZN(n_1_737_2265));
   AOI21_X1 i_1_737_2465 (.A(n_1_737_5337), .B1(n_1_737_854), .B2(n_1_737_2315), 
      .ZN(n_1_737_2266));
   NOR2_X1 i_1_737_2466 (.A1(n_1_737_852), .A2(n_1_737_2267), .ZN(n_199));
   NAND2_X1 i_1_737_2467 (.A1(n_1_737_852), .A2(n_1_737_2267), .ZN(n_200));
   AOI21_X1 i_1_737_2468 (.A(n_1_737_2299), .B1(n_1_737_4615), .B2(n_1_737_3110), 
      .ZN(n_1_737_2267));
   NAND4_X1 i_1_737_2469 (.A1(n_1_737_2276), .A2(n_1_737_2268), .A3(n_1_737_2273), 
      .A4(n_1_737_2281), .ZN(n_201));
   AOI21_X1 i_1_737_2470 (.A(n_1_737_2270), .B1(n_1_737_2279), .B2(n_1_737_2278), 
      .ZN(n_1_737_2268));
   INV_X1 i_1_737_2471 (.A(n_1_737_2270), .ZN(n_1_737_2269));
   OAI22_X1 i_1_737_2472 (.A1(n_1_737_848), .A2(n_1_737_5298), .B1(n_1_737_2272), 
      .B2(n_1_737_2271), .ZN(n_1_737_2270));
   AOI21_X1 i_1_737_2473 (.A(n_1_737_2313), .B1(n_1_737_4632), .B2(n_1_737_3016), 
      .ZN(n_1_737_2271));
   AND2_X1 i_1_737_2474 (.A1(n_1_737_848), .A2(n_1_737_5298), .ZN(n_1_737_2272));
   OAI22_X1 i_1_737_2475 (.A1(n_1_737_5456), .A2(n_1_737_5189), .B1(n_1_737_2275), 
      .B2(n_1_737_2274), .ZN(n_1_737_2273));
   NOR2_X1 i_1_737_2476 (.A1(n_1_737_850), .A2(n_1_737_5190), .ZN(n_1_737_2274));
   OAI21_X1 i_1_737_2477 (.A(n_1_737_2303), .B1(n_1_737_4622), .B2(n_1_737_3005), 
      .ZN(n_1_737_2275));
   OAI21_X1 i_1_737_2478 (.A(n_1_737_2277), .B1(n_1_737_5457), .B2(n_1_737_5235), 
      .ZN(n_1_737_2276));
   OAI221_X1 i_1_737_2479 (.A(n_1_737_2307), .B1(n_1_737_4638), .B2(n_1_737_3010), 
      .C1(n_1_737_849), .C2(n_1_737_5236), .ZN(n_1_737_2277));
   OAI221_X1 i_1_737_2480 (.A(n_1_737_2315), .B1(n_1_737_4626), .B2(n_1_737_3018), 
      .C1(n_1_737_847), .C2(n_1_737_5337), .ZN(n_1_737_2278));
   NAND2_X1 i_1_737_2481 (.A1(n_1_737_847), .A2(n_1_737_5337), .ZN(n_1_737_2279));
   INV_X1 i_1_737_2482 (.A(n_1_737_2281), .ZN(n_1_737_2280));
   OAI21_X1 i_1_737_2483 (.A(n_1_737_2282), .B1(n_1_737_5455), .B2(n_1_737_5365), 
      .ZN(n_1_737_2281));
   OAI221_X1 i_1_737_2484 (.A(n_1_737_2320), .B1(n_1_737_4643), .B2(n_1_737_3022), 
      .C1(n_1_737_851), .C2(n_1_737_5366), .ZN(n_1_737_2282));
   NOR2_X1 i_1_737_2485 (.A1(n_1_737_845), .A2(n_1_737_2283), .ZN(n_202));
   NAND2_X1 i_1_737_2486 (.A1(n_1_737_845), .A2(n_1_737_2283), .ZN(n_203));
   OAI21_X1 i_1_737_2487 (.A(n_1_737_3110), .B1(n_848), .B2(n_1_737_4646), 
      .ZN(n_1_737_2283));
   NAND4_X1 i_1_737_2488 (.A1(n_1_737_2287), .A2(n_1_737_2284), .A3(n_1_737_2293), 
      .A4(n_1_737_2295), .ZN(n_204));
   AOI21_X1 i_1_737_2489 (.A(n_1_737_2290), .B1(n_1_737_2286), .B2(n_1_737_2285), 
      .ZN(n_1_737_2284));
   OAI221_X1 i_1_737_2490 (.A(n_1_737_2315), .B1(n_1_737_4669), .B2(n_1_737_3018), 
      .C1(n_1_737_840), .C2(n_1_737_5337), .ZN(n_1_737_2285));
   NAND2_X1 i_1_737_2491 (.A1(n_1_737_840), .A2(n_1_737_5337), .ZN(n_1_737_2286));
   OAI21_X1 i_1_737_2492 (.A(n_1_737_2288), .B1(n_1_737_5460), .B2(n_1_737_5235), 
      .ZN(n_1_737_2287));
   OAI221_X1 i_1_737_2493 (.A(n_1_737_2307), .B1(n_1_737_4664), .B2(n_1_737_3010), 
      .C1(n_1_737_842), .C2(n_1_737_5236), .ZN(n_1_737_2288));
   INV_X1 i_1_737_2494 (.A(n_1_737_2290), .ZN(n_1_737_2289));
   OAI22_X1 i_1_737_2495 (.A1(n_1_737_841), .A2(n_1_737_5298), .B1(n_1_737_2292), 
      .B2(n_1_737_2291), .ZN(n_1_737_2290));
   AOI21_X1 i_1_737_2496 (.A(n_1_737_2313), .B1(n_1_737_4652), .B2(n_1_737_3016), 
      .ZN(n_1_737_2291));
   AND2_X1 i_1_737_2497 (.A1(n_1_737_841), .A2(n_1_737_5298), .ZN(n_1_737_2292));
   OAI21_X1 i_1_737_2498 (.A(n_1_737_2294), .B1(n_1_737_5459), .B2(n_1_737_5189), 
      .ZN(n_1_737_2293));
   OAI221_X1 i_1_737_2499 (.A(n_1_737_2303), .B1(n_1_737_4658), .B2(n_1_737_3005), 
      .C1(n_1_737_843), .C2(n_1_737_5190), .ZN(n_1_737_2294));
   OAI21_X1 i_1_737_2500 (.A(n_1_737_2296), .B1(n_1_737_5458), .B2(n_1_737_5365), 
      .ZN(n_1_737_2295));
   OAI221_X1 i_1_737_2501 (.A(n_1_737_2320), .B1(n_1_737_4676), .B2(n_1_737_3022), 
      .C1(n_1_737_844), .C2(n_1_737_5366), .ZN(n_1_737_2296));
   NOR2_X1 i_1_737_2502 (.A1(n_1_737_838), .A2(n_1_737_2297), .ZN(n_205));
   NAND2_X1 i_1_737_2503 (.A1(n_1_737_838), .A2(n_1_737_2297), .ZN(n_206));
   OAI21_X1 i_1_737_2504 (.A(n_1_737_3110), .B1(n_848), .B2(n_1_737_4679), 
      .ZN(n_1_737_2297));
   INV_X1 i_1_737_2505 (.A(n_1_737_2299), .ZN(n_1_737_2298));
   NOR2_X1 i_1_737_2506 (.A1(n_1_737_5612), .A2(n_1_737_3756), .ZN(n_1_737_2299));
   OR4_X1 i_1_737_2507 (.A1(n_1_737_2308), .A2(n_1_737_2304), .A3(n_1_737_2300), 
      .A4(n_1_737_2317), .ZN(n_207));
   AOI21_X1 i_1_737_2508 (.A(n_1_737_2301), .B1(n_1_737_836), .B2(n_1_737_5190), 
      .ZN(n_1_737_2300));
   INV_X1 i_1_737_2509 (.A(n_1_737_2302), .ZN(n_1_737_2301));
   OAI221_X1 i_1_737_2510 (.A(n_1_737_2303), .B1(n_1_737_4691), .B2(n_1_737_3005), 
      .C1(n_1_737_836), .C2(n_1_737_5190), .ZN(n_1_737_2302));
   NAND2_X1 i_1_737_2511 (.A1(\out_bs[3] [6]), .A2(n_1_737_3799), .ZN(
      n_1_737_2303));
   AOI21_X1 i_1_737_2512 (.A(n_1_737_2305), .B1(n_1_737_835), .B2(n_1_737_5236), 
      .ZN(n_1_737_2304));
   INV_X1 i_1_737_2513 (.A(n_1_737_2306), .ZN(n_1_737_2305));
   OAI22_X1 i_1_737_2514 (.A1(n_1_737_835), .A2(n_1_737_5236), .B1(n_1_737_4705), 
      .B2(n_1_737_3010), .ZN(n_1_737_2306));
   NAND2_X1 i_1_737_2515 (.A1(\out_bs[2] [6]), .A2(n_1_737_3778), .ZN(
      n_1_737_2307));
   OAI221_X1 i_1_737_2516 (.A(n_1_737_2310), .B1(n_1_737_833), .B2(n_1_737_5337), 
      .C1(n_1_737_2316), .C2(n_1_737_2314), .ZN(n_1_737_2308));
   INV_X1 i_1_737_2517 (.A(n_1_737_2310), .ZN(n_1_737_2309));
   OAI21_X1 i_1_737_2518 (.A(n_1_737_2311), .B1(n_1_737_5461), .B2(n_1_737_5297), 
      .ZN(n_1_737_2310));
   OAI22_X1 i_1_737_2519 (.A1(n_1_737_834), .A2(n_1_737_5298), .B1(n_1_737_4697), 
      .B2(n_1_737_3015), .ZN(n_1_737_2311));
   INV_X1 i_1_737_2520 (.A(n_1_737_2313), .ZN(n_1_737_2312));
   NOR2_X1 i_1_737_2521 (.A1(n_1_737_5664), .A2(n_1_737_3788), .ZN(n_1_737_2313));
   OAI21_X1 i_1_737_2522 (.A(n_1_737_3019), .B1(\out_bs[0] [4]), .B2(
      n_1_737_4686), .ZN(n_1_737_2314));
   NAND2_X1 i_1_737_2523 (.A1(\out_bs[0] [6]), .A2(n_1_737_3769), .ZN(
      n_1_737_2315));
   AND2_X1 i_1_737_2524 (.A1(n_1_737_833), .A2(n_1_737_5337), .ZN(n_1_737_2316));
   AOI21_X1 i_1_737_2525 (.A(n_1_737_2318), .B1(n_1_737_837), .B2(n_1_737_5366), 
      .ZN(n_1_737_2317));
   INV_X1 i_1_737_2526 (.A(n_1_737_2319), .ZN(n_1_737_2318));
   OAI22_X1 i_1_737_2527 (.A1(n_1_737_4713), .A2(n_1_737_3022), .B1(n_1_737_837), 
      .B2(n_1_737_5366), .ZN(n_1_737_2319));
   NAND2_X1 i_1_737_2528 (.A1(\out_bs[4] [6]), .A2(n_1_737_3810), .ZN(
      n_1_737_2320));
   NOR3_X1 i_1_737_2529 (.A1(n_1_737_3696), .A2(n_1_737_3083), .A3(n_1_737_832), 
      .ZN(n_208));
   OAI21_X1 i_1_737_2530 (.A(n_1_737_832), .B1(n_1_737_3696), .B2(n_1_737_3083), 
      .ZN(n_209));
   NOR3_X1 i_1_737_2531 (.A1(n_1_737_4740), .A2(n_1_737_3109), .A3(n_1_737_831), 
      .ZN(n_210));
   OAI21_X1 i_1_737_2532 (.A(n_1_737_831), .B1(n_1_737_4740), .B2(n_1_737_3109), 
      .ZN(n_211));
   OAI211_X1 i_1_737_2533 (.A(n_1_737_2334), .B(n_1_737_2321), .C1(n_1_737_826), 
      .C2(n_1_737_2336), .ZN(n_212));
   NOR4_X1 i_1_737_2534 (.A1(n_1_737_2325), .A2(n_1_737_2322), .A3(n_1_737_2328), 
      .A4(n_1_737_2331), .ZN(n_1_737_2321));
   INV_X1 i_1_737_2535 (.A(n_1_737_2323), .ZN(n_1_737_2322));
   OAI21_X1 i_1_737_2536 (.A(n_1_737_2324), .B1(n_1_737_5463), .B2(n_1_737_5297), 
      .ZN(n_1_737_2323));
   OAI22_X1 i_1_737_2537 (.A1(n_1_737_4752), .A2(n_1_737_3015), .B1(n_1_737_827), 
      .B2(n_1_737_5298), .ZN(n_1_737_2324));
   INV_X1 i_1_737_2538 (.A(n_1_737_2326), .ZN(n_1_737_2325));
   OAI21_X1 i_1_737_2539 (.A(n_1_737_2327), .B1(n_1_737_5462), .B2(n_1_737_5189), 
      .ZN(n_1_737_2326));
   OAI22_X1 i_1_737_2540 (.A1(n_1_737_4762), .A2(n_1_737_3005), .B1(n_1_737_829), 
      .B2(n_1_737_5190), .ZN(n_1_737_2327));
   AOI21_X1 i_1_737_2541 (.A(n_1_737_2329), .B1(n_1_737_828), .B2(n_1_737_5236), 
      .ZN(n_1_737_2328));
   INV_X1 i_1_737_2542 (.A(n_1_737_2330), .ZN(n_1_737_2329));
   OAI22_X1 i_1_737_2543 (.A1(n_1_737_4771), .A2(n_1_737_3010), .B1(n_1_737_828), 
      .B2(n_1_737_5236), .ZN(n_1_737_2330));
   AOI21_X1 i_1_737_2544 (.A(n_1_737_2332), .B1(n_1_737_830), .B2(n_1_737_5366), 
      .ZN(n_1_737_2331));
   INV_X1 i_1_737_2545 (.A(n_1_737_2333), .ZN(n_1_737_2332));
   OAI22_X1 i_1_737_2546 (.A1(n_1_737_4789), .A2(n_1_737_3022), .B1(n_1_737_830), 
      .B2(n_1_737_5366), .ZN(n_1_737_2333));
   INV_X1 i_1_737_2547 (.A(n_1_737_2335), .ZN(n_1_737_2334));
   AOI21_X1 i_1_737_2548 (.A(n_1_737_5337), .B1(n_1_737_826), .B2(n_1_737_2336), 
      .ZN(n_1_737_2335));
   OAI21_X1 i_1_737_2549 (.A(n_1_737_3019), .B1(\out_bs[0] [4]), .B2(
      n_1_737_4780), .ZN(n_1_737_2336));
   NOR3_X1 i_1_737_2550 (.A1(n_1_737_4737), .A2(n_1_737_3109), .A3(n_1_737_824), 
      .ZN(n_213));
   OAI21_X1 i_1_737_2551 (.A(n_1_737_824), .B1(n_1_737_4737), .B2(n_1_737_3109), 
      .ZN(n_214));
   NAND4_X1 i_1_737_2552 (.A1(n_1_737_2339), .A2(n_1_737_2337), .A3(n_1_737_2341), 
      .A4(n_1_737_2350), .ZN(n_215));
   OAI21_X1 i_1_737_2553 (.A(n_1_737_5467), .B1(n_1_737_5336), .B2(n_1_737_2342), 
      .ZN(n_1_737_2337));
   INV_X1 i_1_737_2554 (.A(n_1_737_2339), .ZN(n_1_737_2338));
   OAI21_X1 i_1_737_2555 (.A(n_1_737_2340), .B1(n_1_737_5465), .B2(n_1_737_5235), 
      .ZN(n_1_737_2339));
   OAI22_X1 i_1_737_2556 (.A1(n_1_737_4769), .A2(n_1_737_3010), .B1(n_1_737_821), 
      .B2(n_1_737_5236), .ZN(n_1_737_2340));
   AOI211_X1 i_1_737_2557 (.A(n_1_737_2343), .B(n_1_737_2346), .C1(n_1_737_5336), 
      .C2(n_1_737_2342), .ZN(n_1_737_2341));
   NOR2_X1 i_1_737_2558 (.A1(n_1_737_4777), .A2(n_1_737_3018), .ZN(n_1_737_2342));
   INV_X1 i_1_737_2559 (.A(n_1_737_2344), .ZN(n_1_737_2343));
   OAI21_X1 i_1_737_2560 (.A(n_1_737_2345), .B1(n_1_737_5466), .B2(n_1_737_5297), 
      .ZN(n_1_737_2344));
   OAI22_X1 i_1_737_2561 (.A1(n_1_737_4750), .A2(n_1_737_3015), .B1(n_1_737_820), 
      .B2(n_1_737_5298), .ZN(n_1_737_2345));
   AOI21_X1 i_1_737_2562 (.A(n_1_737_2347), .B1(n_1_737_822), .B2(n_1_737_5190), 
      .ZN(n_1_737_2346));
   INV_X1 i_1_737_2563 (.A(n_1_737_2348), .ZN(n_1_737_2347));
   OAI22_X1 i_1_737_2564 (.A1(n_1_737_4760), .A2(n_1_737_3005), .B1(n_1_737_822), 
      .B2(n_1_737_5190), .ZN(n_1_737_2348));
   INV_X1 i_1_737_2565 (.A(n_1_737_2350), .ZN(n_1_737_2349));
   OAI21_X1 i_1_737_2566 (.A(n_1_737_2351), .B1(n_1_737_5464), .B2(n_1_737_5365), 
      .ZN(n_1_737_2350));
   OAI22_X1 i_1_737_2567 (.A1(n_1_737_4787), .A2(n_1_737_3022), .B1(n_1_737_823), 
      .B2(n_1_737_5366), .ZN(n_1_737_2351));
   NOR2_X1 i_1_737_2568 (.A1(n_1_737_818), .A2(n_1_737_2352), .ZN(n_216));
   NAND2_X1 i_1_737_2569 (.A1(n_1_737_818), .A2(n_1_737_2352), .ZN(n_217));
   NAND2_X1 i_1_737_2570 (.A1(n_1_737_3750), .A2(n_1_737_3084), .ZN(n_1_737_2352));
   NOR2_X1 i_1_737_2571 (.A1(n_1_737_817), .A2(n_1_737_2353), .ZN(n_218));
   NAND2_X1 i_1_737_2572 (.A1(n_1_737_817), .A2(n_1_737_2353), .ZN(n_219));
   NAND2_X1 i_1_737_2573 (.A1(n_1_737_4812), .A2(n_1_737_3110), .ZN(n_1_737_2353));
   NAND4_X1 i_1_737_2574 (.A1(n_1_737_2358), .A2(n_1_737_2356), .A3(n_1_737_2354), 
      .A4(n_1_737_2365), .ZN(n_220));
   OAI21_X1 i_1_737_2575 (.A(n_1_737_2355), .B1(n_1_737_5469), .B2(n_1_737_5189), 
      .ZN(n_1_737_2354));
   OAI22_X1 i_1_737_2576 (.A1(n_1_737_5638), .A2(n_1_737_3798), .B1(n_1_737_815), 
      .B2(n_1_737_5190), .ZN(n_1_737_2355));
   OAI21_X1 i_1_737_2577 (.A(n_1_737_2357), .B1(n_1_737_5470), .B2(n_1_737_5235), 
      .ZN(n_1_737_2356));
   OAI22_X1 i_1_737_2578 (.A1(n_1_737_5651), .A2(n_1_737_3777), .B1(n_1_737_814), 
      .B2(n_1_737_5236), .ZN(n_1_737_2357));
   AOI211_X1 i_1_737_2579 (.A(n_1_737_2359), .B(n_1_737_2362), .C1(n_1_737_5336), 
      .C2(n_1_737_2364), .ZN(n_1_737_2358));
   AOI21_X1 i_1_737_2580 (.A(n_1_737_2360), .B1(n_1_737_813), .B2(n_1_737_5298), 
      .ZN(n_1_737_2359));
   INV_X1 i_1_737_2581 (.A(n_1_737_2361), .ZN(n_1_737_2360));
   OAI22_X1 i_1_737_2582 (.A1(n_1_737_5664), .A2(n_1_737_3787), .B1(n_1_737_813), 
      .B2(n_1_737_5298), .ZN(n_1_737_2361));
   AOI21_X1 i_1_737_2583 (.A(n_1_737_812), .B1(n_1_737_5337), .B2(n_1_737_2363), 
      .ZN(n_1_737_2362));
   INV_X1 i_1_737_2584 (.A(n_1_737_2364), .ZN(n_1_737_2363));
   NOR2_X1 i_1_737_2585 (.A1(n_1_737_5671), .A2(n_1_737_3767), .ZN(n_1_737_2364));
   OAI21_X1 i_1_737_2586 (.A(n_1_737_2366), .B1(n_1_737_5468), .B2(n_1_737_5365), 
      .ZN(n_1_737_2365));
   OAI22_X1 i_1_737_2587 (.A1(n_1_737_5625), .A2(n_1_737_3809), .B1(n_1_737_816), 
      .B2(n_1_737_5366), .ZN(n_1_737_2366));
   NOR2_X1 i_1_737_2588 (.A1(n_1_737_811), .A2(n_1_737_2367), .ZN(n_221));
   NAND2_X1 i_1_737_2589 (.A1(n_1_737_811), .A2(n_1_737_2367), .ZN(n_222));
   OR2_X1 i_1_737_2590 (.A1(n_1_737_3749), .A2(n_1_737_3083), .ZN(n_1_737_2367));
   NOR2_X1 i_1_737_2591 (.A1(n_1_737_810), .A2(n_1_737_2368), .ZN(n_223));
   NAND2_X1 i_1_737_2592 (.A1(n_1_737_810), .A2(n_1_737_2368), .ZN(n_224));
   OR2_X1 i_1_737_2593 (.A1(n_1_737_5612), .A2(n_1_737_3755), .ZN(n_1_737_2368));
   NAND4_X1 i_1_737_2594 (.A1(n_1_737_2373), .A2(n_1_737_2371), .A3(n_1_737_2369), 
      .A4(n_1_737_2380), .ZN(n_225));
   OAI21_X1 i_1_737_2595 (.A(n_1_737_2370), .B1(n_1_737_5472), .B2(n_1_737_5189), 
      .ZN(n_1_737_2369));
   OAI22_X1 i_1_737_2596 (.A1(n_1_737_4829), .A2(n_1_737_3005), .B1(n_1_737_808), 
      .B2(n_1_737_5190), .ZN(n_1_737_2370));
   OAI21_X1 i_1_737_2597 (.A(n_1_737_2372), .B1(n_1_737_5473), .B2(n_1_737_5235), 
      .ZN(n_1_737_2371));
   OAI22_X1 i_1_737_2598 (.A1(n_1_737_4850), .A2(n_1_737_3010), .B1(n_1_737_807), 
      .B2(n_1_737_5236), .ZN(n_1_737_2372));
   AOI211_X1 i_1_737_2599 (.A(n_1_737_2374), .B(n_1_737_2377), .C1(n_1_737_5336), 
      .C2(n_1_737_2378), .ZN(n_1_737_2373));
   AOI21_X1 i_1_737_2600 (.A(n_1_737_2375), .B1(n_1_737_806), .B2(n_1_737_5298), 
      .ZN(n_1_737_2374));
   INV_X1 i_1_737_2601 (.A(n_1_737_2376), .ZN(n_1_737_2375));
   OAI22_X1 i_1_737_2602 (.A1(n_1_737_5664), .A2(n_1_737_3785), .B1(n_1_737_806), 
      .B2(n_1_737_5298), .ZN(n_1_737_2376));
   AOI21_X1 i_1_737_2603 (.A(n_1_737_805), .B1(n_1_737_5337), .B2(n_1_737_2379), 
      .ZN(n_1_737_2377));
   INV_X1 i_1_737_2604 (.A(n_1_737_2379), .ZN(n_1_737_2378));
   OAI211_X1 i_1_737_2605 (.A(\out_bs[0] [5]), .B(\out_bs[0] [6]), .C1(
      \out_bs[0] [4]), .C2(n_1_737_4819), .ZN(n_1_737_2379));
   OAI21_X1 i_1_737_2606 (.A(n_1_737_2381), .B1(n_1_737_5471), .B2(n_1_737_5365), 
      .ZN(n_1_737_2380));
   OAI22_X1 i_1_737_2607 (.A1(n_1_737_5625), .A2(n_1_737_3808), .B1(n_1_737_809), 
      .B2(n_1_737_5366), .ZN(n_1_737_2381));
   NAND4_X1 i_1_737_2608 (.A1(n_1_737_2393), .A2(n_1_737_2382), .A3(n_1_737_2385), 
      .A4(n_1_737_2391), .ZN(n_226));
   AOI211_X1 i_1_737_2609 (.A(n_1_737_2389), .B(n_1_737_2396), .C1(n_1_737_2384), 
      .C2(n_1_737_2383), .ZN(n_1_737_2382));
   NAND2_X1 i_1_737_2610 (.A1(n_1_737_798), .A2(n_1_737_5337), .ZN(n_1_737_2383));
   OAI22_X1 i_1_737_2611 (.A1(n_1_737_5334), .A2(n_1_737_3018), .B1(n_1_737_798), 
      .B2(n_1_737_5337), .ZN(n_1_737_2384));
   INV_X1 i_1_737_2612 (.A(n_1_737_2386), .ZN(n_1_737_2385));
   OAI22_X1 i_1_737_2613 (.A1(n_1_737_802), .A2(n_1_737_2417), .B1(n_1_737_5366), 
      .B2(n_1_737_2387), .ZN(n_1_737_2386));
   AND2_X1 i_1_737_2614 (.A1(n_1_737_802), .A2(n_1_737_2417), .ZN(n_1_737_2387));
   INV_X1 i_1_737_2615 (.A(n_1_737_2389), .ZN(n_1_737_2388));
   OAI22_X1 i_1_737_2616 (.A1(n_1_737_799), .A2(n_1_737_2404), .B1(n_1_737_5298), 
      .B2(n_1_737_2390), .ZN(n_1_737_2389));
   AND2_X1 i_1_737_2617 (.A1(n_1_737_799), .A2(n_1_737_2404), .ZN(n_1_737_2390));
   OAI21_X1 i_1_737_2618 (.A(n_1_737_2392), .B1(n_1_737_5602), .B2(n_1_737_5474), 
      .ZN(n_1_737_2391));
   OAI22_X1 i_1_737_2619 (.A1(n_1_737_5178), .A2(n_1_737_3109), .B1(n_1089), 
      .B2(n_1_737_803), .ZN(n_1_737_2392));
   INV_X1 i_1_737_2620 (.A(n_1_737_2394), .ZN(n_1_737_2393));
   OAI22_X1 i_1_737_2621 (.A1(n_1_737_801), .A2(n_1_737_2409), .B1(n_1_737_5190), 
      .B2(n_1_737_2395), .ZN(n_1_737_2394));
   AND2_X1 i_1_737_2622 (.A1(n_1_737_801), .A2(n_1_737_2409), .ZN(n_1_737_2395));
   OAI22_X1 i_1_737_2623 (.A1(n_1_737_800), .A2(n_1_737_2413), .B1(n_1_737_5236), 
      .B2(n_1_737_2397), .ZN(n_1_737_2396));
   AND2_X1 i_1_737_2624 (.A1(n_1_737_800), .A2(n_1_737_2413), .ZN(n_1_737_2397));
   NOR2_X1 i_1_737_2625 (.A1(n_1_737_797), .A2(n_1_737_2398), .ZN(n_227));
   NAND2_X1 i_1_737_2626 (.A1(n_1_737_797), .A2(n_1_737_2398), .ZN(n_228));
   NAND2_X1 i_1_737_2627 (.A1(n_1_737_3831), .A2(n_1_737_3084), .ZN(n_1_737_2398));
   NOR2_X1 i_1_737_2628 (.A1(n_1_737_796), .A2(n_1_737_2399), .ZN(n_229));
   NAND2_X1 i_1_737_2629 (.A1(n_1_737_796), .A2(n_1_737_2399), .ZN(n_230));
   NAND2_X1 i_1_737_2630 (.A1(n_1_737_4881), .A2(n_1_737_3110), .ZN(n_1_737_2399));
   NAND3_X1 i_1_737_2631 (.A1(n_1_737_2415), .A2(n_1_737_2400), .A3(n_1_737_2418), 
      .ZN(n_231));
   NOR3_X1 i_1_737_2632 (.A1(n_1_737_2406), .A2(n_1_737_2402), .A3(n_1_737_2410), 
      .ZN(n_1_737_2400));
   INV_X1 i_1_737_2633 (.A(n_1_737_2402), .ZN(n_1_737_2401));
   OAI22_X1 i_1_737_2634 (.A1(n_1_737_792), .A2(n_1_737_5298), .B1(n_1_737_2405), 
      .B2(n_1_737_2403), .ZN(n_1_737_2402));
   AOI22_X1 i_1_737_2635 (.A1(\out_bs[1] [6]), .A2(n_1_737_4050), .B1(
      n_1_737_4890), .B2(n_1_737_3016), .ZN(n_1_737_2403));
   NAND2_X1 i_1_737_2636 (.A1(\out_bs[1] [6]), .A2(n_1_737_4050), .ZN(
      n_1_737_2404));
   AND2_X1 i_1_737_2637 (.A1(n_1_737_792), .A2(n_1_737_5298), .ZN(n_1_737_2405));
   AOI21_X1 i_1_737_2638 (.A(n_1_737_2407), .B1(n_1_737_794), .B2(n_1_737_5190), 
      .ZN(n_1_737_2406));
   INV_X1 i_1_737_2639 (.A(n_1_737_2408), .ZN(n_1_737_2407));
   OAI221_X1 i_1_737_2640 (.A(n_1_737_2409), .B1(n_1_737_4895), .B2(n_1_737_3005), 
      .C1(n_1_737_794), .C2(n_1_737_5190), .ZN(n_1_737_2408));
   NAND2_X1 i_1_737_2641 (.A1(\out_bs[3] [6]), .A2(n_1_737_4039), .ZN(
      n_1_737_2409));
   OAI22_X1 i_1_737_2642 (.A1(n_1_737_793), .A2(n_1_737_5236), .B1(n_1_737_2412), 
      .B2(n_1_737_2411), .ZN(n_1_737_2410));
   AND2_X1 i_1_737_2643 (.A1(n_1_737_793), .A2(n_1_737_5236), .ZN(n_1_737_2411));
   AOI22_X1 i_1_737_2644 (.A1(\out_bs[2] [6]), .A2(n_1_737_4062), .B1(
      n_1_737_4901), .B2(n_1_737_3011), .ZN(n_1_737_2412));
   NAND2_X1 i_1_737_2645 (.A1(\out_bs[2] [6]), .A2(n_1_737_4062), .ZN(
      n_1_737_2413));
   INV_X1 i_1_737_2646 (.A(n_1_737_2415), .ZN(n_1_737_2414));
   OAI21_X1 i_1_737_2647 (.A(n_1_737_2416), .B1(n_1_737_5475), .B2(n_1_737_5365), 
      .ZN(n_1_737_2415));
   OAI221_X1 i_1_737_2648 (.A(n_1_737_2417), .B1(n_1_737_4911), .B2(n_1_737_3022), 
      .C1(n_1_737_795), .C2(n_1_737_5366), .ZN(n_1_737_2416));
   NAND2_X1 i_1_737_2649 (.A1(\out_bs[4] [6]), .A2(n_1_737_4073), .ZN(
      n_1_737_2417));
   OAI21_X1 i_1_737_2650 (.A(n_1_737_2419), .B1(n_1_737_5476), .B2(n_1_737_5336), 
      .ZN(n_1_737_2418));
   OAI22_X1 i_1_737_2651 (.A1(n_1_737_4904), .A2(n_1_737_3018), .B1(n_1_737_791), 
      .B2(n_1_737_5337), .ZN(n_1_737_2419));
   NOR3_X1 i_1_737_2652 (.A1(n_1_737_4916), .A2(n_1_737_3083), .A3(n_1_737_790), 
      .ZN(n_232));
   OAI21_X1 i_1_737_2653 (.A(n_1_737_790), .B1(n_1_737_4916), .B2(n_1_737_3083), 
      .ZN(n_233));
   NOR3_X1 i_1_737_2654 (.A1(n_1_737_4923), .A2(n_1_737_3109), .A3(n_1_737_789), 
      .ZN(n_234));
   OAI21_X1 i_1_737_2655 (.A(n_1_737_789), .B1(n_1_737_4923), .B2(n_1_737_3109), 
      .ZN(n_235));
   OAI211_X1 i_1_737_2656 (.A(n_1_737_2433), .B(n_1_737_2420), .C1(n_1_737_784), 
      .C2(n_1_737_2435), .ZN(n_236));
   NOR4_X1 i_1_737_2657 (.A1(n_1_737_2424), .A2(n_1_737_2421), .A3(n_1_737_2427), 
      .A4(n_1_737_2430), .ZN(n_1_737_2420));
   INV_X1 i_1_737_2658 (.A(n_1_737_2422), .ZN(n_1_737_2421));
   OAI21_X1 i_1_737_2659 (.A(n_1_737_2423), .B1(n_1_737_5478), .B2(n_1_737_5297), 
      .ZN(n_1_737_2422));
   OAI22_X1 i_1_737_2660 (.A1(n_1_737_4932), .A2(n_1_737_3015), .B1(n_1_737_785), 
      .B2(n_1_737_5298), .ZN(n_1_737_2423));
   AOI21_X1 i_1_737_2661 (.A(n_1_737_2425), .B1(n_1_737_787), .B2(n_1_737_5190), 
      .ZN(n_1_737_2424));
   INV_X1 i_1_737_2662 (.A(n_1_737_2426), .ZN(n_1_737_2425));
   OAI22_X1 i_1_737_2663 (.A1(n_1_737_4939), .A2(n_1_737_3005), .B1(n_1_737_787), 
      .B2(n_1_737_5190), .ZN(n_1_737_2426));
   AOI21_X1 i_1_737_2664 (.A(n_1_737_2428), .B1(n_1_737_786), .B2(n_1_737_5236), 
      .ZN(n_1_737_2427));
   INV_X1 i_1_737_2665 (.A(n_1_737_2429), .ZN(n_1_737_2428));
   OAI22_X1 i_1_737_2666 (.A1(n_1_737_4953), .A2(n_1_737_3010), .B1(n_1_737_786), 
      .B2(n_1_737_5236), .ZN(n_1_737_2429));
   INV_X1 i_1_737_2667 (.A(n_1_737_2431), .ZN(n_1_737_2430));
   OAI21_X1 i_1_737_2668 (.A(n_1_737_2432), .B1(n_1_737_5477), .B2(n_1_737_5365), 
      .ZN(n_1_737_2431));
   OAI22_X1 i_1_737_2669 (.A1(n_1_737_4960), .A2(n_1_737_3022), .B1(n_1_737_788), 
      .B2(n_1_737_5366), .ZN(n_1_737_2432));
   INV_X1 i_1_737_2670 (.A(n_1_737_2434), .ZN(n_1_737_2433));
   AOI21_X1 i_1_737_2671 (.A(n_1_737_5337), .B1(n_1_737_784), .B2(n_1_737_2435), 
      .ZN(n_1_737_2434));
   NAND2_X1 i_1_737_2672 (.A1(n_1_737_4945), .A2(n_1_737_3019), .ZN(n_1_737_2435));
   NOR2_X1 i_1_737_2673 (.A1(n_1_737_783), .A2(n_1_737_2436), .ZN(n_237));
   NAND2_X1 i_1_737_2674 (.A1(n_1_737_783), .A2(n_1_737_2436), .ZN(n_238));
   NAND2_X1 i_1_737_2675 (.A1(n_1_737_3882), .A2(n_1_737_3084), .ZN(n_1_737_2436));
   NOR2_X1 i_1_737_2676 (.A1(n_1_737_782), .A2(n_1_737_2437), .ZN(n_239));
   NAND2_X1 i_1_737_2677 (.A1(n_1_737_782), .A2(n_1_737_2437), .ZN(n_240));
   NAND2_X1 i_1_737_2678 (.A1(n_1_737_4963), .A2(n_1_737_3110), .ZN(n_1_737_2437));
   NAND3_X1 i_1_737_2679 (.A1(n_1_737_2440), .A2(n_1_737_2438), .A3(n_1_737_2450), 
      .ZN(n_241));
   AOI211_X1 i_1_737_2680 (.A(n_1_737_2447), .B(n_1_737_2443), .C1(n_1_737_2446), 
      .C2(n_1_737_2445), .ZN(n_1_737_2438));
   INV_X1 i_1_737_2681 (.A(n_1_737_2440), .ZN(n_1_737_2439));
   OAI21_X1 i_1_737_2682 (.A(n_1_737_2441), .B1(n_1_737_5480), .B2(n_1_737_5189), 
      .ZN(n_1_737_2440));
   OAI21_X1 i_1_737_2683 (.A(n_1_737_2442), .B1(n_1_737_780), .B2(n_1_737_5190), 
      .ZN(n_1_737_2441));
   OAI21_X1 i_1_737_2684 (.A(\out_bs[3] [6]), .B1(n_1_737_4039), .B2(
      n_1_737_3896), .ZN(n_1_737_2442));
   AOI21_X1 i_1_737_2685 (.A(n_1_737_2444), .B1(n_1_737_779), .B2(n_1_737_5236), 
      .ZN(n_1_737_2443));
   AOI22_X1 i_1_737_2686 (.A1(\out_bs[2] [6]), .A2(n_1_737_3908), .B1(
      n_1_737_5481), .B2(n_1_737_5235), .ZN(n_1_737_2444));
   NAND2_X1 i_1_737_2687 (.A1(n_1_737_777), .A2(n_1_737_5337), .ZN(n_1_737_2445));
   OAI22_X1 i_1_737_2688 (.A1(n_1_737_5671), .A2(n_1_737_3890), .B1(n_1_737_777), 
      .B2(n_1_737_5337), .ZN(n_1_737_2446));
   INV_X1 i_1_737_2689 (.A(n_1_737_2448), .ZN(n_1_737_2447));
   OAI21_X1 i_1_737_2690 (.A(n_1_737_2449), .B1(n_1_737_5482), .B2(n_1_737_5297), 
      .ZN(n_1_737_2448));
   OAI22_X1 i_1_737_2691 (.A1(n_1_737_5664), .A2(n_1_737_3903), .B1(n_1_737_778), 
      .B2(n_1_737_5298), .ZN(n_1_737_2449));
   OAI21_X1 i_1_737_2692 (.A(n_1_737_2451), .B1(n_1_737_5479), .B2(n_1_737_5365), 
      .ZN(n_1_737_2450));
   OAI22_X1 i_1_737_2693 (.A1(n_1_737_5625), .A2(n_1_737_3914), .B1(n_1_737_781), 
      .B2(n_1_737_5366), .ZN(n_1_737_2451));
   NOR3_X1 i_1_737_2694 (.A1(n_1_737_5607), .A2(n_1_737_4011), .A3(n_1_737_776), 
      .ZN(n_242));
   OAI21_X1 i_1_737_2695 (.A(n_1_737_776), .B1(n_1_737_5607), .B2(n_1_737_4011), 
      .ZN(n_243));
   NOR2_X1 i_1_737_2696 (.A1(n_1_737_775), .A2(n_1_737_2452), .ZN(n_244));
   NAND2_X1 i_1_737_2697 (.A1(n_1_737_775), .A2(n_1_737_2452), .ZN(n_245));
   NAND2_X1 i_1_737_2698 (.A1(n_844), .A2(n_1_737_4020), .ZN(n_1_737_2452));
   OR4_X1 i_1_737_2699 (.A1(n_1_737_2455), .A2(n_1_737_2453), .A3(n_1_737_2463), 
      .A4(n_1_737_2466), .ZN(n_246));
   OAI211_X1 i_1_737_2700 (.A(n_1_737_2454), .B(n_1_737_2461), .C1(n_1_737_770), 
      .C2(n_1_737_2458), .ZN(n_1_737_2453));
   OAI21_X1 i_1_737_2701 (.A(n_1_737_5336), .B1(n_1_737_5485), .B2(n_1_737_2459), 
      .ZN(n_1_737_2454));
   AOI21_X1 i_1_737_2702 (.A(n_1_737_2456), .B1(n_1_737_772), .B2(n_1_737_5236), 
      .ZN(n_1_737_2455));
   INV_X1 i_1_737_2703 (.A(n_1_737_2457), .ZN(n_1_737_2456));
   OAI22_X1 i_1_737_2704 (.A1(n_1_737_5651), .A2(n_1_737_4061), .B1(n_1_737_772), 
      .B2(n_1_737_5236), .ZN(n_1_737_2457));
   INV_X1 i_1_737_2705 (.A(n_1_737_2459), .ZN(n_1_737_2458));
   NOR2_X1 i_1_737_2706 (.A1(n_1_737_5671), .A2(n_1_737_4028), .ZN(n_1_737_2459));
   INV_X1 i_1_737_2707 (.A(n_1_737_2461), .ZN(n_1_737_2460));
   OAI21_X1 i_1_737_2708 (.A(n_1_737_2462), .B1(n_1_737_5484), .B2(n_1_737_5297), 
      .ZN(n_1_737_2461));
   OAI22_X1 i_1_737_2709 (.A1(n_1_737_5664), .A2(n_1_737_4048), .B1(n_1_737_771), 
      .B2(n_1_737_5298), .ZN(n_1_737_2462));
   INV_X1 i_1_737_2710 (.A(n_1_737_2464), .ZN(n_1_737_2463));
   OAI21_X1 i_1_737_2711 (.A(n_1_737_2465), .B1(n_1_737_5483), .B2(n_1_737_5189), 
      .ZN(n_1_737_2464));
   OAI22_X1 i_1_737_2712 (.A1(n_1_737_5638), .A2(n_1_737_4038), .B1(n_1_737_773), 
      .B2(n_1_737_5190), .ZN(n_1_737_2465));
   AOI21_X1 i_1_737_2713 (.A(n_1_737_2467), .B1(n_1_737_774), .B2(n_1_737_5366), 
      .ZN(n_1_737_2466));
   INV_X1 i_1_737_2714 (.A(n_1_737_2468), .ZN(n_1_737_2467));
   OAI22_X1 i_1_737_2715 (.A1(n_1_737_5625), .A2(n_1_737_4072), .B1(n_1_737_774), 
      .B2(n_1_737_5366), .ZN(n_1_737_2468));
   NOR2_X1 i_1_737_2716 (.A1(n_1_737_769), .A2(n_1_737_2469), .ZN(n_247));
   NAND2_X1 i_1_737_2717 (.A1(n_1_737_769), .A2(n_1_737_2469), .ZN(n_248));
   OAI21_X1 i_1_737_2718 (.A(\out_bs[6] [6]), .B1(n_1_737_4012), .B2(
      n_1_737_3940), .ZN(n_1_737_2469));
   NOR2_X1 i_1_737_2719 (.A1(n_1_737_768), .A2(n_1_737_2470), .ZN(n_249));
   NAND2_X1 i_1_737_2720 (.A1(n_1_737_768), .A2(n_1_737_2470), .ZN(n_250));
   OAI21_X1 i_1_737_2721 (.A(n_844), .B1(n_1_737_4020), .B2(n_1_737_3945), 
      .ZN(n_1_737_2470));
   OAI211_X1 i_1_737_2722 (.A(n_1_737_2471), .B(n_1_737_2486), .C1(n_1_737_763), 
      .C2(n_1_737_2482), .ZN(n_251));
   NOR3_X1 i_1_737_2723 (.A1(n_1_737_2475), .A2(n_1_737_2472), .A3(n_1_737_2478), 
      .ZN(n_1_737_2471));
   AOI21_X1 i_1_737_2724 (.A(n_1_737_2473), .B1(n_1_737_766), .B2(n_1_737_5190), 
      .ZN(n_1_737_2472));
   INV_X1 i_1_737_2725 (.A(n_1_737_2474), .ZN(n_1_737_2473));
   OAI22_X1 i_1_737_2726 (.A1(n_1_737_5638), .A2(n_1_737_3957), .B1(n_1_737_766), 
      .B2(n_1_737_5190), .ZN(n_1_737_2474));
   AOI21_X1 i_1_737_2727 (.A(n_1_737_2476), .B1(n_1_737_765), .B2(n_1_737_5236), 
      .ZN(n_1_737_2475));
   INV_X1 i_1_737_2728 (.A(n_1_737_2477), .ZN(n_1_737_2476));
   OAI22_X1 i_1_737_2729 (.A1(n_1_737_5651), .A2(n_1_737_3951), .B1(n_1_737_765), 
      .B2(n_1_737_5236), .ZN(n_1_737_2477));
   OAI21_X1 i_1_737_2730 (.A(n_1_737_2480), .B1(n_1_737_5337), .B2(n_1_737_2483), 
      .ZN(n_1_737_2478));
   INV_X1 i_1_737_2731 (.A(n_1_737_2480), .ZN(n_1_737_2479));
   OAI21_X1 i_1_737_2732 (.A(n_1_737_2481), .B1(n_1_737_5487), .B2(n_1_737_5297), 
      .ZN(n_1_737_2480));
   OAI22_X1 i_1_737_2733 (.A1(n_1_737_5664), .A2(n_1_737_3970), .B1(n_1_737_764), 
      .B2(n_1_737_5298), .ZN(n_1_737_2481));
   NOR2_X1 i_1_737_2734 (.A1(n_1_737_5336), .A2(n_1_737_2484), .ZN(n_1_737_2482));
   INV_X1 i_1_737_2735 (.A(n_1_737_2484), .ZN(n_1_737_2483));
   NOR2_X1 i_1_737_2736 (.A1(n_1_737_5671), .A2(n_1_737_3963), .ZN(n_1_737_2484));
   INV_X1 i_1_737_2737 (.A(n_1_737_2486), .ZN(n_1_737_2485));
   OAI21_X1 i_1_737_2738 (.A(n_1_737_2487), .B1(n_1_737_5486), .B2(n_1_737_5365), 
      .ZN(n_1_737_2486));
   OAI22_X1 i_1_737_2739 (.A1(n_1_737_5625), .A2(n_1_737_3977), .B1(n_1_737_767), 
      .B2(n_1_737_5366), .ZN(n_1_737_2487));
   NOR3_X1 i_1_737_2740 (.A1(n_1_737_5072), .A2(n_1_737_3109), .A3(n_1_737_761), 
      .ZN(n_252));
   OAI21_X1 i_1_737_2741 (.A(n_1_737_761), .B1(n_1_737_5072), .B2(n_1_737_3109), 
      .ZN(n_253));
   OAI211_X1 i_1_737_2742 (.A(n_1_737_2501), .B(n_1_737_2488), .C1(n_1_737_756), 
      .C2(n_1_737_2503), .ZN(n_254));
   NOR4_X1 i_1_737_2743 (.A1(n_1_737_2492), .A2(n_1_737_2489), .A3(n_1_737_2495), 
      .A4(n_1_737_2498), .ZN(n_1_737_2488));
   INV_X1 i_1_737_2744 (.A(n_1_737_2490), .ZN(n_1_737_2489));
   OAI21_X1 i_1_737_2745 (.A(n_1_737_2491), .B1(n_1_737_5489), .B2(n_1_737_5297), 
      .ZN(n_1_737_2490));
   OAI22_X1 i_1_737_2746 (.A1(n_1_737_5109), .A2(n_1_737_3015), .B1(n_1_737_757), 
      .B2(n_1_737_5298), .ZN(n_1_737_2491));
   INV_X1 i_1_737_2747 (.A(n_1_737_2493), .ZN(n_1_737_2492));
   OAI21_X1 i_1_737_2748 (.A(n_1_737_2494), .B1(n_1_737_5488), .B2(n_1_737_5189), 
      .ZN(n_1_737_2493));
   OAI22_X1 i_1_737_2749 (.A1(n_1_737_5120), .A2(n_1_737_3005), .B1(n_1_737_759), 
      .B2(n_1_737_5190), .ZN(n_1_737_2494));
   AOI21_X1 i_1_737_2750 (.A(n_1_737_2496), .B1(n_1_737_758), .B2(n_1_737_5236), 
      .ZN(n_1_737_2495));
   INV_X1 i_1_737_2751 (.A(n_1_737_2497), .ZN(n_1_737_2496));
   OAI22_X1 i_1_737_2752 (.A1(n_1_737_5093), .A2(n_1_737_3010), .B1(n_1_737_758), 
      .B2(n_1_737_5236), .ZN(n_1_737_2497));
   AOI21_X1 i_1_737_2753 (.A(n_1_737_2499), .B1(n_1_737_760), .B2(n_1_737_5366), 
      .ZN(n_1_737_2498));
   INV_X1 i_1_737_2754 (.A(n_1_737_2500), .ZN(n_1_737_2499));
   OAI22_X1 i_1_737_2755 (.A1(n_1_737_5128), .A2(n_1_737_3022), .B1(n_1_737_760), 
      .B2(n_1_737_5366), .ZN(n_1_737_2500));
   INV_X1 i_1_737_2756 (.A(n_1_737_2502), .ZN(n_1_737_2501));
   AOI21_X1 i_1_737_2757 (.A(n_1_737_5337), .B1(n_1_737_756), .B2(n_1_737_2503), 
      .ZN(n_1_737_2502));
   OR2_X1 i_1_737_2758 (.A1(n_1_737_5079), .A2(n_1_737_3018), .ZN(n_1_737_2503));
   NOR2_X1 i_1_737_2759 (.A1(n_1_737_755), .A2(n_1_737_2504), .ZN(n_255));
   NAND2_X1 i_1_737_2760 (.A1(n_1_737_755), .A2(n_1_737_2504), .ZN(n_256));
   OR2_X1 i_1_737_2761 (.A1(n_1_737_4013), .A2(n_1_737_3083), .ZN(n_1_737_2504));
   NOR2_X1 i_1_737_2762 (.A1(n_1_737_754), .A2(n_1_737_2505), .ZN(n_257));
   NAND2_X1 i_1_737_2763 (.A1(n_1_737_754), .A2(n_1_737_2505), .ZN(n_258));
   OAI21_X1 i_1_737_2764 (.A(n_844), .B1(n_1_737_4021), .B2(n_1_737_4020), 
      .ZN(n_1_737_2505));
   NAND4_X1 i_1_737_2765 (.A1(n_1_737_2510), .A2(n_1_737_2508), .A3(n_1_737_2506), 
      .A4(n_1_737_2517), .ZN(n_259));
   OAI21_X1 i_1_737_2766 (.A(n_1_737_2507), .B1(n_1_737_5491), .B2(n_1_737_5189), 
      .ZN(n_1_737_2506));
   OAI22_X1 i_1_737_2767 (.A1(n_1_737_5638), .A2(n_1_737_4037), .B1(n_1_737_752), 
      .B2(n_1_737_5190), .ZN(n_1_737_2507));
   OAI21_X1 i_1_737_2768 (.A(n_1_737_2509), .B1(n_1_737_5492), .B2(n_1_737_5235), 
      .ZN(n_1_737_2508));
   OAI22_X1 i_1_737_2769 (.A1(n_1_737_5651), .A2(n_1_737_4060), .B1(n_1_737_751), 
      .B2(n_1_737_5236), .ZN(n_1_737_2509));
   AOI211_X1 i_1_737_2770 (.A(n_1_737_2511), .B(n_1_737_2514), .C1(n_1_737_5336), 
      .C2(n_1_737_2515), .ZN(n_1_737_2510));
   INV_X1 i_1_737_2771 (.A(n_1_737_2512), .ZN(n_1_737_2511));
   OAI21_X1 i_1_737_2772 (.A(n_1_737_2513), .B1(n_1_737_5493), .B2(n_1_737_5297), 
      .ZN(n_1_737_2512));
   OAI22_X1 i_1_737_2773 (.A1(n_1_737_5664), .A2(n_1_737_4047), .B1(n_1_737_750), 
      .B2(n_1_737_5298), .ZN(n_1_737_2513));
   AOI21_X1 i_1_737_2774 (.A(n_1_737_749), .B1(n_1_737_5337), .B2(n_1_737_2516), 
      .ZN(n_1_737_2514));
   INV_X1 i_1_737_2775 (.A(n_1_737_2516), .ZN(n_1_737_2515));
   OAI211_X1 i_1_737_2776 (.A(\out_bs[0] [5]), .B(\out_bs[0] [6]), .C1(
      \out_bs[0] [4]), .C2(n_1_737_5326), .ZN(n_1_737_2516));
   OAI21_X1 i_1_737_2777 (.A(n_1_737_2518), .B1(n_1_737_5490), .B2(n_1_737_5365), 
      .ZN(n_1_737_2517));
   OAI22_X1 i_1_737_2778 (.A1(n_1_737_5625), .A2(n_1_737_4071), .B1(n_1_737_753), 
      .B2(n_1_737_5366), .ZN(n_1_737_2518));
   NAND4_X1 i_1_737_2779 (.A1(n_1_737_2522), .A2(n_1_737_2519), .A3(n_1_737_2531), 
      .A4(n_1_737_2524), .ZN(n_260));
   AOI211_X1 i_1_737_2780 (.A(n_1_737_2526), .B(n_1_737_2529), .C1(n_1_737_2521), 
      .C2(n_1_737_2520), .ZN(n_1_737_2519));
   NAND2_X1 i_1_737_2781 (.A1(n_1_737_742), .A2(n_1_737_5337), .ZN(n_1_737_2520));
   OAI21_X1 i_1_737_2782 (.A(n_1_737_3018), .B1(n_1_737_742), .B2(n_1_737_5337), 
      .ZN(n_1_737_2521));
   OAI21_X1 i_1_737_2783 (.A(n_1_737_2523), .B1(n_1_737_5495), .B2(n_1_737_5189), 
      .ZN(n_1_737_2522));
   OAI21_X1 i_1_737_2784 (.A(n_1_737_3005), .B1(n_1_737_745), .B2(n_1_737_5190), 
      .ZN(n_1_737_2523));
   OAI21_X1 i_1_737_2785 (.A(n_1_737_2525), .B1(n_1_737_5602), .B2(n_1_737_5494), 
      .ZN(n_1_737_2524));
   OAI21_X1 i_1_737_2786 (.A(n_1_737_3109), .B1(n_1089), .B2(n_1_737_747), 
      .ZN(n_1_737_2525));
   OAI22_X1 i_1_737_2787 (.A1(n_1_737_743), .A2(n_1_737_3015), .B1(n_1_737_5298), 
      .B2(n_1_737_2527), .ZN(n_1_737_2526));
   AND2_X1 i_1_737_2788 (.A1(n_1_737_743), .A2(n_1_737_3015), .ZN(n_1_737_2527));
   INV_X1 i_1_737_2789 (.A(n_1_737_2529), .ZN(n_1_737_2528));
   OAI22_X1 i_1_737_2790 (.A1(n_1_737_744), .A2(n_1_737_3010), .B1(n_1_737_5236), 
      .B2(n_1_737_2530), .ZN(n_1_737_2529));
   AND2_X1 i_1_737_2791 (.A1(n_1_737_744), .A2(n_1_737_3010), .ZN(n_1_737_2530));
   INV_X1 i_1_737_2792 (.A(n_1_737_2532), .ZN(n_1_737_2531));
   OAI22_X1 i_1_737_2793 (.A1(n_1_737_746), .A2(n_1_737_3022), .B1(n_1_737_5366), 
      .B2(n_1_737_2533), .ZN(n_1_737_2532));
   AND2_X1 i_1_737_2794 (.A1(n_1_737_746), .A2(n_1_737_3022), .ZN(n_1_737_2533));
   NOR2_X1 i_1_737_2795 (.A1(n_1_737_741), .A2(n_1_737_2534), .ZN(n_261));
   NAND2_X1 i_1_737_2796 (.A1(n_1_737_741), .A2(n_1_737_2534), .ZN(n_262));
   INV_X1 i_1_737_2797 (.A(n_1_737_2535), .ZN(n_1_737_2534));
   AOI21_X1 i_1_737_2798 (.A(n_1_737_2591), .B1(n_1_737_5606), .B2(n_1_737_3943), 
      .ZN(n_1_737_2535));
   NOR2_X1 i_1_737_2799 (.A1(n_1_737_740), .A2(n_1_737_2536), .ZN(n_263));
   NAND2_X1 i_1_737_2800 (.A1(n_1_737_740), .A2(n_1_737_2536), .ZN(n_264));
   OAI21_X1 i_1_737_2801 (.A(n_844), .B1(n_845), .B2(n_1_737_4092), .ZN(
      n_1_737_2536));
   OR4_X1 i_1_737_2802 (.A1(n_1_737_2543), .A2(n_1_737_2540), .A3(n_1_737_2537), 
      .A4(n_1_737_2550), .ZN(n_265));
   INV_X1 i_1_737_2803 (.A(n_1_737_2538), .ZN(n_1_737_2537));
   OAI21_X1 i_1_737_2804 (.A(n_1_737_2539), .B1(n_1_737_5496), .B2(n_1_737_5189), 
      .ZN(n_1_737_2538));
   OAI22_X1 i_1_737_2805 (.A1(n_1_737_5638), .A2(n_1_737_4112), .B1(n_1_737_738), 
      .B2(n_1_737_5190), .ZN(n_1_737_2539));
   AOI21_X1 i_1_737_2806 (.A(n_1_737_2541), .B1(n_1_737_737), .B2(n_1_737_5236), 
      .ZN(n_1_737_2540));
   INV_X1 i_1_737_2807 (.A(n_1_737_2542), .ZN(n_1_737_2541));
   OAI22_X1 i_1_737_2808 (.A1(n_1_737_5651), .A2(n_1_737_4107), .B1(n_1_737_737), 
      .B2(n_1_737_5236), .ZN(n_1_737_2542));
   OAI211_X1 i_1_737_2809 (.A(n_1_737_2545), .B(n_1_737_2547), .C1(n_1_737_5337), 
      .C2(n_1_737_2549), .ZN(n_1_737_2543));
   INV_X1 i_1_737_2810 (.A(n_1_737_2545), .ZN(n_1_737_2544));
   OAI21_X1 i_1_737_2811 (.A(n_1_737_2546), .B1(n_1_737_5497), .B2(n_1_737_5297), 
      .ZN(n_1_737_2545));
   OAI22_X1 i_1_737_2812 (.A1(n_1_737_5664), .A2(n_1_737_4117), .B1(n_1_737_736), 
      .B2(n_1_737_5298), .ZN(n_1_737_2546));
   INV_X1 i_1_737_2813 (.A(n_1_737_2548), .ZN(n_1_737_2547));
   AOI21_X1 i_1_737_2814 (.A(n_1_737_735), .B1(n_1_737_5337), .B2(n_1_737_2549), 
      .ZN(n_1_737_2548));
   OAI21_X1 i_1_737_2815 (.A(\out_bs[0] [6]), .B1(\out_bs[0] [5]), .B2(
      n_1_737_4096), .ZN(n_1_737_2549));
   AOI21_X1 i_1_737_2816 (.A(n_1_737_2551), .B1(n_1_737_739), .B2(n_1_737_5366), 
      .ZN(n_1_737_2550));
   INV_X1 i_1_737_2817 (.A(n_1_737_2552), .ZN(n_1_737_2551));
   OAI22_X1 i_1_737_2818 (.A1(n_1_737_5625), .A2(n_1_737_4100), .B1(n_1_737_739), 
      .B2(n_1_737_5366), .ZN(n_1_737_2552));
   NOR2_X1 i_1_737_2819 (.A1(n_1_737_734), .A2(n_1_737_2553), .ZN(n_266));
   NAND2_X1 i_1_737_2820 (.A1(n_1_737_734), .A2(n_1_737_2553), .ZN(n_267));
   OAI21_X1 i_1_737_2821 (.A(n_1_737_2666), .B1(n_1_737_4921), .B2(n_1_737_3084), 
      .ZN(n_1_737_2553));
   NOR2_X1 i_1_737_2822 (.A1(n_1_737_733), .A2(n_1_737_2554), .ZN(n_268));
   NAND2_X1 i_1_737_2823 (.A1(n_1_737_733), .A2(n_1_737_2554), .ZN(n_269));
   OAI21_X1 i_1_737_2824 (.A(n_844), .B1(n_845), .B2(n_1_737_4120), .ZN(
      n_1_737_2554));
   OR4_X1 i_1_737_2825 (.A1(n_1_737_2556), .A2(n_1_737_2555), .A3(n_1_737_2559), 
      .A4(n_1_737_2569), .ZN(n_270));
   AOI21_X1 i_1_737_2826 (.A(n_1_737_728), .B1(n_1_737_5337), .B2(n_1_737_2560), 
      .ZN(n_1_737_2555));
   AOI21_X1 i_1_737_2827 (.A(n_1_737_2557), .B1(n_1_737_730), .B2(n_1_737_5236), 
      .ZN(n_1_737_2556));
   INV_X1 i_1_737_2828 (.A(n_1_737_2558), .ZN(n_1_737_2557));
   OAI22_X1 i_1_737_2829 (.A1(n_1_737_5651), .A2(n_1_737_4142), .B1(n_1_737_730), 
      .B2(n_1_737_5236), .ZN(n_1_737_2558));
   OAI211_X1 i_1_737_2830 (.A(n_1_737_2562), .B(n_1_737_2566), .C1(n_1_737_5337), 
      .C2(n_1_737_2560), .ZN(n_1_737_2559));
   OAI21_X1 i_1_737_2831 (.A(\out_bs[0] [6]), .B1(\out_bs[0] [5]), .B2(
      n_1_737_4138), .ZN(n_1_737_2560));
   INV_X1 i_1_737_2832 (.A(n_1_737_2562), .ZN(n_1_737_2561));
   OAI21_X1 i_1_737_2833 (.A(n_1_737_2563), .B1(n_1_737_5500), .B2(n_1_737_5297), 
      .ZN(n_1_737_2562));
   OAI21_X1 i_1_737_2834 (.A(n_1_737_2564), .B1(n_1_737_729), .B2(n_1_737_5298), 
      .ZN(n_1_737_2563));
   OAI21_X1 i_1_737_2835 (.A(n_1_737_2673), .B1(\out_bs[1] [5]), .B2(
      n_1_737_4933), .ZN(n_1_737_2564));
   INV_X1 i_1_737_2836 (.A(n_1_737_2566), .ZN(n_1_737_2565));
   OAI21_X1 i_1_737_2837 (.A(n_1_737_2567), .B1(n_1_737_5499), .B2(n_1_737_5189), 
      .ZN(n_1_737_2566));
   OAI21_X1 i_1_737_2838 (.A(n_1_737_2568), .B1(n_1_737_731), .B2(n_1_737_5190), 
      .ZN(n_1_737_2567));
   OAI21_X1 i_1_737_2839 (.A(\out_bs[3] [6]), .B1(\out_bs[3] [5]), .B2(
      n_1_737_4132), .ZN(n_1_737_2568));
   INV_X1 i_1_737_2840 (.A(n_1_737_2570), .ZN(n_1_737_2569));
   OAI21_X1 i_1_737_2841 (.A(n_1_737_2571), .B1(n_1_737_5498), .B2(n_1_737_5365), 
      .ZN(n_1_737_2570));
   OAI22_X1 i_1_737_2842 (.A1(n_1_737_5625), .A2(n_1_737_4149), .B1(n_1_737_732), 
      .B2(n_1_737_5366), .ZN(n_1_737_2571));
   NOR2_X1 i_1_737_2843 (.A1(n_1_737_727), .A2(n_1_737_2572), .ZN(n_271));
   NAND2_X1 i_1_737_2844 (.A1(n_1_737_727), .A2(n_1_737_2572), .ZN(n_272));
   OAI21_X1 i_1_737_2845 (.A(\out_bs[6] [6]), .B1(\out_bs[6] [5]), .B2(
      n_1_737_3195), .ZN(n_1_737_2572));
   NOR2_X1 i_1_737_2846 (.A1(n_1_737_726), .A2(n_1_737_2573), .ZN(n_273));
   NAND2_X1 i_1_737_2847 (.A1(n_1_737_726), .A2(n_1_737_2573), .ZN(n_274));
   OAI21_X1 i_1_737_2848 (.A(n_844), .B1(n_845), .B2(n_1_737_4153), .ZN(
      n_1_737_2573));
   OR4_X1 i_1_737_2849 (.A1(n_1_737_2580), .A2(n_1_737_2577), .A3(n_1_737_2574), 
      .A4(n_1_737_2587), .ZN(n_275));
   AOI21_X1 i_1_737_2850 (.A(n_1_737_2575), .B1(n_1_737_724), .B2(n_1_737_5190), 
      .ZN(n_1_737_2574));
   INV_X1 i_1_737_2851 (.A(n_1_737_2576), .ZN(n_1_737_2575));
   OAI22_X1 i_1_737_2852 (.A1(n_1_737_5638), .A2(n_1_737_4163), .B1(n_1_737_724), 
      .B2(n_1_737_5190), .ZN(n_1_737_2576));
   INV_X1 i_1_737_2853 (.A(n_1_737_2578), .ZN(n_1_737_2577));
   OAI21_X1 i_1_737_2854 (.A(n_1_737_2579), .B1(n_1_737_5501), .B2(n_1_737_5235), 
      .ZN(n_1_737_2578));
   OAI22_X1 i_1_737_2855 (.A1(n_1_737_5651), .A2(n_1_737_4177), .B1(n_1_737_723), 
      .B2(n_1_737_5236), .ZN(n_1_737_2579));
   OAI211_X1 i_1_737_2856 (.A(n_1_737_2582), .B(n_1_737_2584), .C1(n_1_737_5337), 
      .C2(n_1_737_2586), .ZN(n_1_737_2580));
   INV_X1 i_1_737_2857 (.A(n_1_737_2582), .ZN(n_1_737_2581));
   OAI21_X1 i_1_737_2858 (.A(n_1_737_2583), .B1(n_1_737_5502), .B2(n_1_737_5297), 
      .ZN(n_1_737_2582));
   OAI22_X1 i_1_737_2859 (.A1(n_1_737_5664), .A2(n_1_737_4171), .B1(n_1_737_722), 
      .B2(n_1_737_5298), .ZN(n_1_737_2583));
   INV_X1 i_1_737_2860 (.A(n_1_737_2585), .ZN(n_1_737_2584));
   AOI21_X1 i_1_737_2861 (.A(n_1_737_721), .B1(n_1_737_5337), .B2(n_1_737_2586), 
      .ZN(n_1_737_2585));
   OAI21_X1 i_1_737_2862 (.A(\out_bs[0] [6]), .B1(\out_bs[0] [5]), .B2(
      n_1_737_4159), .ZN(n_1_737_2586));
   AOI21_X1 i_1_737_2863 (.A(n_1_737_2588), .B1(n_1_737_725), .B2(n_1_737_5366), 
      .ZN(n_1_737_2587));
   INV_X1 i_1_737_2864 (.A(n_1_737_2589), .ZN(n_1_737_2588));
   OAI21_X1 i_1_737_2865 (.A(n_1_737_2590), .B1(n_1_737_725), .B2(n_1_737_5366), 
      .ZN(n_1_737_2589));
   OAI21_X1 i_1_737_2866 (.A(n_1_737_2609), .B1(\out_bs[4] [5]), .B2(
      n_1_737_5404), .ZN(n_1_737_2590));
   NOR2_X1 i_1_737_2867 (.A1(n_1_737_720), .A2(n_1_737_2591), .ZN(n_276));
   NAND2_X1 i_1_737_2868 (.A1(n_1_737_720), .A2(n_1_737_2591), .ZN(n_277));
   OAI21_X1 i_1_737_2869 (.A(\out_bs[6] [6]), .B1(\out_bs[6] [5]), .B2(
      n_1_737_3223), .ZN(n_1_737_2591));
   NAND3_X1 i_1_737_2870 (.A1(n_1_737_2606), .A2(n_1_737_2604), .A3(n_1_737_2592), 
      .ZN(n_278));
   NOR3_X1 i_1_737_2871 (.A1(n_1_737_2594), .A2(n_1_737_2593), .A3(n_1_737_2597), 
      .ZN(n_1_737_2592));
   AOI21_X1 i_1_737_2872 (.A(n_1_737_5337), .B1(n_1_737_714), .B2(n_1_737_2598), 
      .ZN(n_1_737_2593));
   INV_X1 i_1_737_2873 (.A(n_1_737_2595), .ZN(n_1_737_2594));
   OAI21_X1 i_1_737_2874 (.A(n_1_737_2596), .B1(n_1_737_5505), .B2(n_1_737_5297), 
      .ZN(n_1_737_2595));
   OAI221_X1 i_1_737_2875 (.A(n_1_737_3015), .B1(n_1_737_5664), .B2(n_1_737_4218), 
      .C1(n_1_737_715), .C2(n_1_737_5298), .ZN(n_1_737_2596));
   OAI211_X1 i_1_737_2876 (.A(n_1_737_2599), .B(n_1_737_2602), .C1(n_1_737_714), 
      .C2(n_1_737_2598), .ZN(n_1_737_2597));
   OAI21_X1 i_1_737_2877 (.A(\out_bs[0] [6]), .B1(\out_bs[0] [5]), .B2(
      n_1_737_4243), .ZN(n_1_737_2598));
   INV_X1 i_1_737_2878 (.A(n_1_737_2600), .ZN(n_1_737_2599));
   OAI22_X1 i_1_737_2879 (.A1(n_1089), .A2(n_1_737_719), .B1(n_1_737_2611), 
      .B2(n_1_737_2601), .ZN(n_1_737_2600));
   AND2_X1 i_1_737_2880 (.A1(n_1089), .A2(n_1_737_719), .ZN(n_1_737_2601));
   OAI21_X1 i_1_737_2881 (.A(n_1_737_2603), .B1(n_1_737_5503), .B2(n_1_737_5189), 
      .ZN(n_1_737_2602));
   OAI221_X1 i_1_737_2882 (.A(n_1_737_3005), .B1(n_1_737_5638), .B2(n_1_737_4225), 
      .C1(n_1_737_717), .C2(n_1_737_5190), .ZN(n_1_737_2603));
   OAI21_X1 i_1_737_2883 (.A(n_1_737_2605), .B1(n_1_737_5504), .B2(n_1_737_5235), 
      .ZN(n_1_737_2604));
   OAI221_X1 i_1_737_2884 (.A(n_1_737_3010), .B1(n_1_737_5651), .B2(n_1_737_4234), 
      .C1(n_1_737_716), .C2(n_1_737_5236), .ZN(n_1_737_2605));
   OAI21_X1 i_1_737_2885 (.A(n_1_737_2607), .B1(n_1_737_5365), .B2(n_1_737_2609), 
      .ZN(n_1_737_2606));
   OAI21_X1 i_1_737_2886 (.A(n_1_737_718), .B1(n_1_737_5366), .B2(n_1_737_2608), 
      .ZN(n_1_737_2607));
   INV_X1 i_1_737_2887 (.A(n_1_737_2609), .ZN(n_1_737_2608));
   NOR2_X1 i_1_737_2888 (.A1(n_1_737_5625), .A2(n_1_737_4252), .ZN(n_1_737_2609));
   NOR2_X1 i_1_737_2889 (.A1(n_1_737_712), .A2(n_1_737_2610), .ZN(n_279));
   NAND2_X1 i_1_737_2890 (.A1(n_1_737_712), .A2(n_1_737_2610), .ZN(n_280));
   OAI21_X1 i_1_737_2891 (.A(n_844), .B1(n_845), .B2(n_1_737_4206), .ZN(
      n_1_737_2610));
   OAI21_X1 i_1_737_2892 (.A(n_844), .B1(n_845), .B2(n_1_737_4209), .ZN(
      n_1_737_2611));
   NAND2_X1 i_1_737_2893 (.A1(n_1_737_2618), .A2(n_1_737_2612), .ZN(n_281));
   AOI21_X1 i_1_737_2894 (.A(n_1_737_2615), .B1(n_1_737_2614), .B2(n_1_737_2613), 
      .ZN(n_1_737_2612));
   NAND2_X1 i_1_737_2895 (.A1(n_1_737_707), .A2(n_1_737_5337), .ZN(n_1_737_2613));
   OAI22_X1 i_1_737_2896 (.A1(n_1_737_5671), .A2(n_1_737_4240), .B1(n_1_737_707), 
      .B2(n_1_737_5337), .ZN(n_1_737_2614));
   OAI22_X1 i_1_737_2897 (.A1(n_1_737_711), .A2(n_1_737_5366), .B1(n_1_737_2617), 
      .B2(n_1_737_2616), .ZN(n_1_737_2615));
   OAI21_X1 i_1_737_2898 (.A(\out_bs[4] [6]), .B1(\out_bs[4] [5]), .B2(
      n_1_737_4249), .ZN(n_1_737_2616));
   AND2_X1 i_1_737_2899 (.A1(n_1_737_711), .A2(n_1_737_5366), .ZN(n_1_737_2617));
   NOR3_X1 i_1_737_2900 (.A1(n_1_737_2623), .A2(n_1_737_2620), .A3(n_1_737_2626), 
      .ZN(n_1_737_2618));
   INV_X1 i_1_737_2901 (.A(n_1_737_2620), .ZN(n_1_737_2619));
   OAI22_X1 i_1_737_2902 (.A1(n_1_737_708), .A2(n_1_737_5298), .B1(n_1_737_2622), 
      .B2(n_1_737_2621), .ZN(n_1_737_2620));
   OAI21_X1 i_1_737_2903 (.A(\out_bs[1] [6]), .B1(\out_bs[1] [5]), .B2(
      n_1_737_4217), .ZN(n_1_737_2621));
   AND2_X1 i_1_737_2904 (.A1(n_1_737_708), .A2(n_1_737_5298), .ZN(n_1_737_2622));
   OAI22_X1 i_1_737_2905 (.A1(n_1_737_709), .A2(n_1_737_5236), .B1(n_1_737_2625), 
      .B2(n_1_737_2624), .ZN(n_1_737_2623));
   OAI21_X1 i_1_737_2906 (.A(\out_bs[2] [6]), .B1(\out_bs[2] [5]), .B2(
      n_1_737_4232), .ZN(n_1_737_2624));
   AND2_X1 i_1_737_2907 (.A1(n_1_737_709), .A2(n_1_737_5236), .ZN(n_1_737_2625));
   OAI22_X1 i_1_737_2908 (.A1(n_1_737_710), .A2(n_1_737_5190), .B1(n_1_737_2628), 
      .B2(n_1_737_2627), .ZN(n_1_737_2626));
   AND2_X1 i_1_737_2909 (.A1(n_1_737_710), .A2(n_1_737_5190), .ZN(n_1_737_2627));
   OAI21_X1 i_1_737_2910 (.A(\out_bs[3] [6]), .B1(\out_bs[3] [5]), .B2(
      n_1_737_4223), .ZN(n_1_737_2628));
   NOR2_X1 i_1_737_2911 (.A1(n_1_737_706), .A2(n_1_737_2629), .ZN(n_282));
   NAND2_X1 i_1_737_2912 (.A1(n_1_737_706), .A2(n_1_737_2629), .ZN(n_283));
   OAI21_X1 i_1_737_2913 (.A(n_1_737_2666), .B1(\out_bs[6] [5]), .B2(
      n_1_737_4514), .ZN(n_1_737_2629));
   NOR2_X1 i_1_737_2914 (.A1(n_1_737_705), .A2(n_1_737_2630), .ZN(n_284));
   NAND2_X1 i_1_737_2915 (.A1(n_1_737_705), .A2(n_1_737_2630), .ZN(n_285));
   OAI21_X1 i_1_737_2916 (.A(n_844), .B1(n_845), .B2(n_1_737_4255), .ZN(
      n_1_737_2630));
   OR4_X1 i_1_737_2917 (.A1(n_1_737_2632), .A2(n_1_737_2631), .A3(n_1_737_2635), 
      .A4(n_1_737_2644), .ZN(n_286));
   AOI21_X1 i_1_737_2918 (.A(n_1_737_700), .B1(n_1_737_5337), .B2(n_1_737_2636), 
      .ZN(n_1_737_2631));
   AOI21_X1 i_1_737_2919 (.A(n_1_737_2633), .B1(n_1_737_702), .B2(n_1_737_5236), 
      .ZN(n_1_737_2632));
   INV_X1 i_1_737_2920 (.A(n_1_737_2634), .ZN(n_1_737_2633));
   OAI22_X1 i_1_737_2921 (.A1(n_1_737_5651), .A2(n_1_737_4277), .B1(n_1_737_702), 
      .B2(n_1_737_5236), .ZN(n_1_737_2634));
   OAI211_X1 i_1_737_2922 (.A(n_1_737_2638), .B(n_1_737_2641), .C1(n_1_737_5337), 
      .C2(n_1_737_2636), .ZN(n_1_737_2635));
   OAI21_X1 i_1_737_2923 (.A(\out_bs[0] [6]), .B1(\out_bs[0] [5]), .B2(
      n_1_737_4266), .ZN(n_1_737_2636));
   INV_X1 i_1_737_2924 (.A(n_1_737_2638), .ZN(n_1_737_2637));
   OAI21_X1 i_1_737_2925 (.A(n_1_737_2639), .B1(n_1_737_5507), .B2(n_1_737_5297), 
      .ZN(n_1_737_2638));
   OAI22_X1 i_1_737_2926 (.A1(n_1_737_5664), .A2(n_1_737_4272), .B1(n_1_737_701), 
      .B2(n_1_737_5298), .ZN(n_1_737_2639));
   INV_X1 i_1_737_2927 (.A(n_1_737_2641), .ZN(n_1_737_2640));
   OAI21_X1 i_1_737_2928 (.A(n_1_737_2642), .B1(n_1_737_5506), .B2(n_1_737_5189), 
      .ZN(n_1_737_2641));
   OAI21_X1 i_1_737_2929 (.A(n_1_737_2643), .B1(n_1_737_703), .B2(n_1_737_5190), 
      .ZN(n_1_737_2642));
   OAI21_X1 i_1_737_2930 (.A(\out_bs[3] [6]), .B1(\out_bs[3] [5]), .B2(
      n_1_737_4263), .ZN(n_1_737_2643));
   AOI21_X1 i_1_737_2931 (.A(n_1_737_2645), .B1(n_1_737_704), .B2(n_1_737_5366), 
      .ZN(n_1_737_2644));
   INV_X1 i_1_737_2932 (.A(n_1_737_2646), .ZN(n_1_737_2645));
   OAI21_X1 i_1_737_2933 (.A(n_1_737_2647), .B1(n_1_737_704), .B2(n_1_737_5366), 
      .ZN(n_1_737_2646));
   OAI21_X1 i_1_737_2934 (.A(\out_bs[4] [6]), .B1(\out_bs[4] [5]), .B2(
      n_1_737_4285), .ZN(n_1_737_2647));
   NOR2_X1 i_1_737_2935 (.A1(n_1_737_698), .A2(n_1_737_2648), .ZN(n_287));
   NAND2_X1 i_1_737_2936 (.A1(n_1_737_698), .A2(n_1_737_2648), .ZN(n_288));
   AOI21_X1 i_1_737_2937 (.A(n_1_737_3110), .B1(n_1_737_4810), .B2(n_1_737_3108), 
      .ZN(n_1_737_2648));
   NAND4_X1 i_1_737_2938 (.A1(n_1_737_2655), .A2(n_1_737_2652), .A3(n_1_737_2649), 
      .A4(n_1_737_2663), .ZN(n_289));
   OAI21_X1 i_1_737_2939 (.A(n_1_737_2650), .B1(n_1_737_5509), .B2(n_1_737_5189), 
      .ZN(n_1_737_2649));
   OAI21_X1 i_1_737_2940 (.A(n_1_737_2651), .B1(n_1_737_696), .B2(n_1_737_5190), 
      .ZN(n_1_737_2650));
   OAI21_X1 i_1_737_2941 (.A(\out_bs[3] [6]), .B1(\out_bs[3] [5]), .B2(
      n_1_737_4308), .ZN(n_1_737_2651));
   OAI21_X1 i_1_737_2942 (.A(n_1_737_2653), .B1(n_1_737_5510), .B2(n_1_737_5235), 
      .ZN(n_1_737_2652));
   OAI21_X1 i_1_737_2943 (.A(n_1_737_2654), .B1(n_1_737_695), .B2(n_1_737_5236), 
      .ZN(n_1_737_2653));
   OAI21_X1 i_1_737_2944 (.A(\out_bs[2] [6]), .B1(\out_bs[2] [5]), .B2(
      n_1_737_4297), .ZN(n_1_737_2654));
   AOI211_X1 i_1_737_2945 (.A(n_1_737_2656), .B(n_1_737_2660), .C1(n_1_737_5336), 
      .C2(n_1_737_2661), .ZN(n_1_737_2655));
   AOI21_X1 i_1_737_2946 (.A(n_1_737_2657), .B1(n_1_737_694), .B2(n_1_737_5298), 
      .ZN(n_1_737_2656));
   INV_X1 i_1_737_2947 (.A(n_1_737_2658), .ZN(n_1_737_2657));
   OAI21_X1 i_1_737_2948 (.A(n_1_737_2659), .B1(n_1_737_694), .B2(n_1_737_5298), 
      .ZN(n_1_737_2658));
   OAI21_X1 i_1_737_2949 (.A(\out_bs[1] [6]), .B1(\out_bs[1] [5]), .B2(
      n_1_737_4303), .ZN(n_1_737_2659));
   AOI21_X1 i_1_737_2950 (.A(n_1_737_693), .B1(n_1_737_5337), .B2(n_1_737_2662), 
      .ZN(n_1_737_2660));
   INV_X1 i_1_737_2951 (.A(n_1_737_2662), .ZN(n_1_737_2661));
   OAI21_X1 i_1_737_2952 (.A(\out_bs[0] [6]), .B1(\out_bs[0] [5]), .B2(
      n_1_737_4292), .ZN(n_1_737_2662));
   OAI21_X1 i_1_737_2953 (.A(n_1_737_2664), .B1(n_1_737_5508), .B2(n_1_737_5365), 
      .ZN(n_1_737_2663));
   OAI21_X1 i_1_737_2954 (.A(n_1_737_2665), .B1(n_1_737_697), .B2(n_1_737_5366), 
      .ZN(n_1_737_2664));
   OAI21_X1 i_1_737_2955 (.A(\out_bs[4] [6]), .B1(\out_bs[4] [5]), .B2(
      n_1_737_4314), .ZN(n_1_737_2665));
   NOR2_X1 i_1_737_2956 (.A1(n_1_737_692), .A2(n_1_737_2667), .ZN(n_290));
   NAND2_X1 i_1_737_2957 (.A1(n_1_737_692), .A2(n_1_737_2667), .ZN(n_291));
   INV_X1 i_1_737_2958 (.A(n_1_737_2667), .ZN(n_1_737_2666));
   OAI21_X1 i_1_737_2959 (.A(\out_bs[6] [6]), .B1(\out_bs[6] [5]), .B2(
      n_1_737_3332), .ZN(n_1_737_2667));
   NOR2_X1 i_1_737_2960 (.A1(n_1_737_691), .A2(n_1_737_2728), .ZN(n_292));
   NAND2_X1 i_1_737_2961 (.A1(n_1_737_691), .A2(n_1_737_2728), .ZN(n_293));
   OAI211_X1 i_1_737_2962 (.A(n_1_737_2683), .B(n_1_737_2668), .C1(n_1_737_686), 
      .C2(n_1_737_2684), .ZN(n_294));
   NOR4_X1 i_1_737_2963 (.A1(n_1_737_2674), .A2(n_1_737_2669), .A3(n_1_737_2677), 
      .A4(n_1_737_2680), .ZN(n_1_737_2668));
   INV_X1 i_1_737_2964 (.A(n_1_737_2670), .ZN(n_1_737_2669));
   OAI21_X1 i_1_737_2965 (.A(n_1_737_2671), .B1(n_1_737_5297), .B2(n_1_737_2673), 
      .ZN(n_1_737_2670));
   OAI21_X1 i_1_737_2966 (.A(n_1_737_687), .B1(n_1_737_5298), .B2(n_1_737_2672), 
      .ZN(n_1_737_2671));
   INV_X1 i_1_737_2967 (.A(n_1_737_2673), .ZN(n_1_737_2672));
   NOR2_X1 i_1_737_2968 (.A1(n_1_737_5664), .A2(n_1_737_4449), .ZN(n_1_737_2673));
   AOI21_X1 i_1_737_2969 (.A(n_1_737_2675), .B1(n_1_737_689), .B2(n_1_737_5190), 
      .ZN(n_1_737_2674));
   INV_X1 i_1_737_2970 (.A(n_1_737_2676), .ZN(n_1_737_2675));
   OAI22_X1 i_1_737_2971 (.A1(n_1_737_5638), .A2(n_1_737_4425), .B1(n_1_737_689), 
      .B2(n_1_737_5190), .ZN(n_1_737_2676));
   INV_X1 i_1_737_2972 (.A(n_1_737_2678), .ZN(n_1_737_2677));
   OAI21_X1 i_1_737_2973 (.A(n_1_737_2679), .B1(n_1_737_5512), .B2(n_1_737_5235), 
      .ZN(n_1_737_2678));
   OAI22_X1 i_1_737_2974 (.A1(n_1_737_5651), .A2(n_1_737_4414), .B1(n_1_737_688), 
      .B2(n_1_737_5236), .ZN(n_1_737_2679));
   INV_X1 i_1_737_2975 (.A(n_1_737_2681), .ZN(n_1_737_2680));
   OAI21_X1 i_1_737_2976 (.A(n_1_737_2682), .B1(n_1_737_5511), .B2(n_1_737_5365), 
      .ZN(n_1_737_2681));
   OAI22_X1 i_1_737_2977 (.A1(n_1_737_5625), .A2(n_1_737_4461), .B1(n_1_737_690), 
      .B2(n_1_737_5366), .ZN(n_1_737_2682));
   OAI21_X1 i_1_737_2978 (.A(n_1_737_5336), .B1(n_1_737_5513), .B2(n_1_737_2685), 
      .ZN(n_1_737_2683));
   INV_X1 i_1_737_2979 (.A(n_1_737_2685), .ZN(n_1_737_2684));
   NOR2_X1 i_1_737_2980 (.A1(n_1_737_5671), .A2(n_1_737_4436), .ZN(n_1_737_2685));
   NOR2_X1 i_1_737_2981 (.A1(n_1_737_684), .A2(n_1_737_2686), .ZN(n_295));
   NAND2_X1 i_1_737_2982 (.A1(n_1_737_684), .A2(n_1_737_2686), .ZN(n_296));
   INV_X1 i_1_737_2983 (.A(n_1_737_2687), .ZN(n_1_737_2686));
   OAI21_X1 i_1_737_2984 (.A(n_1_737_2728), .B1(n_1_737_4882), .B2(n_1_737_3107), 
      .ZN(n_1_737_2687));
   NAND4_X1 i_1_737_2985 (.A1(n_1_737_2694), .A2(n_1_737_2688), .A3(n_1_737_2692), 
      .A4(n_1_737_2702), .ZN(n_297));
   AOI21_X1 i_1_737_2986 (.A(n_1_737_2698), .B1(n_1_737_2690), .B2(n_1_737_2689), 
      .ZN(n_1_737_2688));
   NAND2_X1 i_1_737_2987 (.A1(n_1_737_679), .A2(n_1_737_5337), .ZN(n_1_737_2689));
   OAI22_X1 i_1_737_2988 (.A1(n_1_737_4341), .A2(n_1_737_2713), .B1(n_1_737_679), 
      .B2(n_1_737_5337), .ZN(n_1_737_2690));
   INV_X1 i_1_737_2989 (.A(n_1_737_2692), .ZN(n_1_737_2691));
   OAI21_X1 i_1_737_2990 (.A(n_1_737_2693), .B1(n_1_737_5515), .B2(n_1_737_5189), 
      .ZN(n_1_737_2692));
   OAI22_X1 i_1_737_2991 (.A1(n_1_737_5638), .A2(n_1_737_4346), .B1(n_1_737_682), 
      .B2(n_1_737_5190), .ZN(n_1_737_2693));
   INV_X1 i_1_737_2992 (.A(n_1_737_2695), .ZN(n_1_737_2694));
   AOI21_X1 i_1_737_2993 (.A(n_1_737_2696), .B1(n_1_737_681), .B2(n_1_737_5236), 
      .ZN(n_1_737_2695));
   AOI21_X1 i_1_737_2994 (.A(n_1_737_2697), .B1(n_1_737_5516), .B2(n_1_737_5235), 
      .ZN(n_1_737_2696));
   AOI21_X1 i_1_737_2995 (.A(n_1_737_5651), .B1(n_1_737_5650), .B2(n_1_737_4360), 
      .ZN(n_1_737_2697));
   INV_X1 i_1_737_2996 (.A(n_1_737_2699), .ZN(n_1_737_2698));
   OAI21_X1 i_1_737_2997 (.A(n_1_737_2700), .B1(n_1_737_5517), .B2(n_1_737_5297), 
      .ZN(n_1_737_2699));
   OAI21_X1 i_1_737_2998 (.A(n_1_737_2701), .B1(n_1_737_680), .B2(n_1_737_5298), 
      .ZN(n_1_737_2700));
   OAI21_X1 i_1_737_2999 (.A(n_1_737_2718), .B1(\out_bs[1] [0]), .B2(
      n_1_737_4448), .ZN(n_1_737_2701));
   OAI21_X1 i_1_737_3000 (.A(n_1_737_2703), .B1(n_1_737_5514), .B2(n_1_737_5365), 
      .ZN(n_1_737_2702));
   OAI21_X1 i_1_737_3001 (.A(n_1_737_2704), .B1(n_1_737_683), .B2(n_1_737_5366), 
      .ZN(n_1_737_2703));
   OAI21_X1 i_1_737_3002 (.A(n_1_737_2725), .B1(\out_bs[4] [0]), .B2(
      n_1_737_4460), .ZN(n_1_737_2704));
   NOR2_X1 i_1_737_3003 (.A1(n_1_737_677), .A2(n_1_737_2705), .ZN(n_298));
   NAND2_X1 i_1_737_3004 (.A1(n_1_737_677), .A2(n_1_737_2705), .ZN(n_299));
   INV_X1 i_1_737_3005 (.A(n_1_737_2706), .ZN(n_1_737_2705));
   OAI21_X1 i_1_737_3006 (.A(n_1_737_2728), .B1(n_1_737_4925), .B2(n_1_737_3107), 
      .ZN(n_1_737_2706));
   NAND2_X1 i_1_737_3007 (.A1(n_1_737_2722), .A2(n_1_737_2707), .ZN(n_300));
   NOR4_X1 i_1_737_3008 (.A1(n_1_737_2719), .A2(n_1_737_2712), .A3(n_1_737_2709), 
      .A4(n_1_737_2708), .ZN(n_1_737_2707));
   AOI21_X1 i_1_737_3009 (.A(n_1_737_672), .B1(n_1_737_5337), .B2(n_1_737_2713), 
      .ZN(n_1_737_2708));
   AOI21_X1 i_1_737_3010 (.A(n_1_737_2710), .B1(n_1_737_674), .B2(n_1_737_5236), 
      .ZN(n_1_737_2709));
   INV_X1 i_1_737_3011 (.A(n_1_737_2711), .ZN(n_1_737_2710));
   OAI22_X1 i_1_737_3012 (.A1(n_1_737_5651), .A2(n_1_737_4386), .B1(n_1_737_674), 
      .B2(n_1_737_5236), .ZN(n_1_737_2711));
   OAI21_X1 i_1_737_3013 (.A(n_1_737_2715), .B1(n_1_737_5337), .B2(n_1_737_2713), 
      .ZN(n_1_737_2712));
   OAI21_X1 i_1_737_3014 (.A(\out_bs[0] [6]), .B1(n_1_737_4435), .B2(
      n_1_737_4392), .ZN(n_1_737_2713));
   INV_X1 i_1_737_3015 (.A(n_1_737_2715), .ZN(n_1_737_2714));
   OAI21_X1 i_1_737_3016 (.A(n_1_737_2716), .B1(n_1_737_5297), .B2(n_1_737_2718), 
      .ZN(n_1_737_2715));
   OAI21_X1 i_1_737_3017 (.A(n_1_737_673), .B1(n_1_737_5298), .B2(n_1_737_2717), 
      .ZN(n_1_737_2716));
   INV_X1 i_1_737_3018 (.A(n_1_737_2718), .ZN(n_1_737_2717));
   NOR2_X1 i_1_737_3019 (.A1(n_1_737_5664), .A2(n_1_737_4375), .ZN(n_1_737_2718));
   AOI21_X1 i_1_737_3020 (.A(n_1_737_2720), .B1(n_1_737_675), .B2(n_1_737_5190), 
      .ZN(n_1_737_2719));
   INV_X1 i_1_737_3021 (.A(n_1_737_2721), .ZN(n_1_737_2720));
   OAI22_X1 i_1_737_3022 (.A1(n_1_737_5638), .A2(n_1_737_4380), .B1(n_1_737_675), 
      .B2(n_1_737_5190), .ZN(n_1_737_2721));
   OAI21_X1 i_1_737_3023 (.A(n_1_737_2723), .B1(n_1_737_5365), .B2(n_1_737_2725), 
      .ZN(n_1_737_2722));
   OAI21_X1 i_1_737_3024 (.A(n_1_737_676), .B1(n_1_737_5366), .B2(n_1_737_2724), 
      .ZN(n_1_737_2723));
   INV_X1 i_1_737_3025 (.A(n_1_737_2725), .ZN(n_1_737_2724));
   NOR2_X1 i_1_737_3026 (.A1(n_1_737_5625), .A2(n_1_737_4397), .ZN(n_1_737_2725));
   NOR2_X1 i_1_737_3027 (.A1(n_1_737_670), .A2(n_1_737_2726), .ZN(n_301));
   NAND2_X1 i_1_737_3028 (.A1(n_1_737_670), .A2(n_1_737_2726), .ZN(n_302));
   INV_X1 i_1_737_3029 (.A(n_1_737_2727), .ZN(n_1_737_2726));
   OAI21_X1 i_1_737_3030 (.A(n_1_737_2728), .B1(n_1_737_4964), .B2(n_1_737_3107), 
      .ZN(n_1_737_2727));
   OAI21_X1 i_1_737_3031 (.A(n_844), .B1(n_845), .B2(n_1_737_4404), .ZN(
      n_1_737_2728));
   OR4_X1 i_1_737_3032 (.A1(n_1_737_2730), .A2(n_1_737_2729), .A3(n_1_737_2733), 
      .A4(n_1_737_2741), .ZN(n_303));
   AOI21_X1 i_1_737_3033 (.A(n_1_737_665), .B1(n_1_737_5337), .B2(n_1_737_2734), 
      .ZN(n_1_737_2729));
   INV_X1 i_1_737_3034 (.A(n_1_737_2731), .ZN(n_1_737_2730));
   OAI21_X1 i_1_737_3035 (.A(n_1_737_2732), .B1(n_1_737_5519), .B2(n_1_737_5189), 
      .ZN(n_1_737_2731));
   OAI22_X1 i_1_737_3036 (.A1(n_1_737_5638), .A2(n_1_737_4423), .B1(n_1_737_668), 
      .B2(n_1_737_5190), .ZN(n_1_737_2732));
   OAI211_X1 i_1_737_3037 (.A(n_1_737_2736), .B(n_1_737_2739), .C1(n_1_737_5337), 
      .C2(n_1_737_2734), .ZN(n_1_737_2733));
   OAI21_X1 i_1_737_3038 (.A(\out_bs[0] [6]), .B1(n_1_737_4439), .B2(
      n_1_737_4435), .ZN(n_1_737_2734));
   INV_X1 i_1_737_3039 (.A(n_1_737_2736), .ZN(n_1_737_2735));
   OAI21_X1 i_1_737_3040 (.A(n_1_737_2737), .B1(n_1_737_5521), .B2(n_1_737_5297), 
      .ZN(n_1_737_2736));
   OAI22_X1 i_1_737_3041 (.A1(n_1_737_5664), .A2(n_1_737_4447), .B1(n_1_737_666), 
      .B2(n_1_737_5298), .ZN(n_1_737_2737));
   INV_X1 i_1_737_3042 (.A(n_1_737_2739), .ZN(n_1_737_2738));
   OAI21_X1 i_1_737_3043 (.A(n_1_737_2740), .B1(n_1_737_5520), .B2(n_1_737_5235), 
      .ZN(n_1_737_2739));
   OAI22_X1 i_1_737_3044 (.A1(n_1_737_5651), .A2(n_1_737_4411), .B1(n_1_737_667), 
      .B2(n_1_737_5236), .ZN(n_1_737_2740));
   AOI21_X1 i_1_737_3045 (.A(n_1_737_2742), .B1(n_1_737_669), .B2(n_1_737_5366), 
      .ZN(n_1_737_2741));
   AOI22_X1 i_1_737_3046 (.A1(\out_bs[4] [6]), .A2(n_1_737_4459), .B1(
      n_1_737_5518), .B2(n_1_737_5365), .ZN(n_1_737_2742));
   NOR2_X1 i_1_737_3047 (.A1(n_1_737_664), .A2(n_1_737_2743), .ZN(n_304));
   NAND2_X1 i_1_737_3048 (.A1(n_1_737_664), .A2(n_1_737_2743), .ZN(n_305));
   INV_X1 i_1_737_3049 (.A(n_1_737_2744), .ZN(n_1_737_2743));
   AOI21_X1 i_1_737_3050 (.A(n_1_737_3082), .B1(n_1_737_5606), .B2(n_1_737_4513), 
      .ZN(n_1_737_2744));
   NOR2_X1 i_1_737_3051 (.A1(n_1_737_663), .A2(n_1_737_2780), .ZN(n_306));
   NAND2_X1 i_1_737_3052 (.A1(n_1_737_663), .A2(n_1_737_2780), .ZN(n_307));
   NAND4_X1 i_1_737_3053 (.A1(n_1_737_2749), .A2(n_1_737_2745), .A3(n_1_737_2747), 
      .A4(n_1_737_2756), .ZN(n_308));
   OAI21_X1 i_1_737_3054 (.A(n_1_737_2746), .B1(n_1_737_5524), .B2(n_1_737_5235), 
      .ZN(n_1_737_2745));
   OAI22_X1 i_1_737_3055 (.A1(n_1_737_5651), .A2(n_1_737_4553), .B1(n_1_737_660), 
      .B2(n_1_737_5236), .ZN(n_1_737_2746));
   OAI21_X1 i_1_737_3056 (.A(n_1_737_2748), .B1(n_1_737_5523), .B2(n_1_737_5189), 
      .ZN(n_1_737_2747));
   OAI21_X1 i_1_737_3057 (.A(n_1_737_2793), .B1(n_1_737_661), .B2(n_1_737_5190), 
      .ZN(n_1_737_2748));
   AOI21_X1 i_1_737_3058 (.A(n_1_737_2750), .B1(n_1_737_5336), .B2(n_1_737_2754), 
      .ZN(n_1_737_2749));
   OAI21_X1 i_1_737_3059 (.A(n_1_737_2752), .B1(n_1_737_658), .B2(n_1_737_2755), 
      .ZN(n_1_737_2750));
   INV_X1 i_1_737_3060 (.A(n_1_737_2752), .ZN(n_1_737_2751));
   OAI21_X1 i_1_737_3061 (.A(n_1_737_2753), .B1(n_1_737_5525), .B2(n_1_737_5297), 
      .ZN(n_1_737_2752));
   OAI221_X1 i_1_737_3062 (.A(n_1_737_3015), .B1(n_1_737_5664), .B2(n_1_737_4528), 
      .C1(n_1_737_659), .C2(n_1_737_5298), .ZN(n_1_737_2753));
   NAND2_X1 i_1_737_3063 (.A1(n_1_737_658), .A2(n_1_737_2755), .ZN(n_1_737_2754));
   OAI21_X1 i_1_737_3064 (.A(\out_bs[0] [6]), .B1(\out_bs[0] [5]), .B2(
      n_1_737_4544), .ZN(n_1_737_2755));
   OAI21_X1 i_1_737_3065 (.A(n_1_737_2757), .B1(n_1_737_5522), .B2(n_1_737_5365), 
      .ZN(n_1_737_2756));
   OAI22_X1 i_1_737_3066 (.A1(n_1_737_5625), .A2(n_1_737_4563), .B1(n_1_737_662), 
      .B2(n_1_737_5366), .ZN(n_1_737_2757));
   NOR2_X1 i_1_737_3067 (.A1(n_1_737_656), .A2(n_1_737_2758), .ZN(n_309));
   NAND2_X1 i_1_737_3068 (.A1(n_1_737_656), .A2(n_1_737_2758), .ZN(n_310));
   AOI21_X1 i_1_737_3069 (.A(n_1_737_3110), .B1(n_1_737_5020), .B2(n_1_737_3108), 
      .ZN(n_1_737_2758));
   NAND3_X1 i_1_737_3070 (.A1(n_1_737_2761), .A2(n_1_737_2759), .A3(n_1_737_2775), 
      .ZN(n_311));
   NOR3_X1 i_1_737_3071 (.A1(n_1_737_2773), .A2(n_1_737_2768), .A3(n_1_737_2764), 
      .ZN(n_1_737_2759));
   INV_X1 i_1_737_3072 (.A(n_1_737_2761), .ZN(n_1_737_2760));
   OAI21_X1 i_1_737_3073 (.A(n_1_737_2762), .B1(n_1_737_5527), .B2(n_1_737_5189), 
      .ZN(n_1_737_2761));
   OAI21_X1 i_1_737_3074 (.A(n_1_737_2763), .B1(n_1_737_654), .B2(n_1_737_5190), 
      .ZN(n_1_737_2762));
   OAI21_X1 i_1_737_3075 (.A(\out_bs[3] [6]), .B1(\out_bs[3] [5]), .B2(
      n_1_737_4491), .ZN(n_1_737_2763));
   AOI21_X1 i_1_737_3076 (.A(n_1_737_2765), .B1(n_1_737_653), .B2(n_1_737_5236), 
      .ZN(n_1_737_2764));
   INV_X1 i_1_737_3077 (.A(n_1_737_2766), .ZN(n_1_737_2765));
   OAI21_X1 i_1_737_3078 (.A(n_1_737_2767), .B1(n_1_737_653), .B2(n_1_737_5236), 
      .ZN(n_1_737_2766));
   OAI21_X1 i_1_737_3079 (.A(\out_bs[2] [6]), .B1(\out_bs[2] [5]), .B2(
      n_1_737_4504), .ZN(n_1_737_2767));
   OAI21_X1 i_1_737_3080 (.A(n_1_737_2770), .B1(n_1_737_5337), .B2(n_1_737_2774), 
      .ZN(n_1_737_2768));
   INV_X1 i_1_737_3081 (.A(n_1_737_2770), .ZN(n_1_737_2769));
   OAI21_X1 i_1_737_3082 (.A(n_1_737_2771), .B1(n_1_737_5528), .B2(n_1_737_5297), 
      .ZN(n_1_737_2770));
   OAI21_X1 i_1_737_3083 (.A(n_1_737_2772), .B1(n_1_737_652), .B2(n_1_737_5298), 
      .ZN(n_1_737_2771));
   OAI21_X1 i_1_737_3084 (.A(\out_bs[1] [6]), .B1(\out_bs[1] [5]), .B2(
      n_1_737_4498), .ZN(n_1_737_2772));
   AOI21_X1 i_1_737_3085 (.A(n_1_737_651), .B1(n_1_737_5337), .B2(n_1_737_2774), 
      .ZN(n_1_737_2773));
   OAI21_X1 i_1_737_3086 (.A(\out_bs[0] [6]), .B1(\out_bs[0] [5]), .B2(
      n_1_737_4486), .ZN(n_1_737_2774));
   OAI21_X1 i_1_737_3087 (.A(n_1_737_2776), .B1(n_1_737_5526), .B2(n_1_737_5365), 
      .ZN(n_1_737_2775));
   OAI21_X1 i_1_737_3088 (.A(n_1_737_2777), .B1(n_1_737_655), .B2(n_1_737_5366), 
      .ZN(n_1_737_2776));
   OAI21_X1 i_1_737_3089 (.A(\out_bs[4] [6]), .B1(\out_bs[4] [5]), .B2(
      n_1_737_4510), .ZN(n_1_737_2777));
   NOR2_X1 i_1_737_3090 (.A1(n_1_737_650), .A2(n_1_737_2778), .ZN(n_312));
   NAND2_X1 i_1_737_3091 (.A1(n_1_737_650), .A2(n_1_737_2778), .ZN(n_313));
   OAI21_X1 i_1_737_3092 (.A(\out_bs[6] [6]), .B1(\out_bs[6] [5]), .B2(
      n_1_737_4512), .ZN(n_1_737_2778));
   NOR2_X1 i_1_737_3093 (.A1(n_1_737_649), .A2(n_1_737_2779), .ZN(n_314));
   NAND2_X1 i_1_737_3094 (.A1(n_1_737_649), .A2(n_1_737_2779), .ZN(n_315));
   OAI21_X1 i_1_737_3095 (.A(n_844), .B1(n_845), .B2(n_1_737_4516), .ZN(
      n_1_737_2779));
   OAI21_X1 i_1_737_3096 (.A(n_844), .B1(n_845), .B2(n_1_737_4519), .ZN(
      n_1_737_2780));
   NAND3_X1 i_1_737_3097 (.A1(n_1_737_2789), .A2(n_1_737_2786), .A3(n_1_737_2781), 
      .ZN(n_316));
   AOI211_X1 i_1_737_3098 (.A(n_1_737_2794), .B(n_1_737_2784), .C1(n_1_737_2783), 
      .C2(n_1_737_2782), .ZN(n_1_737_2781));
   NAND2_X1 i_1_737_3099 (.A1(n_1_737_644), .A2(n_1_737_5337), .ZN(n_1_737_2782));
   OAI22_X1 i_1_737_3100 (.A1(n_1_737_5671), .A2(n_1_737_4541), .B1(n_1_737_644), 
      .B2(n_1_737_5337), .ZN(n_1_737_2783));
   AOI21_X1 i_1_737_3101 (.A(n_1_737_2785), .B1(n_1_737_646), .B2(n_1_737_5236), 
      .ZN(n_1_737_2784));
   AOI22_X1 i_1_737_3102 (.A1(\out_bs[2] [6]), .A2(n_1_737_4550), .B1(
      n_1_737_5529), .B2(n_1_737_5235), .ZN(n_1_737_2785));
   INV_X1 i_1_737_3103 (.A(n_1_737_2787), .ZN(n_1_737_2786));
   AOI21_X1 i_1_737_3104 (.A(n_1_737_2788), .B1(n_1_737_645), .B2(n_1_737_5298), 
      .ZN(n_1_737_2787));
   AOI22_X1 i_1_737_3105 (.A1(\out_bs[1] [6]), .A2(n_1_737_4526), .B1(
      n_1_737_5530), .B2(n_1_737_5297), .ZN(n_1_737_2788));
   INV_X1 i_1_737_3106 (.A(n_1_737_2790), .ZN(n_1_737_2789));
   OAI21_X1 i_1_737_3107 (.A(n_1_737_2791), .B1(n_1_737_647), .B2(n_1_737_5190), 
      .ZN(n_1_737_2790));
   INV_X1 i_1_737_3108 (.A(n_1_737_2792), .ZN(n_1_737_2791));
   AOI221_X1 i_1_737_3109 (.A(n_1_737_5638), .B1(n_1_737_5637), .B2(n_1_737_4532), 
      .C1(n_1_737_647), .C2(n_1_737_5190), .ZN(n_1_737_2792));
   OAI21_X1 i_1_737_3110 (.A(\out_bs[3] [6]), .B1(\out_bs[3] [5]), .B2(
      n_1_737_4535), .ZN(n_1_737_2793));
   OAI22_X1 i_1_737_3111 (.A1(n_1_737_648), .A2(n_1_737_5366), .B1(n_1_737_2796), 
      .B2(n_1_737_2795), .ZN(n_1_737_2794));
   OAI21_X1 i_1_737_3112 (.A(\out_bs[4] [6]), .B1(\out_bs[4] [5]), .B2(
      n_1_737_4560), .ZN(n_1_737_2795));
   AND2_X1 i_1_737_3113 (.A1(n_1_737_648), .A2(n_1_737_5366), .ZN(n_1_737_2796));
   NOR2_X1 i_1_737_3114 (.A1(n_1_737_642), .A2(n_1_737_2797), .ZN(n_317));
   NAND2_X1 i_1_737_3115 (.A1(n_1_737_642), .A2(n_1_737_2797), .ZN(n_318));
   AOI21_X1 i_1_737_3116 (.A(n_1_737_3110), .B1(n_1_737_5172), .B2(n_1_737_3108), 
      .ZN(n_1_737_2797));
   NAND3_X1 i_1_737_3117 (.A1(n_1_737_2800), .A2(n_1_737_2798), .A3(n_1_737_2814), 
      .ZN(n_319));
   NOR3_X1 i_1_737_3118 (.A1(n_1_737_2812), .A2(n_1_737_2807), .A3(n_1_737_2803), 
      .ZN(n_1_737_2798));
   INV_X1 i_1_737_3119 (.A(n_1_737_2800), .ZN(n_1_737_2799));
   OAI21_X1 i_1_737_3120 (.A(n_1_737_2801), .B1(n_1_737_5532), .B2(n_1_737_5189), 
      .ZN(n_1_737_2800));
   OAI21_X1 i_1_737_3121 (.A(n_1_737_2802), .B1(n_1_737_640), .B2(n_1_737_5190), 
      .ZN(n_1_737_2801));
   OAI21_X1 i_1_737_3122 (.A(\out_bs[3] [6]), .B1(\out_bs[3] [5]), .B2(
      n_1_737_4576), .ZN(n_1_737_2802));
   AOI21_X1 i_1_737_3123 (.A(n_1_737_2804), .B1(n_1_737_639), .B2(n_1_737_5236), 
      .ZN(n_1_737_2803));
   INV_X1 i_1_737_3124 (.A(n_1_737_2805), .ZN(n_1_737_2804));
   OAI21_X1 i_1_737_3125 (.A(n_1_737_2806), .B1(n_1_737_639), .B2(n_1_737_5236), 
      .ZN(n_1_737_2805));
   OAI21_X1 i_1_737_3126 (.A(\out_bs[2] [6]), .B1(\out_bs[2] [5]), .B2(
      n_1_737_4588), .ZN(n_1_737_2806));
   OAI21_X1 i_1_737_3127 (.A(n_1_737_2809), .B1(n_1_737_5337), .B2(n_1_737_2813), 
      .ZN(n_1_737_2807));
   INV_X1 i_1_737_3128 (.A(n_1_737_2809), .ZN(n_1_737_2808));
   OAI21_X1 i_1_737_3129 (.A(n_1_737_2810), .B1(n_1_737_5533), .B2(n_1_737_5297), 
      .ZN(n_1_737_2809));
   OAI21_X1 i_1_737_3130 (.A(n_1_737_2811), .B1(n_1_737_638), .B2(n_1_737_5298), 
      .ZN(n_1_737_2810));
   OAI21_X1 i_1_737_3131 (.A(\out_bs[1] [6]), .B1(\out_bs[1] [5]), .B2(
      n_1_737_4583), .ZN(n_1_737_2811));
   AOI21_X1 i_1_737_3132 (.A(n_1_737_637), .B1(n_1_737_5337), .B2(n_1_737_2813), 
      .ZN(n_1_737_2812));
   OAI21_X1 i_1_737_3133 (.A(\out_bs[0] [6]), .B1(\out_bs[0] [5]), .B2(
      n_1_737_4571), .ZN(n_1_737_2813));
   OAI21_X1 i_1_737_3134 (.A(n_1_737_2815), .B1(n_1_737_5531), .B2(n_1_737_5365), 
      .ZN(n_1_737_2814));
   OAI21_X1 i_1_737_3135 (.A(n_1_737_2816), .B1(n_1_737_641), .B2(n_1_737_5366), 
      .ZN(n_1_737_2815));
   OAI21_X1 i_1_737_3136 (.A(\out_bs[4] [6]), .B1(\out_bs[4] [5]), .B2(
      n_1_737_4594), .ZN(n_1_737_2816));
   NOR2_X1 i_1_737_3137 (.A1(n_1_737_636), .A2(n_1_737_3082), .ZN(n_320));
   NAND2_X1 i_1_737_3138 (.A1(n_1_737_636), .A2(n_1_737_3082), .ZN(n_321));
   NOR2_X1 i_1_737_3139 (.A1(n_1_737_635), .A2(n_1_737_3106), .ZN(n_322));
   NAND2_X1 i_1_737_3140 (.A1(n_1_737_635), .A2(n_1_737_3106), .ZN(n_323));
   OAI211_X1 i_1_737_3141 (.A(n_1_737_2830), .B(n_1_737_2817), .C1(n_1_737_630), 
      .C2(n_1_737_2832), .ZN(n_324));
   NOR4_X1 i_1_737_3142 (.A1(n_1_737_2821), .A2(n_1_737_2818), .A3(n_1_737_2824), 
      .A4(n_1_737_2827), .ZN(n_1_737_2817));
   INV_X1 i_1_737_3143 (.A(n_1_737_2819), .ZN(n_1_737_2818));
   OAI21_X1 i_1_737_3144 (.A(n_1_737_2820), .B1(n_1_737_5535), .B2(n_1_737_5297), 
      .ZN(n_1_737_2819));
   OAI22_X1 i_1_737_3145 (.A1(n_1_737_5664), .A2(n_1_737_5293), .B1(n_1_737_631), 
      .B2(n_1_737_5298), .ZN(n_1_737_2820));
   AOI21_X1 i_1_737_3146 (.A(n_1_737_2822), .B1(n_1_737_633), .B2(n_1_737_5190), 
      .ZN(n_1_737_2821));
   INV_X1 i_1_737_3147 (.A(n_1_737_2823), .ZN(n_1_737_2822));
   OAI22_X1 i_1_737_3148 (.A1(n_1_737_5638), .A2(n_1_737_5229), .B1(n_1_737_633), 
      .B2(n_1_737_5190), .ZN(n_1_737_2823));
   AOI21_X1 i_1_737_3149 (.A(n_1_737_2825), .B1(n_1_737_632), .B2(n_1_737_5236), 
      .ZN(n_1_737_2824));
   INV_X1 i_1_737_3150 (.A(n_1_737_2826), .ZN(n_1_737_2825));
   OAI22_X1 i_1_737_3151 (.A1(n_1_737_5651), .A2(n_1_737_5260), .B1(n_1_737_632), 
      .B2(n_1_737_5236), .ZN(n_1_737_2826));
   INV_X1 i_1_737_3152 (.A(n_1_737_2828), .ZN(n_1_737_2827));
   OAI21_X1 i_1_737_3153 (.A(n_1_737_2829), .B1(n_1_737_5534), .B2(n_1_737_5365), 
      .ZN(n_1_737_2828));
   OAI22_X1 i_1_737_3154 (.A1(n_1_737_5625), .A2(n_1_737_5401), .B1(n_1_737_634), 
      .B2(n_1_737_5366), .ZN(n_1_737_2829));
   INV_X1 i_1_737_3155 (.A(n_1_737_2831), .ZN(n_1_737_2830));
   AOI21_X1 i_1_737_3156 (.A(n_1_737_5337), .B1(n_1_737_630), .B2(n_1_737_2832), 
      .ZN(n_1_737_2831));
   NAND2_X1 i_1_737_3157 (.A1(\out_bs[0] [6]), .A2(n_1_737_5331), .ZN(
      n_1_737_2832));
   NOR2_X1 i_1_737_3158 (.A1(n_1_737_628), .A2(n_1_737_2833), .ZN(n_325));
   NAND2_X1 i_1_737_3159 (.A1(n_1_737_628), .A2(n_1_737_2833), .ZN(n_326));
   AOI211_X1 i_1_737_3160 (.A(n_1_737_3110), .B(n_1_737_3108), .C1(n_844), 
      .C2(n_1_737_4615), .ZN(n_1_737_2833));
   OR4_X1 i_1_737_3161 (.A1(n_1_737_2835), .A2(n_1_737_2834), .A3(n_1_737_2839), 
      .A4(n_1_737_2848), .ZN(n_327));
   AOI21_X1 i_1_737_3162 (.A(n_1_737_623), .B1(n_1_737_5337), .B2(n_1_737_2840), 
      .ZN(n_1_737_2834));
   INV_X1 i_1_737_3163 (.A(n_1_737_2836), .ZN(n_1_737_2835));
   OAI21_X1 i_1_737_3164 (.A(n_1_737_2837), .B1(n_1_737_5538), .B2(n_1_737_5235), 
      .ZN(n_1_737_2836));
   OAI21_X1 i_1_737_3165 (.A(n_1_737_2838), .B1(n_1_737_625), .B2(n_1_737_5236), 
      .ZN(n_1_737_2837));
   OAI21_X1 i_1_737_3166 (.A(\out_bs[2] [6]), .B1(n_1_737_5259), .B2(
      n_1_737_4637), .ZN(n_1_737_2838));
   OAI211_X1 i_1_737_3167 (.A(n_1_737_2842), .B(n_1_737_2845), .C1(n_1_737_5337), 
      .C2(n_1_737_2840), .ZN(n_1_737_2839));
   OAI21_X1 i_1_737_3168 (.A(\out_bs[0] [6]), .B1(n_1_737_5331), .B2(
      n_1_737_4625), .ZN(n_1_737_2840));
   INV_X1 i_1_737_3169 (.A(n_1_737_2842), .ZN(n_1_737_2841));
   OAI21_X1 i_1_737_3170 (.A(n_1_737_2843), .B1(n_1_737_5539), .B2(n_1_737_5297), 
      .ZN(n_1_737_2842));
   OAI21_X1 i_1_737_3171 (.A(n_1_737_2844), .B1(n_1_737_624), .B2(n_1_737_5298), 
      .ZN(n_1_737_2843));
   OAI21_X1 i_1_737_3172 (.A(\out_bs[1] [6]), .B1(n_1_737_5292), .B2(
      n_1_737_4632), .ZN(n_1_737_2844));
   OAI21_X1 i_1_737_3173 (.A(n_1_737_2846), .B1(n_1_737_5537), .B2(n_1_737_5189), 
      .ZN(n_1_737_2845));
   OAI21_X1 i_1_737_3174 (.A(n_1_737_2847), .B1(n_1_737_626), .B2(n_1_737_5190), 
      .ZN(n_1_737_2846));
   OAI21_X1 i_1_737_3175 (.A(\out_bs[3] [6]), .B1(n_1_737_5228), .B2(
      n_1_737_4623), .ZN(n_1_737_2847));
   INV_X1 i_1_737_3176 (.A(n_1_737_2849), .ZN(n_1_737_2848));
   OAI21_X1 i_1_737_3177 (.A(n_1_737_2850), .B1(n_1_737_5536), .B2(n_1_737_5365), 
      .ZN(n_1_737_2849));
   OAI21_X1 i_1_737_3178 (.A(n_1_737_2851), .B1(n_1_737_627), .B2(n_1_737_5366), 
      .ZN(n_1_737_2850));
   OAI21_X1 i_1_737_3179 (.A(\out_bs[4] [6]), .B1(n_1_737_5400), .B2(
      n_1_737_4644), .ZN(n_1_737_2851));
   NOR2_X1 i_1_737_3180 (.A1(n_1_737_621), .A2(n_1_737_2852), .ZN(n_328));
   NAND2_X1 i_1_737_3181 (.A1(n_1_737_621), .A2(n_1_737_2852), .ZN(n_329));
   AOI211_X1 i_1_737_3182 (.A(n_1_737_3110), .B(n_1_737_3108), .C1(n_844), 
      .C2(n_1_737_4646), .ZN(n_1_737_2852));
   NAND4_X1 i_1_737_3183 (.A1(n_1_737_2856), .A2(n_1_737_2853), .A3(n_1_737_2864), 
      .A4(n_1_737_2867), .ZN(n_330));
   AOI21_X1 i_1_737_3184 (.A(n_1_737_2860), .B1(n_1_737_2855), .B2(n_1_737_2854), 
      .ZN(n_1_737_2853));
   NAND2_X1 i_1_737_3185 (.A1(n_1_737_616), .A2(n_1_737_5337), .ZN(n_1_737_2854));
   OAI21_X1 i_1_737_3186 (.A(n_1_737_2859), .B1(n_1_737_616), .B2(n_1_737_5337), 
      .ZN(n_1_737_2855));
   OAI21_X1 i_1_737_3187 (.A(n_1_737_2857), .B1(n_1_737_5542), .B2(n_1_737_5235), 
      .ZN(n_1_737_2856));
   OAI21_X1 i_1_737_3188 (.A(n_1_737_2858), .B1(n_1_737_618), .B2(n_1_737_5236), 
      .ZN(n_1_737_2857));
   OAI21_X1 i_1_737_3189 (.A(\out_bs[2] [6]), .B1(n_1_737_5259), .B2(
      n_1_737_4665), .ZN(n_1_737_2858));
   OAI21_X1 i_1_737_3190 (.A(\out_bs[0] [6]), .B1(n_1_737_5331), .B2(
      n_1_737_4670), .ZN(n_1_737_2859));
   INV_X1 i_1_737_3191 (.A(n_1_737_2861), .ZN(n_1_737_2860));
   OAI21_X1 i_1_737_3192 (.A(n_1_737_2862), .B1(n_1_737_5543), .B2(n_1_737_5297), 
      .ZN(n_1_737_2861));
   OAI21_X1 i_1_737_3193 (.A(n_1_737_2863), .B1(n_1_737_617), .B2(n_1_737_5298), 
      .ZN(n_1_737_2862));
   OAI21_X1 i_1_737_3194 (.A(\out_bs[1] [6]), .B1(n_1_737_5292), .B2(
      n_1_737_4652), .ZN(n_1_737_2863));
   OAI21_X1 i_1_737_3195 (.A(n_1_737_2865), .B1(n_1_737_5541), .B2(n_1_737_5189), 
      .ZN(n_1_737_2864));
   OAI21_X1 i_1_737_3196 (.A(n_1_737_2866), .B1(n_1_737_619), .B2(n_1_737_5190), 
      .ZN(n_1_737_2865));
   OAI21_X1 i_1_737_3197 (.A(\out_bs[3] [6]), .B1(n_1_737_5228), .B2(
      n_1_737_4659), .ZN(n_1_737_2866));
   OAI21_X1 i_1_737_3198 (.A(n_1_737_2868), .B1(n_1_737_5540), .B2(n_1_737_5365), 
      .ZN(n_1_737_2867));
   OAI21_X1 i_1_737_3199 (.A(n_1_737_2869), .B1(n_1_737_620), .B2(n_1_737_5366), 
      .ZN(n_1_737_2868));
   OAI21_X1 i_1_737_3200 (.A(\out_bs[4] [6]), .B1(n_1_737_5400), .B2(
      n_1_737_4677), .ZN(n_1_737_2869));
   NOR2_X1 i_1_737_3201 (.A1(n_1_737_614), .A2(n_1_737_2870), .ZN(n_331));
   NAND2_X1 i_1_737_3202 (.A1(n_1_737_614), .A2(n_1_737_2870), .ZN(n_332));
   AOI211_X1 i_1_737_3203 (.A(n_1_737_3110), .B(n_1_737_3108), .C1(n_844), 
      .C2(n_1_737_4679), .ZN(n_1_737_2870));
   NAND3_X1 i_1_737_3204 (.A1(n_1_737_2873), .A2(n_1_737_2871), .A3(n_1_737_2887), 
      .ZN(n_333));
   NOR3_X1 i_1_737_3205 (.A1(n_1_737_2885), .A2(n_1_737_2880), .A3(n_1_737_2876), 
      .ZN(n_1_737_2871));
   INV_X1 i_1_737_3206 (.A(n_1_737_2873), .ZN(n_1_737_2872));
   OAI21_X1 i_1_737_3207 (.A(n_1_737_2874), .B1(n_1_737_5545), .B2(n_1_737_5189), 
      .ZN(n_1_737_2873));
   OAI21_X1 i_1_737_3208 (.A(n_1_737_2875), .B1(n_1_737_612), .B2(n_1_737_5190), 
      .ZN(n_1_737_2874));
   OAI21_X1 i_1_737_3209 (.A(\out_bs[3] [6]), .B1(n_1_737_5228), .B2(
      n_1_737_4692), .ZN(n_1_737_2875));
   AOI21_X1 i_1_737_3210 (.A(n_1_737_2877), .B1(n_1_737_611), .B2(n_1_737_5236), 
      .ZN(n_1_737_2876));
   INV_X1 i_1_737_3211 (.A(n_1_737_2878), .ZN(n_1_737_2877));
   OAI21_X1 i_1_737_3212 (.A(n_1_737_2879), .B1(n_1_737_611), .B2(n_1_737_5236), 
      .ZN(n_1_737_2878));
   OAI21_X1 i_1_737_3213 (.A(\out_bs[2] [6]), .B1(n_1_737_5259), .B2(
      n_1_737_4707), .ZN(n_1_737_2879));
   OAI21_X1 i_1_737_3214 (.A(n_1_737_2882), .B1(n_1_737_5337), .B2(n_1_737_2886), 
      .ZN(n_1_737_2880));
   INV_X1 i_1_737_3215 (.A(n_1_737_2882), .ZN(n_1_737_2881));
   OAI21_X1 i_1_737_3216 (.A(n_1_737_2883), .B1(n_1_737_5546), .B2(n_1_737_5297), 
      .ZN(n_1_737_2882));
   OAI21_X1 i_1_737_3217 (.A(n_1_737_2884), .B1(n_1_737_610), .B2(n_1_737_5298), 
      .ZN(n_1_737_2883));
   OAI21_X1 i_1_737_3218 (.A(\out_bs[1] [6]), .B1(n_1_737_5292), .B2(
      n_1_737_4699), .ZN(n_1_737_2884));
   AOI21_X1 i_1_737_3219 (.A(n_1_737_609), .B1(n_1_737_5337), .B2(n_1_737_2886), 
      .ZN(n_1_737_2885));
   OAI21_X1 i_1_737_3220 (.A(\out_bs[0] [6]), .B1(n_1_737_5331), .B2(
      n_1_737_4686), .ZN(n_1_737_2886));
   OAI21_X1 i_1_737_3221 (.A(n_1_737_2888), .B1(n_1_737_5544), .B2(n_1_737_5365), 
      .ZN(n_1_737_2887));
   OAI21_X1 i_1_737_3222 (.A(n_1_737_2889), .B1(n_1_737_613), .B2(n_1_737_5366), 
      .ZN(n_1_737_2888));
   OAI21_X1 i_1_737_3223 (.A(\out_bs[4] [6]), .B1(n_1_737_5400), .B2(
      n_1_737_4715), .ZN(n_1_737_2889));
   NOR2_X1 i_1_737_3224 (.A1(n_1_737_608), .A2(n_1_737_2903), .ZN(n_334));
   NAND2_X1 i_1_737_3225 (.A1(n_1_737_608), .A2(n_1_737_2903), .ZN(n_335));
   NOR2_X1 i_1_737_3226 (.A1(n_1_737_607), .A2(n_1_737_2905), .ZN(n_336));
   NAND2_X1 i_1_737_3227 (.A1(n_1_737_607), .A2(n_1_737_2905), .ZN(n_337));
   NAND4_X1 i_1_737_3228 (.A1(n_1_737_2898), .A2(n_1_737_2890), .A3(n_1_737_2894), 
      .A4(n_1_737_2896), .ZN(n_338));
   AOI21_X1 i_1_737_3229 (.A(n_1_737_2891), .B1(n_1_737_2901), .B2(n_1_737_2900), 
      .ZN(n_1_737_2890));
   INV_X1 i_1_737_3230 (.A(n_1_737_2892), .ZN(n_1_737_2891));
   OAI21_X1 i_1_737_3231 (.A(n_1_737_2893), .B1(n_1_737_5550), .B2(n_1_737_5297), 
      .ZN(n_1_737_2892));
   OAI22_X1 i_1_737_3232 (.A1(n_1_737_5664), .A2(n_1_737_4749), .B1(n_1_737_603), 
      .B2(n_1_737_5298), .ZN(n_1_737_2893));
   OAI21_X1 i_1_737_3233 (.A(n_1_737_2895), .B1(n_1_737_5548), .B2(n_1_737_5189), 
      .ZN(n_1_737_2894));
   OAI22_X1 i_1_737_3234 (.A1(n_1_737_5638), .A2(n_1_737_4759), .B1(n_1_737_605), 
      .B2(n_1_737_5190), .ZN(n_1_737_2895));
   OAI22_X1 i_1_737_3235 (.A1(n_1_737_2921), .A2(n_1_737_2897), .B1(n_1_737_5547), 
      .B2(n_1_737_5365), .ZN(n_1_737_2896));
   NOR2_X1 i_1_737_3236 (.A1(n_1_737_606), .A2(n_1_737_5366), .ZN(n_1_737_2897));
   OAI21_X1 i_1_737_3237 (.A(n_1_737_2899), .B1(n_1_737_5549), .B2(n_1_737_5235), 
      .ZN(n_1_737_2898));
   OAI22_X1 i_1_737_3238 (.A1(n_1_737_5651), .A2(n_1_737_4768), .B1(n_1_737_604), 
      .B2(n_1_737_5236), .ZN(n_1_737_2899));
   NAND2_X1 i_1_737_3239 (.A1(n_1_737_602), .A2(n_1_737_5337), .ZN(n_1_737_2900));
   OAI22_X1 i_1_737_3240 (.A1(n_1_737_5671), .A2(n_1_737_4776), .B1(n_1_737_602), 
      .B2(n_1_737_5337), .ZN(n_1_737_2901));
   NOR2_X1 i_1_737_3241 (.A1(n_1_737_601), .A2(n_1_737_2902), .ZN(n_339));
   NAND2_X1 i_1_737_3242 (.A1(n_1_737_601), .A2(n_1_737_2902), .ZN(n_340));
   OAI21_X1 i_1_737_3243 (.A(\out_bs[6] [6]), .B1(\out_bs[6] [5]), .B2(
      n_1_737_3695), .ZN(n_1_737_2902));
   OAI21_X1 i_1_737_3244 (.A(\out_bs[6] [6]), .B1(\out_bs[6] [5]), .B2(
      n_1_737_3697), .ZN(n_1_737_2903));
   NOR2_X1 i_1_737_3245 (.A1(n_1_737_600), .A2(n_1_737_2904), .ZN(n_341));
   NAND2_X1 i_1_737_3246 (.A1(n_1_737_600), .A2(n_1_737_2904), .ZN(n_342));
   OAI21_X1 i_1_737_3247 (.A(n_844), .B1(n_845), .B2(n_1_737_4738), .ZN(
      n_1_737_2904));
   OAI21_X1 i_1_737_3248 (.A(n_844), .B1(n_845), .B2(n_1_737_4741), .ZN(
      n_1_737_2905));
   NAND4_X1 i_1_737_3249 (.A1(n_1_737_2911), .A2(n_1_737_2906), .A3(n_1_737_2915), 
      .A4(n_1_737_2917), .ZN(n_343));
   AOI21_X1 i_1_737_3250 (.A(n_1_737_2908), .B1(n_1_737_2923), .B2(n_1_737_2922), 
      .ZN(n_1_737_2906));
   INV_X1 i_1_737_3251 (.A(n_1_737_2908), .ZN(n_1_737_2907));
   OAI22_X1 i_1_737_3252 (.A1(n_1_737_596), .A2(n_1_737_5298), .B1(n_1_737_2910), 
      .B2(n_1_737_2909), .ZN(n_1_737_2908));
   OAI21_X1 i_1_737_3253 (.A(\out_bs[1] [6]), .B1(\out_bs[1] [5]), .B2(
      n_1_737_4751), .ZN(n_1_737_2909));
   AND2_X1 i_1_737_3254 (.A1(n_1_737_596), .A2(n_1_737_5298), .ZN(n_1_737_2910));
   INV_X1 i_1_737_3255 (.A(n_1_737_2912), .ZN(n_1_737_2911));
   OAI22_X1 i_1_737_3256 (.A1(n_1_737_597), .A2(n_1_737_5236), .B1(n_1_737_2914), 
      .B2(n_1_737_2913), .ZN(n_1_737_2912));
   OAI21_X1 i_1_737_3257 (.A(\out_bs[2] [6]), .B1(\out_bs[2] [5]), .B2(
      n_1_737_4770), .ZN(n_1_737_2913));
   AND2_X1 i_1_737_3258 (.A1(n_1_737_597), .A2(n_1_737_5236), .ZN(n_1_737_2914));
   OAI21_X1 i_1_737_3259 (.A(n_1_737_2916), .B1(n_1_737_5551), .B2(n_1_737_5189), 
      .ZN(n_1_737_2915));
   OAI221_X1 i_1_737_3260 (.A(n_1_737_3005), .B1(n_1_737_5638), .B2(n_1_737_4760), 
      .C1(n_1_737_598), .C2(n_1_737_5190), .ZN(n_1_737_2916));
   INV_X1 i_1_737_3261 (.A(n_1_737_2918), .ZN(n_1_737_2917));
   OAI22_X1 i_1_737_3262 (.A1(n_1_737_599), .A2(n_1_737_5366), .B1(n_1_737_2920), 
      .B2(n_1_737_2919), .ZN(n_1_737_2918));
   AND2_X1 i_1_737_3263 (.A1(n_1_737_599), .A2(n_1_737_5366), .ZN(n_1_737_2919));
   OAI21_X1 i_1_737_3264 (.A(\out_bs[4] [6]), .B1(\out_bs[4] [5]), .B2(
      n_1_737_4788), .ZN(n_1_737_2920));
   NOR2_X1 i_1_737_3265 (.A1(n_1_737_5625), .A2(n_1_737_4786), .ZN(n_1_737_2921));
   NAND2_X1 i_1_737_3266 (.A1(n_1_737_595), .A2(n_1_737_5337), .ZN(n_1_737_2922));
   OAI221_X1 i_1_737_3267 (.A(n_1_737_3018), .B1(n_1_737_5671), .B2(n_1_737_4777), 
      .C1(n_1_737_595), .C2(n_1_737_5337), .ZN(n_1_737_2923));
   NOR2_X1 i_1_737_3268 (.A1(n_1_737_594), .A2(n_1_737_2924), .ZN(n_344));
   NAND2_X1 i_1_737_3269 (.A1(n_1_737_594), .A2(n_1_737_2924), .ZN(n_345));
   OAI21_X1 i_1_737_3270 (.A(\out_bs[6] [6]), .B1(\out_bs[6] [5]), .B2(
      n_1_737_3750), .ZN(n_1_737_2924));
   NOR2_X1 i_1_737_3271 (.A1(n_1_737_593), .A2(n_1_737_2925), .ZN(n_346));
   NAND2_X1 i_1_737_3272 (.A1(n_1_737_593), .A2(n_1_737_2925), .ZN(n_347));
   OAI21_X1 i_1_737_3273 (.A(n_844), .B1(n_845), .B2(n_1_737_4812), .ZN(
      n_1_737_2925));
   NAND4_X1 i_1_737_3274 (.A1(n_1_737_2931), .A2(n_1_737_2926), .A3(n_1_737_2929), 
      .A4(n_1_737_2936), .ZN(n_348));
   AOI21_X1 i_1_737_3275 (.A(n_1_737_2933), .B1(n_1_737_2928), .B2(n_1_737_2927), 
      .ZN(n_1_737_2926));
   NAND2_X1 i_1_737_3276 (.A1(n_1_737_588), .A2(n_1_737_5337), .ZN(n_1_737_2927));
   OAI21_X1 i_1_737_3277 (.A(n_1_737_2956), .B1(n_1_737_588), .B2(n_1_737_5337), 
      .ZN(n_1_737_2928));
   OAI21_X1 i_1_737_3278 (.A(n_1_737_2930), .B1(n_1_737_5553), .B2(n_1_737_5189), 
      .ZN(n_1_737_2929));
   OAI21_X1 i_1_737_3279 (.A(n_1_737_2945), .B1(n_1_737_591), .B2(n_1_737_5190), 
      .ZN(n_1_737_2930));
   OAI21_X1 i_1_737_3280 (.A(n_1_737_2932), .B1(n_1_737_5554), .B2(n_1_737_5235), 
      .ZN(n_1_737_2931));
   OAI21_X1 i_1_737_3281 (.A(n_1_737_2949), .B1(n_1_737_590), .B2(n_1_737_5236), 
      .ZN(n_1_737_2932));
   AOI21_X1 i_1_737_3282 (.A(n_1_737_2934), .B1(n_1_737_589), .B2(n_1_737_5298), 
      .ZN(n_1_737_2933));
   INV_X1 i_1_737_3283 (.A(n_1_737_2935), .ZN(n_1_737_2934));
   OAI21_X1 i_1_737_3284 (.A(n_1_737_2954), .B1(n_1_737_589), .B2(n_1_737_5298), 
      .ZN(n_1_737_2935));
   OAI21_X1 i_1_737_3285 (.A(n_1_737_2937), .B1(n_1_737_5552), .B2(n_1_737_5365), 
      .ZN(n_1_737_2936));
   OAI21_X1 i_1_737_3286 (.A(n_1_737_2959), .B1(n_1_737_592), .B2(n_1_737_5366), 
      .ZN(n_1_737_2937));
   NOR2_X1 i_1_737_3287 (.A1(n_1_737_586), .A2(n_1_737_2938), .ZN(n_349));
   NAND2_X1 i_1_737_3288 (.A1(n_1_737_586), .A2(n_1_737_2938), .ZN(n_350));
   AOI211_X1 i_1_737_3289 (.A(n_1_737_3110), .B(n_1_737_3108), .C1(n_844), 
      .C2(n_1_737_4810), .ZN(n_1_737_2938));
   OR4_X1 i_1_737_3290 (.A1(n_1_737_2946), .A2(n_1_737_2939), .A3(n_1_737_2942), 
      .A4(n_1_737_2957), .ZN(n_351));
   OAI211_X1 i_1_737_3291 (.A(n_1_737_2940), .B(n_1_737_2951), .C1(n_1_737_581), 
      .C2(n_1_737_2955), .ZN(n_1_737_2939));
   INV_X1 i_1_737_3292 (.A(n_1_737_2941), .ZN(n_1_737_2940));
   AOI21_X1 i_1_737_3293 (.A(n_1_737_5337), .B1(n_1_737_581), .B2(n_1_737_2955), 
      .ZN(n_1_737_2941));
   AOI21_X1 i_1_737_3294 (.A(n_1_737_2943), .B1(n_1_737_584), .B2(n_1_737_5190), 
      .ZN(n_1_737_2942));
   AOI21_X1 i_1_737_3295 (.A(n_1_737_2944), .B1(n_1_737_5555), .B2(n_1_737_5189), 
      .ZN(n_1_737_2943));
   AOI21_X1 i_1_737_3296 (.A(n_1_737_5638), .B1(n_1_737_5637), .B2(n_1_737_4829), 
      .ZN(n_1_737_2944));
   OAI21_X1 i_1_737_3297 (.A(\out_bs[3] [6]), .B1(n_1_737_5228), .B2(
      n_1_737_4835), .ZN(n_1_737_2945));
   AOI21_X1 i_1_737_3298 (.A(n_1_737_2947), .B1(n_1_737_583), .B2(n_1_737_5236), 
      .ZN(n_1_737_2946));
   AOI21_X1 i_1_737_3299 (.A(n_1_737_2948), .B1(n_1_737_5556), .B2(n_1_737_5235), 
      .ZN(n_1_737_2947));
   AOI21_X1 i_1_737_3300 (.A(n_1_737_5651), .B1(n_1_737_5650), .B2(n_1_737_4850), 
      .ZN(n_1_737_2948));
   OAI21_X1 i_1_737_3301 (.A(\out_bs[2] [6]), .B1(n_1_737_5259), .B2(
      n_1_737_4854), .ZN(n_1_737_2949));
   INV_X1 i_1_737_3302 (.A(n_1_737_2951), .ZN(n_1_737_2950));
   OAI21_X1 i_1_737_3303 (.A(n_1_737_2952), .B1(n_1_737_5557), .B2(n_1_737_5297), 
      .ZN(n_1_737_2951));
   OAI21_X1 i_1_737_3304 (.A(n_1_737_2953), .B1(n_1_737_582), .B2(n_1_737_5298), 
      .ZN(n_1_737_2952));
   OAI21_X1 i_1_737_3305 (.A(\out_bs[1] [6]), .B1(n_1_737_5292), .B2(
      n_1_737_4841), .ZN(n_1_737_2953));
   OAI21_X1 i_1_737_3306 (.A(\out_bs[1] [6]), .B1(n_1_737_5292), .B2(
      n_1_737_4845), .ZN(n_1_737_2954));
   OAI21_X1 i_1_737_3307 (.A(\out_bs[0] [6]), .B1(n_1_737_5331), .B2(
      n_1_737_4819), .ZN(n_1_737_2955));
   OAI21_X1 i_1_737_3308 (.A(\out_bs[0] [6]), .B1(n_1_737_5331), .B2(
      n_1_737_4823), .ZN(n_1_737_2956));
   OAI22_X1 i_1_737_3309 (.A1(n_1_737_585), .A2(n_1_737_5366), .B1(n_1_737_2960), 
      .B2(n_1_737_2958), .ZN(n_1_737_2957));
   OAI21_X1 i_1_737_3310 (.A(\out_bs[4] [6]), .B1(n_1_737_5400), .B2(
      n_1_737_4860), .ZN(n_1_737_2958));
   OAI21_X1 i_1_737_3311 (.A(\out_bs[4] [6]), .B1(n_1_737_5400), .B2(
      n_1_737_4863), .ZN(n_1_737_2959));
   AND2_X1 i_1_737_3312 (.A1(n_1_737_585), .A2(n_1_737_5366), .ZN(n_1_737_2960));
   NOR2_X1 i_1_737_3313 (.A1(n_1_737_580), .A2(n_1_737_3081), .ZN(n_352));
   NAND2_X1 i_1_737_3314 (.A1(n_1_737_580), .A2(n_1_737_3081), .ZN(n_353));
   NOR2_X1 i_1_737_3315 (.A1(n_1_737_579), .A2(n_1_737_3086), .ZN(n_354));
   NAND2_X1 i_1_737_3316 (.A1(n_1_737_579), .A2(n_1_737_3086), .ZN(n_355));
   OAI211_X1 i_1_737_3317 (.A(n_1_737_2972), .B(n_1_737_2961), .C1(n_1_737_574), 
      .C2(n_1_737_3094), .ZN(n_356));
   NOR4_X1 i_1_737_3318 (.A1(n_1_737_2965), .A2(n_1_737_2962), .A3(n_1_737_2967), 
      .A4(n_1_737_2970), .ZN(n_1_737_2961));
   INV_X1 i_1_737_3319 (.A(n_1_737_2963), .ZN(n_1_737_2962));
   OAI21_X1 i_1_737_3320 (.A(n_1_737_2964), .B1(n_1_737_5559), .B2(n_1_737_5297), 
      .ZN(n_1_737_2963));
   OAI22_X1 i_1_737_3321 (.A1(n_1_737_5664), .A2(n_1_737_5291), .B1(n_1_737_575), 
      .B2(n_1_737_5298), .ZN(n_1_737_2964));
   AOI21_X1 i_1_737_3322 (.A(n_1_737_2966), .B1(n_1_737_577), .B2(n_1_737_5190), 
      .ZN(n_1_737_2965));
   AOI21_X1 i_1_737_3323 (.A(n_1_737_3101), .B1(n_1_737_5558), .B2(n_1_737_5189), 
      .ZN(n_1_737_2966));
   OAI22_X1 i_1_737_3324 (.A1(n_1_737_576), .A2(n_1_737_3091), .B1(n_1_737_5236), 
      .B2(n_1_737_2968), .ZN(n_1_737_2967));
   AND2_X1 i_1_737_3325 (.A1(n_1_737_576), .A2(n_1_737_3091), .ZN(n_1_737_2968));
   INV_X1 i_1_737_3326 (.A(n_1_737_2970), .ZN(n_1_737_2969));
   OAI22_X1 i_1_737_3327 (.A1(n_1_737_578), .A2(n_1_737_3104), .B1(n_1_737_5366), 
      .B2(n_1_737_2971), .ZN(n_1_737_2970));
   AND2_X1 i_1_737_3328 (.A1(n_1_737_578), .A2(n_1_737_3104), .ZN(n_1_737_2971));
   INV_X1 i_1_737_3329 (.A(n_1_737_2973), .ZN(n_1_737_2972));
   AOI21_X1 i_1_737_3330 (.A(n_1_737_5337), .B1(n_1_737_574), .B2(n_1_737_3094), 
      .ZN(n_1_737_2973));
   NOR2_X1 i_1_737_3331 (.A1(n_1_737_573), .A2(n_1_737_2974), .ZN(n_357));
   NAND2_X1 i_1_737_3332 (.A1(n_1_737_573), .A2(n_1_737_2974), .ZN(n_358));
   OAI21_X1 i_1_737_3333 (.A(\out_bs[6] [6]), .B1(\out_bs[6] [5]), .B2(
      n_1_737_3831), .ZN(n_1_737_2974));
   NOR2_X1 i_1_737_3334 (.A1(n_1_737_572), .A2(n_1_737_2975), .ZN(n_359));
   NAND2_X1 i_1_737_3335 (.A1(n_1_737_572), .A2(n_1_737_2975), .ZN(n_360));
   OAI21_X1 i_1_737_3336 (.A(n_844), .B1(n_845), .B2(n_1_737_4881), .ZN(
      n_1_737_2975));
   NAND3_X1 i_1_737_3337 (.A1(n_1_737_2991), .A2(n_1_737_2976), .A3(n_1_737_2994), 
      .ZN(n_361));
   NOR3_X1 i_1_737_3338 (.A1(n_1_737_2986), .A2(n_1_737_2977), .A3(n_1_737_2980), 
      .ZN(n_1_737_2976));
   AOI21_X1 i_1_737_3339 (.A(n_1_737_2978), .B1(n_1_737_567), .B2(n_1_737_5337), 
      .ZN(n_1_737_2977));
   INV_X1 i_1_737_3340 (.A(n_1_737_2979), .ZN(n_1_737_2978));
   OAI21_X1 i_1_737_3341 (.A(n_1_737_2984), .B1(n_1_737_567), .B2(n_1_737_5337), 
      .ZN(n_1_737_2979));
   AOI21_X1 i_1_737_3342 (.A(n_1_737_2981), .B1(n_1_737_569), .B2(n_1_737_5236), 
      .ZN(n_1_737_2980));
   INV_X1 i_1_737_3343 (.A(n_1_737_2982), .ZN(n_1_737_2981));
   OAI21_X1 i_1_737_3344 (.A(n_1_737_2983), .B1(n_1_737_569), .B2(n_1_737_5236), 
      .ZN(n_1_737_2982));
   OAI21_X1 i_1_737_3345 (.A(\out_bs[2] [6]), .B1(n_1_737_5258), .B2(
      n_1_737_4901), .ZN(n_1_737_2983));
   INV_X1 i_1_737_3346 (.A(n_1_737_2985), .ZN(n_1_737_2984));
   AOI21_X1 i_1_737_3347 (.A(n_1_737_5671), .B1(n_1_737_5670), .B2(n_1_737_4904), 
      .ZN(n_1_737_2985));
   INV_X1 i_1_737_3348 (.A(n_1_737_2987), .ZN(n_1_737_2986));
   OAI21_X1 i_1_737_3349 (.A(n_1_737_2988), .B1(n_1_737_5562), .B2(n_1_737_5297), 
      .ZN(n_1_737_2987));
   OAI21_X1 i_1_737_3350 (.A(n_1_737_2989), .B1(n_1_737_568), .B2(n_1_737_5298), 
      .ZN(n_1_737_2988));
   OAI21_X1 i_1_737_3351 (.A(\out_bs[1] [6]), .B1(n_1_737_5290), .B2(
      n_1_737_4890), .ZN(n_1_737_2989));
   INV_X1 i_1_737_3352 (.A(n_1_737_2991), .ZN(n_1_737_2990));
   OAI21_X1 i_1_737_3353 (.A(n_1_737_2992), .B1(n_1_737_5561), .B2(n_1_737_5189), 
      .ZN(n_1_737_2991));
   OAI21_X1 i_1_737_3354 (.A(n_1_737_2993), .B1(n_1_737_570), .B2(n_1_737_5190), 
      .ZN(n_1_737_2992));
   OAI21_X1 i_1_737_3355 (.A(\out_bs[3] [6]), .B1(n_1_737_5226), .B2(
      n_1_737_4896), .ZN(n_1_737_2993));
   OAI21_X1 i_1_737_3356 (.A(n_1_737_2995), .B1(n_1_737_5560), .B2(n_1_737_5365), 
      .ZN(n_1_737_2994));
   OAI21_X1 i_1_737_3357 (.A(n_1_737_2996), .B1(n_1_737_571), .B2(n_1_737_5366), 
      .ZN(n_1_737_2995));
   OAI21_X1 i_1_737_3358 (.A(\out_bs[4] [6]), .B1(n_1_737_5399), .B2(
      n_1_737_4912), .ZN(n_1_737_2996));
   NOR2_X1 i_1_737_3359 (.A1(n_1_737_566), .A2(n_1_737_2997), .ZN(n_362));
   NAND2_X1 i_1_737_3360 (.A1(n_1_737_566), .A2(n_1_737_2997), .ZN(n_363));
   OAI21_X1 i_1_737_3361 (.A(\out_bs[6] [6]), .B1(\out_bs[6] [5]), .B2(
      n_1_737_4917), .ZN(n_1_737_2997));
   NOR2_X1 i_1_737_3362 (.A1(n_1_737_565), .A2(n_1_737_2998), .ZN(n_364));
   NAND2_X1 i_1_737_3363 (.A1(n_1_737_565), .A2(n_1_737_2998), .ZN(n_365));
   OAI21_X1 i_1_737_3364 (.A(n_844), .B1(n_845), .B2(n_1_737_4922), .ZN(
      n_1_737_2998));
   NAND3_X1 i_1_737_3365 (.A1(n_1_737_3003), .A2(n_1_737_2999), .A3(n_1_737_3020), 
      .ZN(n_366));
   AOI211_X1 i_1_737_3366 (.A(n_1_737_3013), .B(n_1_737_3007), .C1(n_1_737_3001), 
      .C2(n_1_737_3000), .ZN(n_1_737_2999));
   NAND2_X1 i_1_737_3367 (.A1(n_1_737_560), .A2(n_1_737_5337), .ZN(n_1_737_3000));
   OAI221_X1 i_1_737_3368 (.A(n_1_737_3018), .B1(n_1_737_5671), .B2(n_1_737_4946), 
      .C1(n_1_737_560), .C2(n_1_737_5337), .ZN(n_1_737_3001));
   INV_X1 i_1_737_3369 (.A(n_1_737_3003), .ZN(n_1_737_3002));
   OAI21_X1 i_1_737_3370 (.A(n_1_737_3004), .B1(n_1_737_5564), .B2(n_1_737_5189), 
      .ZN(n_1_737_3003));
   OAI221_X1 i_1_737_3371 (.A(n_1_737_3005), .B1(n_1_737_5638), .B2(n_1_737_4939), 
      .C1(n_1_737_563), .C2(n_1_737_5190), .ZN(n_1_737_3004));
   INV_X1 i_1_737_3372 (.A(n_1_737_3006), .ZN(n_1_737_3005));
   NOR2_X1 i_1_737_3373 (.A1(n_1_737_5638), .A2(n_1_737_5637), .ZN(n_1_737_3006));
   AOI21_X1 i_1_737_3374 (.A(n_1_737_3008), .B1(n_1_737_562), .B2(n_1_737_5236), 
      .ZN(n_1_737_3007));
   INV_X1 i_1_737_3375 (.A(n_1_737_3009), .ZN(n_1_737_3008));
   OAI221_X1 i_1_737_3376 (.A(n_1_737_3010), .B1(n_1_737_5651), .B2(n_1_737_4953), 
      .C1(n_1_737_562), .C2(n_1_737_5236), .ZN(n_1_737_3009));
   INV_X1 i_1_737_3377 (.A(n_1_737_3011), .ZN(n_1_737_3010));
   NOR2_X1 i_1_737_3378 (.A1(n_1_737_5651), .A2(n_1_737_5650), .ZN(n_1_737_3011));
   INV_X1 i_1_737_3379 (.A(n_1_737_3013), .ZN(n_1_737_3012));
   OAI22_X1 i_1_737_3380 (.A1(n_1_737_561), .A2(n_1_737_5298), .B1(n_1_737_3017), 
      .B2(n_1_737_3014), .ZN(n_1_737_3013));
   OAI21_X1 i_1_737_3381 (.A(\out_bs[1] [6]), .B1(\out_bs[1] [5]), .B2(
      n_1_737_4931), .ZN(n_1_737_3014));
   INV_X1 i_1_737_3382 (.A(n_1_737_3016), .ZN(n_1_737_3015));
   NOR2_X1 i_1_737_3383 (.A1(n_1_737_5664), .A2(n_1_737_5663), .ZN(n_1_737_3016));
   AND2_X1 i_1_737_3384 (.A1(n_1_737_561), .A2(n_1_737_5298), .ZN(n_1_737_3017));
   INV_X1 i_1_737_3385 (.A(n_1_737_3019), .ZN(n_1_737_3018));
   NOR2_X1 i_1_737_3386 (.A1(n_1_737_5671), .A2(n_1_737_5670), .ZN(n_1_737_3019));
   OAI21_X1 i_1_737_3387 (.A(n_1_737_3021), .B1(n_1_737_5563), .B2(n_1_737_5365), 
      .ZN(n_1_737_3020));
   OAI221_X1 i_1_737_3388 (.A(n_1_737_3022), .B1(n_1_737_5625), .B2(n_1_737_4960), 
      .C1(n_1_737_564), .C2(n_1_737_5366), .ZN(n_1_737_3021));
   INV_X1 i_1_737_3389 (.A(n_1_737_3023), .ZN(n_1_737_3022));
   NOR2_X1 i_1_737_3390 (.A1(n_1_737_5625), .A2(n_1_737_5624), .ZN(n_1_737_3023));
   NOR2_X1 i_1_737_3391 (.A1(n_1_737_559), .A2(n_1_737_3024), .ZN(n_367));
   NAND2_X1 i_1_737_3392 (.A1(n_1_737_559), .A2(n_1_737_3024), .ZN(n_368));
   OAI21_X1 i_1_737_3393 (.A(\out_bs[6] [6]), .B1(\out_bs[6] [5]), .B2(
      n_1_737_3882), .ZN(n_1_737_3024));
   NOR2_X1 i_1_737_3394 (.A1(n_1_737_558), .A2(n_1_737_3025), .ZN(n_369));
   NAND2_X1 i_1_737_3395 (.A1(n_1_737_558), .A2(n_1_737_3025), .ZN(n_370));
   OAI21_X1 i_1_737_3396 (.A(n_844), .B1(n_845), .B2(n_1_737_4963), .ZN(
      n_1_737_3025));
   NAND4_X1 i_1_737_3397 (.A1(n_1_737_3029), .A2(n_1_737_3026), .A3(n_1_737_3037), 
      .A4(n_1_737_3040), .ZN(n_371));
   AOI21_X1 i_1_737_3398 (.A(n_1_737_3033), .B1(n_1_737_3028), .B2(n_1_737_3027), 
      .ZN(n_1_737_3026));
   NAND2_X1 i_1_737_3399 (.A1(n_1_737_553), .A2(n_1_737_5337), .ZN(n_1_737_3027));
   OAI21_X1 i_1_737_3400 (.A(n_1_737_3032), .B1(n_1_737_553), .B2(n_1_737_5337), 
      .ZN(n_1_737_3028));
   OAI21_X1 i_1_737_3401 (.A(n_1_737_3030), .B1(n_1_737_5567), .B2(n_1_737_5235), 
      .ZN(n_1_737_3029));
   OAI21_X1 i_1_737_3402 (.A(n_1_737_3031), .B1(n_1_737_555), .B2(n_1_737_5236), 
      .ZN(n_1_737_3030));
   OAI21_X1 i_1_737_3403 (.A(\out_bs[2] [6]), .B1(n_1_737_5258), .B2(
      n_1_737_4987), .ZN(n_1_737_3031));
   OAI21_X1 i_1_737_3404 (.A(\out_bs[0] [6]), .B1(n_1_737_5330), .B2(
      n_1_737_4993), .ZN(n_1_737_3032));
   INV_X1 i_1_737_3405 (.A(n_1_737_3034), .ZN(n_1_737_3033));
   OAI21_X1 i_1_737_3406 (.A(n_1_737_3035), .B1(n_1_737_5568), .B2(n_1_737_5297), 
      .ZN(n_1_737_3034));
   OAI21_X1 i_1_737_3407 (.A(n_1_737_3036), .B1(n_1_737_554), .B2(n_1_737_5298), 
      .ZN(n_1_737_3035));
   OAI21_X1 i_1_737_3408 (.A(\out_bs[1] [6]), .B1(n_1_737_5290), .B2(
      n_1_737_4972), .ZN(n_1_737_3036));
   OAI21_X1 i_1_737_3409 (.A(n_1_737_3038), .B1(n_1_737_5566), .B2(n_1_737_5189), 
      .ZN(n_1_737_3037));
   OAI21_X1 i_1_737_3410 (.A(n_1_737_3039), .B1(n_1_737_556), .B2(n_1_737_5190), 
      .ZN(n_1_737_3038));
   OAI21_X1 i_1_737_3411 (.A(\out_bs[3] [6]), .B1(n_1_737_5226), .B2(
      n_1_737_4980), .ZN(n_1_737_3039));
   OAI21_X1 i_1_737_3412 (.A(n_1_737_3041), .B1(n_1_737_5565), .B2(n_1_737_5365), 
      .ZN(n_1_737_3040));
   OAI21_X1 i_1_737_3413 (.A(n_1_737_3042), .B1(n_1_737_557), .B2(n_1_737_5366), 
      .ZN(n_1_737_3041));
   OAI21_X1 i_1_737_3414 (.A(\out_bs[4] [6]), .B1(n_1_737_5399), .B2(
      n_1_737_5001), .ZN(n_1_737_3042));
   NOR2_X1 i_1_737_3415 (.A1(n_1_737_551), .A2(n_1_737_3043), .ZN(n_372));
   NAND2_X1 i_1_737_3416 (.A1(n_1_737_551), .A2(n_1_737_3043), .ZN(n_373));
   AOI211_X1 i_1_737_3417 (.A(n_1_737_3110), .B(n_1_737_3108), .C1(n_844), 
      .C2(n_1_737_5174), .ZN(n_1_737_3043));
   NAND4_X1 i_1_737_3418 (.A1(n_1_737_3046), .A2(n_1_737_3044), .A3(n_1_737_3048), 
      .A4(n_1_737_3057), .ZN(n_374));
   OAI21_X1 i_1_737_3419 (.A(n_1_737_5572), .B1(n_1_737_5336), .B2(n_1_737_3049), 
      .ZN(n_1_737_3044));
   INV_X1 i_1_737_3420 (.A(n_1_737_3046), .ZN(n_1_737_3045));
   OAI21_X1 i_1_737_3421 (.A(n_1_737_3047), .B1(n_1_737_5570), .B2(n_1_737_5235), 
      .ZN(n_1_737_3046));
   OAI22_X1 i_1_737_3422 (.A1(n_1_737_5651), .A2(n_1_737_5255), .B1(n_1_737_548), 
      .B2(n_1_737_5236), .ZN(n_1_737_3047));
   AOI211_X1 i_1_737_3423 (.A(n_1_737_3050), .B(n_1_737_3053), .C1(n_1_737_5336), 
      .C2(n_1_737_3049), .ZN(n_1_737_3048));
   NOR2_X1 i_1_737_3424 (.A1(n_1_737_5671), .A2(n_1_737_5327), .ZN(n_1_737_3049));
   INV_X1 i_1_737_3425 (.A(n_1_737_3051), .ZN(n_1_737_3050));
   OAI21_X1 i_1_737_3426 (.A(n_1_737_3052), .B1(n_1_737_5571), .B2(n_1_737_5297), 
      .ZN(n_1_737_3051));
   OAI22_X1 i_1_737_3427 (.A1(n_1_737_5664), .A2(n_1_737_5288), .B1(n_1_737_547), 
      .B2(n_1_737_5298), .ZN(n_1_737_3052));
   AOI21_X1 i_1_737_3428 (.A(n_1_737_3054), .B1(n_1_737_549), .B2(n_1_737_5190), 
      .ZN(n_1_737_3053));
   INV_X1 i_1_737_3429 (.A(n_1_737_3055), .ZN(n_1_737_3054));
   OAI21_X1 i_1_737_3430 (.A(n_1_737_3066), .B1(n_1_737_549), .B2(n_1_737_5190), 
      .ZN(n_1_737_3055));
   INV_X1 i_1_737_3431 (.A(n_1_737_3057), .ZN(n_1_737_3056));
   OAI21_X1 i_1_737_3432 (.A(n_1_737_3058), .B1(n_1_737_5569), .B2(n_1_737_5365), 
      .ZN(n_1_737_3057));
   OAI22_X1 i_1_737_3433 (.A1(n_1_737_5625), .A2(n_1_737_5396), .B1(n_1_737_550), 
      .B2(n_1_737_5366), .ZN(n_1_737_3058));
   NOR2_X1 i_1_737_3434 (.A1(n_1_737_544), .A2(n_1_737_3059), .ZN(n_375));
   NAND2_X1 i_1_737_3435 (.A1(n_1_737_544), .A2(n_1_737_3059), .ZN(n_376));
   AOI211_X1 i_1_737_3436 (.A(n_1_737_3110), .B(n_1_737_3108), .C1(n_844), 
      .C2(n_1_737_5020), .ZN(n_1_737_3059));
   OR4_X1 i_1_737_3437 (.A1(n_1_737_3067), .A2(n_1_737_3060), .A3(n_1_737_3063), 
      .A4(n_1_737_3076), .ZN(n_377));
   OAI211_X1 i_1_737_3438 (.A(n_1_737_3061), .B(n_1_737_3072), .C1(n_1_737_539), 
      .C2(n_1_737_3075), .ZN(n_1_737_3060));
   INV_X1 i_1_737_3439 (.A(n_1_737_3062), .ZN(n_1_737_3061));
   AOI21_X1 i_1_737_3440 (.A(n_1_737_5337), .B1(n_1_737_539), .B2(n_1_737_3075), 
      .ZN(n_1_737_3062));
   INV_X1 i_1_737_3441 (.A(n_1_737_3064), .ZN(n_1_737_3063));
   OAI21_X1 i_1_737_3442 (.A(n_1_737_3065), .B1(n_1_737_5573), .B2(n_1_737_5189), 
      .ZN(n_1_737_3064));
   OAI221_X1 i_1_737_3443 (.A(n_1_737_3066), .B1(n_1_737_5638), .B2(n_1_737_5039), 
      .C1(n_1_737_542), .C2(n_1_737_5190), .ZN(n_1_737_3065));
   OAI21_X1 i_1_737_3444 (.A(\out_bs[3] [6]), .B1(\out_bs[3] [2]), .B2(
      n_1_737_5226), .ZN(n_1_737_3066));
   INV_X1 i_1_737_3445 (.A(n_1_737_3068), .ZN(n_1_737_3067));
   OAI21_X1 i_1_737_3446 (.A(n_1_737_3069), .B1(n_1_737_5574), .B2(n_1_737_5235), 
      .ZN(n_1_737_3068));
   OAI21_X1 i_1_737_3447 (.A(n_1_737_3070), .B1(n_1_737_541), .B2(n_1_737_5236), 
      .ZN(n_1_737_3069));
   OAI21_X1 i_1_737_3448 (.A(\out_bs[2] [6]), .B1(n_1_737_5259), .B2(
      n_1_737_5053), .ZN(n_1_737_3070));
   INV_X1 i_1_737_3449 (.A(n_1_737_3072), .ZN(n_1_737_3071));
   OAI21_X1 i_1_737_3450 (.A(n_1_737_3073), .B1(n_1_737_5575), .B2(n_1_737_5297), 
      .ZN(n_1_737_3072));
   OAI21_X1 i_1_737_3451 (.A(n_1_737_3074), .B1(n_1_737_540), .B2(n_1_737_5298), 
      .ZN(n_1_737_3073));
   OAI21_X1 i_1_737_3452 (.A(\out_bs[1] [6]), .B1(n_1_737_5292), .B2(
      n_1_737_5046), .ZN(n_1_737_3074));
   OAI21_X1 i_1_737_3453 (.A(\out_bs[0] [6]), .B1(n_1_737_5331), .B2(
      n_1_737_5027), .ZN(n_1_737_3075));
   OAI22_X1 i_1_737_3454 (.A1(n_1_737_543), .A2(n_1_737_5366), .B1(n_1_737_3078), 
      .B2(n_1_737_3077), .ZN(n_1_737_3076));
   OAI21_X1 i_1_737_3455 (.A(\out_bs[4] [6]), .B1(n_1_737_5400), .B2(
      n_1_737_5062), .ZN(n_1_737_3077));
   AND2_X1 i_1_737_3456 (.A1(n_1_737_543), .A2(n_1_737_5366), .ZN(n_1_737_3078));
   NOR2_X1 i_1_737_3457 (.A1(n_1_737_538), .A2(n_1_737_3079), .ZN(n_378));
   NAND2_X1 i_1_737_3458 (.A1(n_1_737_538), .A2(n_1_737_3079), .ZN(n_379));
   INV_X1 i_1_737_3459 (.A(n_1_737_3080), .ZN(n_1_737_3079));
   OAI21_X1 i_1_737_3460 (.A(n_1_737_3081), .B1(n_1_737_5607), .B2(n_1_737_4515), 
      .ZN(n_1_737_3080));
   OAI21_X1 i_1_737_3461 (.A(\out_bs[6] [6]), .B1(\out_bs[6] [5]), .B2(
      n_1_737_4918), .ZN(n_1_737_3081));
   OAI21_X1 i_1_737_3462 (.A(\out_bs[6] [6]), .B1(\out_bs[6] [5]), .B2(
      \out_bs[6] [4]), .ZN(n_1_737_3082));
   INV_X1 i_1_737_3463 (.A(n_1_737_3084), .ZN(n_1_737_3083));
   NOR2_X1 i_1_737_3464 (.A1(n_1_737_5607), .A2(n_1_737_5606), .ZN(n_1_737_3084));
   NOR2_X1 i_1_737_3465 (.A1(n_1_737_537), .A2(n_1_737_3085), .ZN(n_380));
   NAND2_X1 i_1_737_3466 (.A1(n_1_737_537), .A2(n_1_737_3085), .ZN(n_381));
   OAI21_X1 i_1_737_3467 (.A(n_844), .B1(n_845), .B2(n_1_737_5071), .ZN(
      n_1_737_3085));
   OAI21_X1 i_1_737_3468 (.A(n_844), .B1(n_845), .B2(n_1_737_5177), .ZN(
      n_1_737_3086));
   NAND4_X1 i_1_737_3469 (.A1(n_1_737_3089), .A2(n_1_737_3087), .A3(n_1_737_3092), 
      .A4(n_1_737_3102), .ZN(n_382));
   OAI21_X1 i_1_737_3470 (.A(n_1_737_5579), .B1(n_1_737_5336), .B2(n_1_737_3093), 
      .ZN(n_1_737_3087));
   INV_X1 i_1_737_3471 (.A(n_1_737_3089), .ZN(n_1_737_3088));
   OAI21_X1 i_1_737_3472 (.A(n_1_737_3090), .B1(n_1_737_5578), .B2(n_1_737_5235), 
      .ZN(n_1_737_3089));
   OAI221_X1 i_1_737_3473 (.A(n_1_737_3091), .B1(n_1_737_5651), .B2(n_1_737_5097), 
      .C1(n_1_737_534), .C2(n_1_737_5236), .ZN(n_1_737_3090));
   NAND2_X1 i_1_737_3474 (.A1(\out_bs[2] [6]), .A2(n_1_737_5258), .ZN(
      n_1_737_3091));
   AOI211_X1 i_1_737_3475 (.A(n_1_737_3096), .B(n_1_737_3099), .C1(n_1_737_5336), 
      .C2(n_1_737_3093), .ZN(n_1_737_3092));
   AOI21_X1 i_1_737_3476 (.A(n_1_737_5671), .B1(n_1_737_5670), .B2(n_1_737_5079), 
      .ZN(n_1_737_3093));
   NAND2_X1 i_1_737_3477 (.A1(\out_bs[0] [6]), .A2(n_1_737_5330), .ZN(
      n_1_737_3094));
   INV_X1 i_1_737_3478 (.A(n_1_737_3096), .ZN(n_1_737_3095));
   OAI22_X1 i_1_737_3479 (.A1(n_1_737_533), .A2(n_1_737_5298), .B1(n_1_737_3098), 
      .B2(n_1_737_3097), .ZN(n_1_737_3096));
   OAI21_X1 i_1_737_3480 (.A(\out_bs[1] [6]), .B1(n_1_737_5290), .B2(
      n_1_737_5112), .ZN(n_1_737_3097));
   AND2_X1 i_1_737_3481 (.A1(n_1_737_533), .A2(n_1_737_5298), .ZN(n_1_737_3098));
   AOI21_X1 i_1_737_3482 (.A(n_1_737_3100), .B1(n_1_737_535), .B2(n_1_737_5190), 
      .ZN(n_1_737_3099));
   AOI221_X1 i_1_737_3483 (.A(n_1_737_3101), .B1(\out_bs[3] [6]), .B2(
      n_1_737_5123), .C1(n_1_737_5577), .C2(n_1_737_5189), .ZN(n_1_737_3100));
   NOR2_X1 i_1_737_3484 (.A1(n_1_737_5638), .A2(n_1_737_5227), .ZN(n_1_737_3101));
   OAI21_X1 i_1_737_3485 (.A(n_1_737_3103), .B1(n_1_737_5576), .B2(n_1_737_5365), 
      .ZN(n_1_737_3102));
   OAI221_X1 i_1_737_3486 (.A(n_1_737_3104), .B1(n_1_737_5625), .B2(n_1_737_5132), 
      .C1(n_1_737_536), .C2(n_1_737_5366), .ZN(n_1_737_3103));
   NAND2_X1 i_1_737_3487 (.A1(\out_bs[4] [6]), .A2(n_1_737_5399), .ZN(
      n_1_737_3104));
   NOR2_X1 i_1_737_3488 (.A1(n_1_737_530), .A2(n_1_737_3105), .ZN(n_383));
   NAND2_X1 i_1_737_3489 (.A1(n_1_737_530), .A2(n_1_737_3105), .ZN(n_384));
   AOI211_X1 i_1_737_3490 (.A(n_1_737_3110), .B(n_1_737_3108), .C1(n_844), 
      .C2(n_1_737_5172), .ZN(n_1_737_3105));
   NOR2_X1 i_1_737_3491 (.A1(n_1_737_3110), .A2(n_1_737_3108), .ZN(n_1_737_3106));
   INV_X1 i_1_737_3492 (.A(n_1_737_3108), .ZN(n_1_737_3107));
   NOR2_X1 i_1_737_3493 (.A1(n_1_737_5612), .A2(n_1_737_5610), .ZN(n_1_737_3108));
   INV_X1 i_1_737_3494 (.A(n_1_737_3110), .ZN(n_1_737_3109));
   NAND3_X1 i_1_737_3496 (.A1(n_1_737_3113), .A2(n_1_737_3111), .A3(n_1_737_3127), 
      .ZN(n_385));
   NOR3_X1 i_1_737_3497 (.A1(n_1_737_3125), .A2(n_1_737_3120), .A3(n_1_737_3116), 
      .ZN(n_1_737_3111));
   INV_X1 i_1_737_3498 (.A(n_1_737_3113), .ZN(n_1_737_3112));
   OAI21_X1 i_1_737_3499 (.A(n_1_737_3114), .B1(n_1_737_5581), .B2(n_1_737_5189), 
      .ZN(n_1_737_3113));
   OAI21_X1 i_1_737_3500 (.A(n_1_737_3115), .B1(n_1_737_528), .B2(n_1_737_5190), 
      .ZN(n_1_737_3114));
   OAI21_X1 i_1_737_3501 (.A(\out_bs[3] [6]), .B1(n_1_737_5228), .B2(
      n_1_737_5223), .ZN(n_1_737_3115));
   AOI21_X1 i_1_737_3502 (.A(n_1_737_3117), .B1(n_1_737_527), .B2(n_1_737_5236), 
      .ZN(n_1_737_3116));
   INV_X1 i_1_737_3503 (.A(n_1_737_3118), .ZN(n_1_737_3117));
   OAI21_X1 i_1_737_3504 (.A(n_1_737_3119), .B1(n_1_737_527), .B2(n_1_737_5236), 
      .ZN(n_1_737_3118));
   OAI21_X1 i_1_737_3505 (.A(\out_bs[2] [6]), .B1(n_1_737_5259), .B2(
      n_1_737_5254), .ZN(n_1_737_3119));
   OAI21_X1 i_1_737_3506 (.A(n_1_737_3122), .B1(n_1_737_5337), .B2(n_1_737_3126), 
      .ZN(n_1_737_3120));
   INV_X1 i_1_737_3507 (.A(n_1_737_3122), .ZN(n_1_737_3121));
   OAI21_X1 i_1_737_3508 (.A(n_1_737_3123), .B1(n_1_737_5582), .B2(n_1_737_5297), 
      .ZN(n_1_737_3122));
   OAI21_X1 i_1_737_3509 (.A(n_1_737_3124), .B1(n_1_737_526), .B2(n_1_737_5298), 
      .ZN(n_1_737_3123));
   OAI21_X1 i_1_737_3510 (.A(\out_bs[1] [6]), .B1(n_1_737_5292), .B2(
      n_1_737_5287), .ZN(n_1_737_3124));
   AOI21_X1 i_1_737_3511 (.A(n_1_737_525), .B1(n_1_737_5337), .B2(n_1_737_3126), 
      .ZN(n_1_737_3125));
   OAI21_X1 i_1_737_3512 (.A(\out_bs[0] [6]), .B1(n_1_737_5331), .B2(
      n_1_737_5326), .ZN(n_1_737_3126));
   OAI21_X1 i_1_737_3513 (.A(n_1_737_3128), .B1(n_1_737_5580), .B2(n_1_737_5365), 
      .ZN(n_1_737_3127));
   OAI21_X1 i_1_737_3514 (.A(n_1_737_3129), .B1(n_1_737_529), .B2(n_1_737_5366), 
      .ZN(n_1_737_3128));
   OAI21_X1 i_1_737_3515 (.A(\out_bs[4] [6]), .B1(n_1_737_5400), .B2(
      n_1_737_5394), .ZN(n_1_737_3129));
   NOR2_X1 i_1_737_3516 (.A1(n_1_737_5607), .A2(n_1_737_524), .ZN(n_386));
   NAND2_X1 i_1_737_3517 (.A1(n_1_737_5607), .A2(n_1_737_524), .ZN(n_387));
   NOR2_X1 i_1_737_3518 (.A1(n_1_737_5612), .A2(n_1_737_523), .ZN(n_388));
   NAND2_X1 i_1_737_3519 (.A1(n_1_737_5612), .A2(n_1_737_523), .ZN(n_389));
   NAND2_X1 i_1_737_3520 (.A1(n_1_737_3135), .A2(n_1_737_3130), .ZN(n_390));
   AOI21_X1 i_1_737_3521 (.A(n_1_737_3133), .B1(n_1_737_3132), .B2(n_1_737_3131), 
      .ZN(n_1_737_3130));
   OAI21_X1 i_1_737_3522 (.A(n_1_737_5337), .B1(n_1_737_518), .B2(n_1_737_5338), 
      .ZN(n_1_737_3131));
   NAND2_X1 i_1_737_3523 (.A1(n_1_737_5671), .A2(n_1_737_518), .ZN(n_1_737_3132));
   OAI21_X1 i_1_737_3524 (.A(n_1_737_3134), .B1(n_1_737_522), .B2(n_1_737_5367), 
      .ZN(n_1_737_3133));
   OAI21_X1 i_1_737_3525 (.A(n_1_737_5365), .B1(\out_bs[4] [6]), .B2(
      n_1_737_5583), .ZN(n_1_737_3134));
   NOR3_X1 i_1_737_3526 (.A1(n_1_737_3141), .A2(n_1_737_3137), .A3(n_1_737_3139), 
      .ZN(n_1_737_3135));
   INV_X1 i_1_737_3527 (.A(n_1_737_3137), .ZN(n_1_737_3136));
   OAI21_X1 i_1_737_3528 (.A(n_1_737_3138), .B1(n_1_737_519), .B2(n_1_737_5299), 
      .ZN(n_1_737_3137));
   OAI21_X1 i_1_737_3529 (.A(n_1_737_5297), .B1(\out_bs[1] [6]), .B2(
      n_1_737_5586), .ZN(n_1_737_3138));
   OAI21_X1 i_1_737_3530 (.A(n_1_737_3140), .B1(n_1_737_521), .B2(n_1_737_5191), 
      .ZN(n_1_737_3139));
   OAI21_X1 i_1_737_3531 (.A(n_1_737_5189), .B1(\out_bs[3] [6]), .B2(
      n_1_737_5584), .ZN(n_1_737_3140));
   OAI21_X1 i_1_737_3532 (.A(n_1_737_3142), .B1(n_1_737_520), .B2(n_1_737_5237), 
      .ZN(n_1_737_3141));
   OAI21_X1 i_1_737_3533 (.A(n_1_737_5235), .B1(\out_bs[2] [6]), .B2(
      n_1_737_5585), .ZN(n_1_737_3142));
   NOR2_X1 i_1_737_3534 (.A1(\out_as[6] [6]), .A2(n_1_737_3143), .ZN(n_391));
   NAND2_X1 i_1_737_3535 (.A1(\out_as[6] [6]), .A2(n_1_737_3143), .ZN(n_392));
   AOI21_X1 i_1_737_3536 (.A(\out_bs[6] [6]), .B1(n_1_737_3940), .B2(
      n_1_737_3223), .ZN(n_1_737_3143));
   NOR2_X1 i_1_737_3537 (.A1(\out_as[5] [6]), .A2(n_1_737_3144), .ZN(n_393));
   NAND2_X1 i_1_737_3538 (.A1(\out_as[5] [6]), .A2(n_1_737_3144), .ZN(n_394));
   AOI21_X1 i_1_737_3539 (.A(n_844), .B1(n_845), .B2(n_1_737_4092), .ZN(
      n_1_737_3144));
   NAND4_X1 i_1_737_3540 (.A1(n_1_737_3156), .A2(n_1_737_3145), .A3(n_1_737_3147), 
      .A4(n_1_737_3165), .ZN(n_395));
   INV_X1 i_1_737_3541 (.A(n_1_737_3146), .ZN(n_1_737_3145));
   OAI211_X1 i_1_737_3542 (.A(n_1_737_3161), .B(n_1_737_3151), .C1(
      \out_as[0] [6]), .C2(n_1_737_5337), .ZN(n_1_737_3146));
   AOI22_X1 i_1_737_3543 (.A1(n_1_737_5631), .A2(n_1_737_3149), .B1(n_1_737_5189), 
      .B2(n_1_737_3148), .ZN(n_1_737_3147));
   NAND3_X1 i_1_737_3544 (.A1(n_1_737_5638), .A2(n_1_737_3150), .A3(
      \out_as[3] [6]), .ZN(n_1_737_3148));
   NAND2_X1 i_1_737_3545 (.A1(n_1_737_5638), .A2(n_1_737_3150), .ZN(n_1_737_3149));
   NAND2_X1 i_1_737_3546 (.A1(\out_bs[3] [5]), .A2(n_1_737_4113), .ZN(
      n_1_737_3150));
   INV_X1 i_1_737_3547 (.A(n_1_737_3152), .ZN(n_1_737_3151));
   OAI21_X1 i_1_737_3548 (.A(n_1_737_3153), .B1(\out_as[1] [6]), .B2(
      n_1_737_5298), .ZN(n_1_737_3152));
   OAI21_X1 i_1_737_3549 (.A(n_1_737_3154), .B1(n_1_737_5658), .B2(n_1_737_5297), 
      .ZN(n_1_737_3153));
   NAND2_X1 i_1_737_3550 (.A1(n_1_737_5664), .A2(n_1_737_3155), .ZN(n_1_737_3154));
   NAND2_X1 i_1_737_3551 (.A1(\out_bs[1] [5]), .A2(n_1_737_4118), .ZN(
      n_1_737_3155));
   OAI21_X1 i_1_737_3552 (.A(n_1_737_3157), .B1(n_1_737_5235), .B2(n_1_737_3159), 
      .ZN(n_1_737_3156));
   OAI21_X1 i_1_737_3553 (.A(\out_as[2] [6]), .B1(n_1_737_5236), .B2(
      n_1_737_3158), .ZN(n_1_737_3157));
   INV_X1 i_1_737_3554 (.A(n_1_737_3159), .ZN(n_1_737_3158));
   NAND2_X1 i_1_737_3555 (.A1(n_1_737_5651), .A2(n_1_737_3160), .ZN(n_1_737_3159));
   NAND2_X1 i_1_737_3556 (.A1(\out_bs[2] [5]), .A2(n_1_737_4108), .ZN(
      n_1_737_3160));
   OAI22_X1 i_1_737_3557 (.A1(\out_bs[0] [6]), .A2(n_1_737_3162), .B1(
      n_1_737_5678), .B2(n_1_737_5336), .ZN(n_1_737_3161));
   INV_X1 i_1_737_3558 (.A(n_1_737_3163), .ZN(n_1_737_3162));
   NAND2_X1 i_1_737_3559 (.A1(\out_bs[0] [5]), .A2(n_1_737_4096), .ZN(
      n_1_737_3163));
   INV_X1 i_1_737_3560 (.A(n_1_737_3165), .ZN(n_1_737_3164));
   OAI21_X1 i_1_737_3561 (.A(n_1_737_3166), .B1(n_1_737_5365), .B2(n_1_737_3168), 
      .ZN(n_1_737_3165));
   OAI21_X1 i_1_737_3562 (.A(\out_as[4] [6]), .B1(n_1_737_5366), .B2(
      n_1_737_3167), .ZN(n_1_737_3166));
   INV_X1 i_1_737_3563 (.A(n_1_737_3168), .ZN(n_1_737_3167));
   NAND2_X1 i_1_737_3564 (.A1(n_1_737_5625), .A2(n_1_737_3169), .ZN(n_1_737_3168));
   NAND2_X1 i_1_737_3565 (.A1(\out_bs[4] [5]), .A2(n_1_737_4101), .ZN(
      n_1_737_3169));
   NOR3_X1 i_1_737_3566 (.A1(\out_as[6] [6]), .A2(n_1_737_517), .A3(n_1_737_3170), 
      .ZN(n_396));
   OAI21_X1 i_1_737_3567 (.A(n_1_737_3170), .B1(\out_as[6] [6]), .B2(n_1_737_517), 
      .ZN(n_397));
   AOI21_X1 i_1_737_3568 (.A(\out_bs[6] [6]), .B1(n_1311), .B2(n_1_737_3222), 
      .ZN(n_1_737_3170));
   NOR3_X1 i_1_737_3569 (.A1(\out_as[5] [6]), .A2(n_1_737_516), .A3(n_1_737_3171), 
      .ZN(n_398));
   OAI21_X1 i_1_737_3570 (.A(n_1_737_3171), .B1(\out_as[5] [6]), .B2(n_1_737_516), 
      .ZN(n_399));
   AOI21_X1 i_1_737_3571 (.A(n_844), .B1(n_845), .B2(n_1_737_4120), .ZN(
      n_1_737_3171));
   NAND4_X1 i_1_737_3572 (.A1(n_1_737_3178), .A2(n_1_737_3172), .A3(n_1_737_3186), 
      .A4(n_1_737_3190), .ZN(n_400));
   AOI211_X1 i_1_737_3573 (.A(n_1_737_3183), .B(n_1_737_3173), .C1(n_1_737_5336), 
      .C2(n_1_737_3185), .ZN(n_1_737_3172));
   INV_X1 i_1_737_3574 (.A(n_1_737_3174), .ZN(n_1_737_3173));
   OAI22_X1 i_1_737_3575 (.A1(n_1_737_3177), .A2(n_1_737_3175), .B1(n_1_737_5297), 
      .B2(n_1_737_3176), .ZN(n_1_737_3174));
   AND2_X1 i_1_737_3576 (.A1(n_1_737_5297), .A2(n_1_737_3176), .ZN(n_1_737_3175));
   NOR2_X1 i_1_737_3577 (.A1(\out_as[1] [6]), .A2(n_1_737_512), .ZN(n_1_737_3176));
   OAI21_X1 i_1_737_3578 (.A(n_1_737_5664), .B1(n_1_737_4653), .B2(n_1_737_3788), 
      .ZN(n_1_737_3177));
   AOI22_X1 i_1_737_3579 (.A1(n_1_737_3182), .A2(n_1_737_3180), .B1(n_1_737_5189), 
      .B2(n_1_737_3179), .ZN(n_1_737_3178));
   OAI21_X1 i_1_737_3580 (.A(n_1_737_3181), .B1(\out_as[3] [6]), .B2(n_1_737_514), 
      .ZN(n_1_737_3179));
   INV_X1 i_1_737_3581 (.A(n_1_737_3181), .ZN(n_1_737_3180));
   AOI21_X1 i_1_737_3582 (.A(\out_bs[3] [6]), .B1(\out_bs[3] [5]), .B2(
      n_1_737_4132), .ZN(n_1_737_3181));
   NOR2_X1 i_1_737_3583 (.A1(\out_as[3] [6]), .A2(n_1_737_514), .ZN(n_1_737_3182));
   AOI221_X1 i_1_737_3584 (.A(n_1_737_3426), .B1(n_1_737_5671), .B2(n_1_737_4947), 
      .C1(n_1_737_5337), .C2(n_1_737_3184), .ZN(n_1_737_3183));
   INV_X1 i_1_737_3585 (.A(n_1_737_3185), .ZN(n_1_737_3184));
   NOR2_X1 i_1_737_3586 (.A1(\out_as[0] [6]), .A2(n_1_737_511), .ZN(n_1_737_3185));
   OAI21_X1 i_1_737_3587 (.A(n_1_737_3187), .B1(n_1_737_5235), .B2(n_1_737_3188), 
      .ZN(n_1_737_3186));
   OAI22_X1 i_1_737_3588 (.A1(\out_as[2] [6]), .A2(n_1_737_513), .B1(
      n_1_737_5236), .B2(n_1_737_3189), .ZN(n_1_737_3187));
   INV_X1 i_1_737_3589 (.A(n_1_737_3189), .ZN(n_1_737_3188));
   AOI21_X1 i_1_737_3590 (.A(\out_bs[2] [6]), .B1(\out_bs[2] [5]), .B2(
      n_1_737_4143), .ZN(n_1_737_3189));
   OAI21_X1 i_1_737_3591 (.A(n_1_737_3191), .B1(n_1_737_5365), .B2(n_1_737_3192), 
      .ZN(n_1_737_3190));
   OAI22_X1 i_1_737_3592 (.A1(\out_as[4] [6]), .A2(n_1_737_515), .B1(
      n_1_737_5366), .B2(n_1_737_3193), .ZN(n_1_737_3191));
   INV_X1 i_1_737_3593 (.A(n_1_737_3193), .ZN(n_1_737_3192));
   AOI21_X1 i_1_737_3594 (.A(\out_bs[4] [6]), .B1(\out_bs[4] [5]), .B2(
      n_1_737_4150), .ZN(n_1_737_3193));
   NOR3_X1 i_1_737_3595 (.A1(\out_as[6] [6]), .A2(n_1_737_510), .A3(n_1_737_3194), 
      .ZN(n_401));
   OAI21_X1 i_1_737_3596 (.A(n_1_737_3194), .B1(\out_as[6] [6]), .B2(n_1_737_510), 
      .ZN(n_402));
   AOI21_X1 i_1_737_3597 (.A(\out_bs[6] [6]), .B1(\out_bs[6] [5]), .B2(
      n_1_737_3195), .ZN(n_1_737_3194));
   NOR2_X1 i_1_737_3598 (.A1(n_1_737_3884), .A2(n_1_737_3331), .ZN(n_1_737_3195));
   NOR3_X1 i_1_737_3599 (.A1(\out_as[5] [6]), .A2(n_1_737_509), .A3(n_1_737_3196), 
      .ZN(n_403));
   OAI21_X1 i_1_737_3600 (.A(n_1_737_3196), .B1(\out_as[5] [6]), .B2(n_1_737_509), 
      .ZN(n_404));
   AOI21_X1 i_1_737_3601 (.A(n_844), .B1(n_845), .B2(n_1_737_4153), .ZN(
      n_1_737_3196));
   NAND3_X1 i_1_737_3602 (.A1(n_1_737_3211), .A2(n_1_737_3202), .A3(n_1_737_3197), 
      .ZN(n_405));
   NOR3_X1 i_1_737_3603 (.A1(n_1_737_3206), .A2(n_1_737_3198), .A3(n_1_737_3216), 
      .ZN(n_1_737_3197));
   OAI21_X1 i_1_737_3604 (.A(n_1_737_3199), .B1(n_1_737_5337), .B2(n_1_737_3200), 
      .ZN(n_1_737_3198));
   OAI221_X1 i_1_737_3605 (.A(n_1_737_3764), .B1(\out_bs[0] [6]), .B2(
      n_1_737_4686), .C1(n_1_737_5336), .C2(n_1_737_3201), .ZN(n_1_737_3199));
   INV_X1 i_1_737_3606 (.A(n_1_737_3201), .ZN(n_1_737_3200));
   NOR2_X1 i_1_737_3607 (.A1(\out_as[0] [6]), .A2(n_1_737_504), .ZN(n_1_737_3201));
   OAI21_X1 i_1_737_3608 (.A(n_1_737_3203), .B1(n_1_737_5235), .B2(n_1_737_3205), 
      .ZN(n_1_737_3202));
   INV_X1 i_1_737_3609 (.A(n_1_737_3204), .ZN(n_1_737_3203));
   AOI221_X1 i_1_737_3610 (.A(\out_bs[2] [6]), .B1(\out_bs[2] [5]), .B2(
      n_1_737_4178), .C1(n_1_737_5235), .C2(n_1_737_3205), .ZN(n_1_737_3204));
   NOR2_X1 i_1_737_3611 (.A1(\out_as[2] [6]), .A2(n_1_737_506), .ZN(n_1_737_3205));
   INV_X1 i_1_737_3612 (.A(n_1_737_3207), .ZN(n_1_737_3206));
   OAI21_X1 i_1_737_3613 (.A(n_1_737_3208), .B1(n_1_737_5297), .B2(n_1_737_3210), 
      .ZN(n_1_737_3207));
   INV_X1 i_1_737_3614 (.A(n_1_737_3209), .ZN(n_1_737_3208));
   AOI221_X1 i_1_737_3615 (.A(\out_bs[1] [6]), .B1(\out_bs[1] [5]), .B2(
      n_1_737_4172), .C1(n_1_737_5297), .C2(n_1_737_3210), .ZN(n_1_737_3209));
   NOR2_X1 i_1_737_3616 (.A1(\out_as[1] [6]), .A2(n_1_737_505), .ZN(n_1_737_3210));
   OAI21_X1 i_1_737_3617 (.A(n_1_737_3212), .B1(n_1_737_5189), .B2(n_1_737_3213), 
      .ZN(n_1_737_3211));
   OAI22_X1 i_1_737_3618 (.A1(\out_as[3] [6]), .A2(n_1_737_507), .B1(
      n_1_737_5190), .B2(n_1_737_3214), .ZN(n_1_737_3212));
   INV_X1 i_1_737_3619 (.A(n_1_737_3214), .ZN(n_1_737_3213));
   AOI21_X1 i_1_737_3620 (.A(\out_bs[3] [6]), .B1(\out_bs[3] [5]), .B2(
      n_1_737_4164), .ZN(n_1_737_3214));
   INV_X1 i_1_737_3621 (.A(n_1_737_3216), .ZN(n_1_737_3215));
   OAI21_X1 i_1_737_3622 (.A(n_1_737_3217), .B1(n_1_737_5366), .B2(n_1_737_3218), 
      .ZN(n_1_737_3216));
   OAI21_X1 i_1_737_3623 (.A(n_1_737_3220), .B1(n_1_737_5365), .B2(n_1_737_3219), 
      .ZN(n_1_737_3217));
   INV_X1 i_1_737_3624 (.A(n_1_737_3219), .ZN(n_1_737_3218));
   NOR2_X1 i_1_737_3625 (.A1(\out_as[4] [6]), .A2(n_1_737_508), .ZN(n_1_737_3219));
   OAI21_X1 i_1_737_3626 (.A(n_1_737_5625), .B1(n_1_737_5000), .B2(n_1_737_3457), 
      .ZN(n_1_737_3220));
   NOR3_X1 i_1_737_3627 (.A1(\out_as[6] [6]), .A2(n_1_737_503), .A3(n_1_737_3221), 
      .ZN(n_406));
   OAI21_X1 i_1_737_3628 (.A(n_1_737_3221), .B1(\out_as[6] [6]), .B2(n_1_737_503), 
      .ZN(n_407));
   NOR2_X1 i_1_737_3629 (.A1(\out_bs[6] [6]), .A2(n_1_737_3222), .ZN(
      n_1_737_3221));
   AND2_X1 i_1_737_3630 (.A1(\out_bs[6] [5]), .A2(n_1_737_3223), .ZN(
      n_1_737_3222));
   NOR2_X1 i_1_737_3631 (.A1(n_1_737_5603), .A2(n_1_737_3331), .ZN(n_1_737_3223));
   NOR3_X1 i_1_737_3632 (.A1(\out_as[5] [6]), .A2(n_1_737_502), .A3(n_1_737_3224), 
      .ZN(n_408));
   OAI21_X1 i_1_737_3633 (.A(n_1_737_3224), .B1(\out_as[5] [6]), .B2(n_1_737_502), 
      .ZN(n_409));
   AOI21_X1 i_1_737_3634 (.A(n_844), .B1(n_845), .B2(n_1_737_4209), .ZN(
      n_1_737_3224));
   OAI211_X1 i_1_737_3635 (.A(n_1_737_3226), .B(n_1_737_3225), .C1(n_1_737_5337), 
      .C2(n_1_737_3237), .ZN(n_410));
   AND4_X1 i_1_737_3636 (.A1(n_1_737_3232), .A2(n_1_737_3228), .A3(n_1_737_3243), 
      .A4(n_1_737_3239), .ZN(n_1_737_3225));
   OAI221_X1 i_1_737_3637 (.A(n_1_737_3764), .B1(\out_bs[0] [6]), .B2(
      n_1_737_4780), .C1(n_1_737_5336), .C2(n_1_737_3238), .ZN(n_1_737_3226));
   INV_X1 i_1_737_3638 (.A(n_1_737_3228), .ZN(n_1_737_3227));
   OAI22_X1 i_1_737_3639 (.A1(n_1_737_3231), .A2(n_1_737_3229), .B1(n_1_737_5297), 
      .B2(n_1_737_3230), .ZN(n_1_737_3228));
   AND2_X1 i_1_737_3640 (.A1(n_1_737_5297), .A2(n_1_737_3230), .ZN(n_1_737_3229));
   NOR2_X1 i_1_737_3641 (.A1(\out_as[1] [6]), .A2(n_1_737_498), .ZN(n_1_737_3230));
   OAI21_X1 i_1_737_3642 (.A(n_1_737_5664), .B1(n_1_737_5663), .B2(n_1_737_4218), 
      .ZN(n_1_737_3231));
   AOI22_X1 i_1_737_3643 (.A1(n_1_737_3236), .A2(n_1_737_3234), .B1(n_1_737_5365), 
      .B2(n_1_737_3233), .ZN(n_1_737_3232));
   OAI21_X1 i_1_737_3644 (.A(n_1_737_3235), .B1(\out_as[4] [6]), .B2(n_1_737_501), 
      .ZN(n_1_737_3233));
   INV_X1 i_1_737_3645 (.A(n_1_737_3235), .ZN(n_1_737_3234));
   AOI21_X1 i_1_737_3646 (.A(\out_bs[4] [6]), .B1(\out_bs[4] [5]), .B2(
      n_1_737_4253), .ZN(n_1_737_3235));
   NOR2_X1 i_1_737_3647 (.A1(\out_as[4] [6]), .A2(n_1_737_501), .ZN(n_1_737_3236));
   INV_X1 i_1_737_3648 (.A(n_1_737_3238), .ZN(n_1_737_3237));
   NOR2_X1 i_1_737_3649 (.A1(\out_as[0] [6]), .A2(n_1_737_497), .ZN(n_1_737_3238));
   AOI22_X1 i_1_737_3650 (.A1(n_1_737_3242), .A2(n_1_737_3241), .B1(n_1_737_5235), 
      .B2(n_1_737_3240), .ZN(n_1_737_3239));
   OR2_X1 i_1_737_3651 (.A1(n_1_737_3242), .A2(n_1_737_3241), .ZN(n_1_737_3240));
   OAI21_X1 i_1_737_3652 (.A(n_1_737_5651), .B1(n_1_737_5650), .B2(n_1_737_4234), 
      .ZN(n_1_737_3241));
   NOR2_X1 i_1_737_3653 (.A1(\out_as[2] [6]), .A2(n_1_737_499), .ZN(n_1_737_3242));
   AOI22_X1 i_1_737_3654 (.A1(n_1_737_3246), .A2(n_1_737_3245), .B1(n_1_737_5189), 
      .B2(n_1_737_3244), .ZN(n_1_737_3243));
   OR2_X1 i_1_737_3655 (.A1(n_1_737_3246), .A2(n_1_737_3245), .ZN(n_1_737_3244));
   OAI21_X1 i_1_737_3656 (.A(n_1_737_5638), .B1(n_1_737_5637), .B2(n_1_737_4225), 
      .ZN(n_1_737_3245));
   NOR2_X1 i_1_737_3657 (.A1(\out_as[3] [6]), .A2(n_1_737_500), .ZN(n_1_737_3246));
   NOR3_X1 i_1_737_3658 (.A1(\out_as[6] [6]), .A2(n_1_737_496), .A3(n_1_737_3247), 
      .ZN(n_411));
   OAI21_X1 i_1_737_3659 (.A(n_1_737_3247), .B1(\out_as[6] [6]), .B2(n_1_737_496), 
      .ZN(n_412));
   OAI21_X1 i_1_737_3660 (.A(n_1_737_3328), .B1(\out_bs[6] [6]), .B2(
      n_1_737_3942), .ZN(n_1_737_3247));
   NOR3_X1 i_1_737_3661 (.A1(\out_as[5] [6]), .A2(n_1_737_495), .A3(n_1_737_3248), 
      .ZN(n_413));
   OAI21_X1 i_1_737_3662 (.A(n_1_737_3248), .B1(\out_as[5] [6]), .B2(n_1_737_495), 
      .ZN(n_414));
   AOI21_X1 i_1_737_3663 (.A(n_844), .B1(n_845), .B2(n_1_737_4206), .ZN(
      n_1_737_3248));
   OR3_X1 i_1_737_3664 (.A1(n_1_737_3264), .A2(n_1_737_3254), .A3(n_1_737_3249), 
      .ZN(n_415));
   OAI211_X1 i_1_737_3665 (.A(n_1_737_3269), .B(n_1_737_3258), .C1(n_1_737_3251), 
      .C2(n_1_737_3250), .ZN(n_1_737_3249));
   NOR2_X1 i_1_737_3666 (.A1(n_1_737_3253), .A2(n_1_737_3252), .ZN(n_1_737_3250));
   AOI21_X1 i_1_737_3667 (.A(n_1_737_5336), .B1(n_1_737_3253), .B2(n_1_737_3252), 
      .ZN(n_1_737_3251));
   NOR2_X1 i_1_737_3668 (.A1(\out_as[0] [6]), .A2(n_1_737_490), .ZN(n_1_737_3252));
   OAI21_X1 i_1_737_3669 (.A(n_1_737_5671), .B1(n_1_737_5670), .B2(n_1_737_4242), 
      .ZN(n_1_737_3253));
   AOI21_X1 i_1_737_3670 (.A(n_1_737_3255), .B1(n_1_737_5190), .B2(n_1_737_3257), 
      .ZN(n_1_737_3254));
   INV_X1 i_1_737_3671 (.A(n_1_737_3256), .ZN(n_1_737_3255));
   OAI22_X1 i_1_737_3672 (.A1(\out_as[3] [6]), .A2(n_1_737_493), .B1(
      n_1_737_5190), .B2(n_1_737_3257), .ZN(n_1_737_3256));
   AOI21_X1 i_1_737_3673 (.A(\out_bs[3] [6]), .B1(\out_bs[3] [5]), .B2(
      n_1_737_4223), .ZN(n_1_737_3257));
   INV_X1 i_1_737_3674 (.A(n_1_737_3259), .ZN(n_1_737_3258));
   OAI21_X1 i_1_737_3675 (.A(n_1_737_3260), .B1(n_1_737_5298), .B2(n_1_737_3261), 
      .ZN(n_1_737_3259));
   OAI21_X1 i_1_737_3676 (.A(n_1_737_3263), .B1(n_1_737_5297), .B2(n_1_737_3262), 
      .ZN(n_1_737_3260));
   INV_X1 i_1_737_3677 (.A(n_1_737_3262), .ZN(n_1_737_3261));
   NOR2_X1 i_1_737_3678 (.A1(\out_as[1] [6]), .A2(n_1_737_491), .ZN(n_1_737_3262));
   OAI21_X1 i_1_737_3679 (.A(n_1_737_5664), .B1(n_1_737_5663), .B2(n_1_737_4216), 
      .ZN(n_1_737_3263));
   OAI21_X1 i_1_737_3680 (.A(n_1_737_3265), .B1(n_1_737_5236), .B2(n_1_737_3266), 
      .ZN(n_1_737_3264));
   OAI21_X1 i_1_737_3681 (.A(n_1_737_3268), .B1(n_1_737_5235), .B2(n_1_737_3267), 
      .ZN(n_1_737_3265));
   INV_X1 i_1_737_3682 (.A(n_1_737_3267), .ZN(n_1_737_3266));
   NOR2_X1 i_1_737_3683 (.A1(\out_as[2] [6]), .A2(n_1_737_492), .ZN(n_1_737_3267));
   OAI21_X1 i_1_737_3684 (.A(n_1_737_5651), .B1(n_1_737_5650), .B2(n_1_737_4231), 
      .ZN(n_1_737_3268));
   INV_X1 i_1_737_3685 (.A(n_1_737_3270), .ZN(n_1_737_3269));
   OAI21_X1 i_1_737_3686 (.A(n_1_737_3271), .B1(n_1_737_5366), .B2(n_1_737_3272), 
      .ZN(n_1_737_3270));
   OAI21_X1 i_1_737_3687 (.A(n_1_737_3274), .B1(n_1_737_5365), .B2(n_1_737_3273), 
      .ZN(n_1_737_3271));
   INV_X1 i_1_737_3688 (.A(n_1_737_3273), .ZN(n_1_737_3272));
   NOR2_X1 i_1_737_3689 (.A1(\out_as[4] [6]), .A2(n_1_737_494), .ZN(n_1_737_3273));
   OAI21_X1 i_1_737_3690 (.A(n_1_737_5625), .B1(n_1_737_5624), .B2(n_1_737_4250), 
      .ZN(n_1_737_3274));
   NOR3_X1 i_1_737_3691 (.A1(\out_as[6] [6]), .A2(n_1_737_489), .A3(n_1_737_3275), 
      .ZN(n_416));
   OAI21_X1 i_1_737_3692 (.A(n_1_737_3275), .B1(\out_as[6] [6]), .B2(n_1_737_489), 
      .ZN(n_417));
   OAI21_X1 i_1_737_3693 (.A(n_1_737_3328), .B1(\out_bs[6] [6]), .B2(
      n_1_737_4514), .ZN(n_1_737_3275));
   NOR3_X1 i_1_737_3694 (.A1(\out_as[5] [6]), .A2(n_1_737_488), .A3(n_1_737_3276), 
      .ZN(n_418));
   OAI21_X1 i_1_737_3695 (.A(n_1_737_3276), .B1(\out_as[5] [6]), .B2(n_1_737_488), 
      .ZN(n_419));
   AOI21_X1 i_1_737_3696 (.A(n_844), .B1(n_845), .B2(n_1_737_4255), .ZN(
      n_1_737_3276));
   NAND3_X1 i_1_737_3697 (.A1(n_1_737_3292), .A2(n_1_737_3283), .A3(n_1_737_3277), 
      .ZN(n_420));
   AND4_X1 i_1_737_3698 (.A1(n_1_737_3289), .A2(n_1_737_3288), .A3(n_1_737_3296), 
      .A4(n_1_737_3279), .ZN(n_1_737_3277));
   INV_X1 i_1_737_3699 (.A(n_1_737_3279), .ZN(n_1_737_3278));
   OAI21_X1 i_1_737_3700 (.A(n_1_737_3280), .B1(n_1_737_5297), .B2(n_1_737_3282), 
      .ZN(n_1_737_3279));
   INV_X1 i_1_737_3701 (.A(n_1_737_3281), .ZN(n_1_737_3280));
   AOI221_X1 i_1_737_3702 (.A(\out_bs[1] [6]), .B1(\out_bs[1] [5]), .B2(
      n_1_737_4273), .C1(n_1_737_5297), .C2(n_1_737_3282), .ZN(n_1_737_3281));
   NOR2_X1 i_1_737_3703 (.A1(\out_as[1] [6]), .A2(n_1_737_484), .ZN(n_1_737_3282));
   AOI22_X1 i_1_737_3704 (.A1(n_1_737_3287), .A2(n_1_737_3285), .B1(n_1_737_5189), 
      .B2(n_1_737_3284), .ZN(n_1_737_3283));
   OAI21_X1 i_1_737_3705 (.A(n_1_737_3286), .B1(\out_as[3] [6]), .B2(n_1_737_486), 
      .ZN(n_1_737_3284));
   INV_X1 i_1_737_3706 (.A(n_1_737_3286), .ZN(n_1_737_3285));
   AOI21_X1 i_1_737_3707 (.A(\out_bs[3] [6]), .B1(\out_bs[3] [5]), .B2(
      n_1_737_4263), .ZN(n_1_737_3286));
   NOR2_X1 i_1_737_3708 (.A1(\out_as[3] [6]), .A2(n_1_737_486), .ZN(n_1_737_3287));
   NAND2_X1 i_1_737_3709 (.A1(n_1_737_5336), .A2(n_1_737_3290), .ZN(n_1_737_3288));
   OAI21_X1 i_1_737_3710 (.A(n_1_737_3291), .B1(n_1_737_5336), .B2(n_1_737_3290), 
      .ZN(n_1_737_3289));
   NOR2_X1 i_1_737_3711 (.A1(\out_as[0] [6]), .A2(n_1_737_483), .ZN(n_1_737_3290));
   OAI21_X1 i_1_737_3712 (.A(n_1_737_5671), .B1(n_1_737_4822), .B2(n_1_737_3768), 
      .ZN(n_1_737_3291));
   OAI21_X1 i_1_737_3713 (.A(n_1_737_3293), .B1(n_1_737_5235), .B2(n_1_737_3294), 
      .ZN(n_1_737_3292));
   OAI22_X1 i_1_737_3714 (.A1(\out_as[2] [6]), .A2(n_1_737_485), .B1(
      n_1_737_5236), .B2(n_1_737_3295), .ZN(n_1_737_3293));
   INV_X1 i_1_737_3715 (.A(n_1_737_3295), .ZN(n_1_737_3294));
   AOI21_X1 i_1_737_3716 (.A(\out_bs[2] [6]), .B1(\out_bs[2] [5]), .B2(
      n_1_737_4278), .ZN(n_1_737_3295));
   OAI21_X1 i_1_737_3717 (.A(n_1_737_3297), .B1(n_1_737_5365), .B2(n_1_737_3298), 
      .ZN(n_1_737_3296));
   OAI22_X1 i_1_737_3718 (.A1(\out_as[4] [6]), .A2(n_1_737_487), .B1(
      n_1_737_5366), .B2(n_1_737_3299), .ZN(n_1_737_3297));
   INV_X1 i_1_737_3719 (.A(n_1_737_3299), .ZN(n_1_737_3298));
   AOI21_X1 i_1_737_3720 (.A(\out_bs[4] [6]), .B1(\out_bs[4] [5]), .B2(
      n_1_737_4285), .ZN(n_1_737_3299));
   NOR3_X1 i_1_737_3721 (.A1(\out_as[6] [6]), .A2(n_1_737_482), .A3(n_1_737_3300), 
      .ZN(n_421));
   OAI21_X1 i_1_737_3722 (.A(n_1_737_3300), .B1(\out_as[6] [6]), .B2(n_1_737_482), 
      .ZN(n_422));
   OAI21_X1 i_1_737_3723 (.A(n_1_737_3328), .B1(\out_bs[6] [6]), .B2(
      n_1_737_4015), .ZN(n_1_737_3300));
   NOR3_X1 i_1_737_3724 (.A1(\out_as[5] [6]), .A2(n_1_737_481), .A3(n_1_737_3301), 
      .ZN(n_423));
   OAI21_X1 i_1_737_3725 (.A(n_1_737_3301), .B1(\out_as[5] [6]), .B2(n_1_737_481), 
      .ZN(n_424));
   AOI21_X1 i_1_737_3726 (.A(n_844), .B1(n_1_737_4810), .B2(n_1_737_3757), 
      .ZN(n_1_737_3301));
   OR3_X1 i_1_737_3727 (.A1(n_1_737_3318), .A2(n_1_737_3307), .A3(n_1_737_3302), 
      .ZN(n_425));
   OAI211_X1 i_1_737_3728 (.A(n_1_737_3323), .B(n_1_737_3313), .C1(n_1_737_3304), 
      .C2(n_1_737_3303), .ZN(n_1_737_3302));
   NOR2_X1 i_1_737_3729 (.A1(n_1_737_3306), .A2(n_1_737_3305), .ZN(n_1_737_3303));
   AOI21_X1 i_1_737_3730 (.A(n_1_737_5336), .B1(n_1_737_3306), .B2(n_1_737_3305), 
      .ZN(n_1_737_3304));
   NOR2_X1 i_1_737_3731 (.A1(\out_as[0] [6]), .A2(n_1_737_476), .ZN(n_1_737_3305));
   OAI21_X1 i_1_737_3732 (.A(n_1_737_5671), .B1(n_1_737_4820), .B2(n_1_737_3768), 
      .ZN(n_1_737_3306));
   INV_X1 i_1_737_3733 (.A(n_1_737_3308), .ZN(n_1_737_3307));
   OAI21_X1 i_1_737_3734 (.A(n_1_737_3309), .B1(n_1_737_5189), .B2(n_1_737_3310), 
      .ZN(n_1_737_3308));
   OAI22_X1 i_1_737_3735 (.A1(\out_as[3] [6]), .A2(n_1_737_479), .B1(
      n_1_737_5190), .B2(n_1_737_3311), .ZN(n_1_737_3309));
   INV_X1 i_1_737_3736 (.A(n_1_737_3311), .ZN(n_1_737_3310));
   AOI21_X1 i_1_737_3737 (.A(\out_bs[3] [6]), .B1(\out_bs[3] [5]), .B2(
      n_1_737_4308), .ZN(n_1_737_3311));
   INV_X1 i_1_737_3738 (.A(n_1_737_3313), .ZN(n_1_737_3312));
   AOI21_X1 i_1_737_3739 (.A(n_1_737_3314), .B1(n_1_737_5297), .B2(n_1_737_3316), 
      .ZN(n_1_737_3313));
   AOI21_X1 i_1_737_3740 (.A(n_1_737_3317), .B1(n_1_737_5298), .B2(n_1_737_3315), 
      .ZN(n_1_737_3314));
   INV_X1 i_1_737_3741 (.A(n_1_737_3316), .ZN(n_1_737_3315));
   NOR2_X1 i_1_737_3742 (.A1(\out_as[1] [6]), .A2(n_1_737_477), .ZN(n_1_737_3316));
   AOI21_X1 i_1_737_3743 (.A(\out_bs[1] [6]), .B1(\out_bs[1] [5]), .B2(
      n_1_737_4303), .ZN(n_1_737_3317));
   OAI22_X1 i_1_737_3744 (.A1(n_1_737_3322), .A2(n_1_737_3319), .B1(n_1_737_5236), 
      .B2(n_1_737_3320), .ZN(n_1_737_3318));
   NOR2_X1 i_1_737_3745 (.A1(n_1_737_5235), .A2(n_1_737_3321), .ZN(n_1_737_3319));
   INV_X1 i_1_737_3746 (.A(n_1_737_3321), .ZN(n_1_737_3320));
   NOR2_X1 i_1_737_3747 (.A1(\out_as[2] [6]), .A2(n_1_737_478), .ZN(n_1_737_3321));
   AOI21_X1 i_1_737_3748 (.A(\out_bs[2] [6]), .B1(\out_bs[2] [5]), .B2(
      n_1_737_4297), .ZN(n_1_737_3322));
   AOI21_X1 i_1_737_3749 (.A(n_1_737_3324), .B1(n_1_737_5365), .B2(n_1_737_3326), 
      .ZN(n_1_737_3323));
   AOI21_X1 i_1_737_3750 (.A(n_1_737_3327), .B1(n_1_737_5366), .B2(n_1_737_3325), 
      .ZN(n_1_737_3324));
   INV_X1 i_1_737_3751 (.A(n_1_737_3326), .ZN(n_1_737_3325));
   NOR2_X1 i_1_737_3752 (.A1(\out_as[4] [6]), .A2(n_1_737_480), .ZN(n_1_737_3326));
   AOI21_X1 i_1_737_3753 (.A(\out_bs[4] [6]), .B1(\out_bs[4] [5]), .B2(
      n_1_737_4314), .ZN(n_1_737_3327));
   NOR3_X1 i_1_737_3754 (.A1(\out_as[6] [6]), .A2(n_1_737_475), .A3(n_1_737_3329), 
      .ZN(n_426));
   OAI21_X1 i_1_737_3755 (.A(n_1_737_3329), .B1(\out_as[6] [6]), .B2(n_1_737_475), 
      .ZN(n_427));
   INV_X1 i_1_737_3756 (.A(n_1_737_3329), .ZN(n_1_737_3328));
   NOR2_X1 i_1_737_3757 (.A1(\out_bs[6] [6]), .A2(n_1_737_3330), .ZN(
      n_1_737_3329));
   NOR2_X1 i_1_737_3758 (.A1(n_1_737_5606), .A2(n_1_737_3331), .ZN(n_1_737_3330));
   INV_X1 i_1_737_3759 (.A(n_1_737_3332), .ZN(n_1_737_3331));
   NOR2_X1 i_1_737_3760 (.A1(n_1_737_5605), .A2(n_1_737_5604), .ZN(n_1_737_3332));
   NOR3_X1 i_1_737_3761 (.A1(\out_as[5] [6]), .A2(n_1_737_474), .A3(n_1_737_3419), 
      .ZN(n_428));
   OAI21_X1 i_1_737_3762 (.A(n_1_737_3419), .B1(\out_as[5] [6]), .B2(n_1_737_474), 
      .ZN(n_429));
   NAND4_X1 i_1_737_3763 (.A1(n_1_737_3343), .A2(n_1_737_3338), .A3(n_1_737_3335), 
      .A4(n_1_737_3333), .ZN(n_430));
   AOI211_X1 i_1_737_3764 (.A(n_1_737_3334), .B(n_1_737_3346), .C1(n_1_737_5336), 
      .C2(n_1_737_3342), .ZN(n_1_737_3333));
   AOI21_X1 i_1_737_3765 (.A(n_1_737_3426), .B1(n_1_737_5337), .B2(n_1_737_3341), 
      .ZN(n_1_737_3334));
   AOI22_X1 i_1_737_3766 (.A1(n_1_737_3432), .A2(n_1_737_3337), .B1(n_1_737_5189), 
      .B2(n_1_737_3336), .ZN(n_1_737_3335));
   OR2_X1 i_1_737_3767 (.A1(n_1_737_3432), .A2(n_1_737_3337), .ZN(n_1_737_3336));
   NOR2_X1 i_1_737_3768 (.A1(\out_as[3] [6]), .A2(n_1_737_472), .ZN(n_1_737_3337));
   AOI22_X1 i_1_737_3769 (.A1(n_1_737_3452), .A2(n_1_737_3340), .B1(n_1_737_5365), 
      .B2(n_1_737_3339), .ZN(n_1_737_3338));
   OAI21_X1 i_1_737_3770 (.A(n_1_737_3453), .B1(\out_as[4] [6]), .B2(n_1_737_473), 
      .ZN(n_1_737_3339));
   NOR2_X1 i_1_737_3771 (.A1(\out_as[4] [6]), .A2(n_1_737_473), .ZN(n_1_737_3340));
   INV_X1 i_1_737_3772 (.A(n_1_737_3342), .ZN(n_1_737_3341));
   NOR2_X1 i_1_737_3773 (.A1(\out_as[0] [6]), .A2(n_1_737_469), .ZN(n_1_737_3342));
   AOI22_X1 i_1_737_3774 (.A1(n_1_737_3446), .A2(n_1_737_3345), .B1(n_1_737_5235), 
      .B2(n_1_737_3344), .ZN(n_1_737_3343));
   OR2_X1 i_1_737_3775 (.A1(n_1_737_3446), .A2(n_1_737_3345), .ZN(n_1_737_3344));
   NOR2_X1 i_1_737_3776 (.A1(\out_as[2] [6]), .A2(n_1_737_471), .ZN(n_1_737_3345));
   INV_X1 i_1_737_3777 (.A(n_1_737_3347), .ZN(n_1_737_3346));
   OAI21_X1 i_1_737_3778 (.A(n_1_737_3348), .B1(n_1_737_5297), .B2(n_1_737_3350), 
      .ZN(n_1_737_3347));
   OAI21_X1 i_1_737_3779 (.A(n_1_737_3439), .B1(n_1_737_5298), .B2(n_1_737_3349), 
      .ZN(n_1_737_3348));
   INV_X1 i_1_737_3780 (.A(n_1_737_3350), .ZN(n_1_737_3349));
   NOR2_X1 i_1_737_3781 (.A1(\out_as[1] [6]), .A2(n_1_737_470), .ZN(n_1_737_3350));
   NOR2_X1 i_1_737_3782 (.A1(\out_as[6] [6]), .A2(n_1_737_468), .ZN(n_431));
   NOR3_X1 i_1_737_3783 (.A1(\out_as[5] [6]), .A2(n_1_737_467), .A3(n_1_737_3351), 
      .ZN(n_432));
   OAI21_X1 i_1_737_3784 (.A(n_1_737_3351), .B1(\out_as[5] [6]), .B2(n_1_737_467), 
      .ZN(n_433));
   AOI21_X1 i_1_737_3785 (.A(n_1_737_3420), .B1(n_1_737_4883), .B2(n_1_737_3757), 
      .ZN(n_1_737_3351));
   OR4_X1 i_1_737_3786 (.A1(n_1_737_3370), .A2(n_1_737_3365), .A3(n_1_737_3352), 
      .A4(n_1_737_3377), .ZN(n_434));
   OAI211_X1 i_1_737_3787 (.A(n_1_737_3353), .B(n_1_737_3359), .C1(n_1_737_5337), 
      .C2(n_1_737_3354), .ZN(n_1_737_3352));
   OAI22_X1 i_1_737_3788 (.A1(\out_bs[0] [6]), .A2(n_1_737_3356), .B1(
      n_1_737_5336), .B2(n_1_737_3355), .ZN(n_1_737_3353));
   INV_X1 i_1_737_3789 (.A(n_1_737_3355), .ZN(n_1_737_3354));
   NOR2_X1 i_1_737_3790 (.A1(\out_as[0] [6]), .A2(n_1_737_462), .ZN(n_1_737_3355));
   INV_X1 i_1_737_3791 (.A(n_1_737_3357), .ZN(n_1_737_3356));
   OR2_X1 i_1_737_3792 (.A1(n_1_737_5670), .A2(n_1_737_4340), .ZN(n_1_737_3357));
   INV_X1 i_1_737_3793 (.A(n_1_737_3359), .ZN(n_1_737_3358));
   OAI21_X1 i_1_737_3794 (.A(n_1_737_3360), .B1(n_1_737_5189), .B2(n_1_737_3362), 
      .ZN(n_1_737_3359));
   OAI22_X1 i_1_737_3795 (.A1(\out_as[3] [6]), .A2(n_1_737_465), .B1(
      n_1_737_5190), .B2(n_1_737_3361), .ZN(n_1_737_3360));
   INV_X1 i_1_737_3796 (.A(n_1_737_3362), .ZN(n_1_737_3361));
   NAND2_X1 i_1_737_3797 (.A1(n_1_737_5638), .A2(n_1_737_3363), .ZN(n_1_737_3362));
   OR2_X1 i_1_737_3798 (.A1(n_1_737_5637), .A2(n_1_737_4347), .ZN(n_1_737_3363));
   INV_X1 i_1_737_3799 (.A(n_1_737_3365), .ZN(n_1_737_3364));
   OAI21_X1 i_1_737_3800 (.A(n_1_737_3366), .B1(n_1_737_5298), .B2(n_1_737_3367), 
      .ZN(n_1_737_3365));
   OAI21_X1 i_1_737_3801 (.A(n_1_737_3369), .B1(n_1_737_5297), .B2(n_1_737_3368), 
      .ZN(n_1_737_3366));
   INV_X1 i_1_737_3802 (.A(n_1_737_3368), .ZN(n_1_737_3367));
   NOR2_X1 i_1_737_3803 (.A1(\out_as[1] [6]), .A2(n_1_737_463), .ZN(n_1_737_3368));
   OAI21_X1 i_1_737_3804 (.A(n_1_737_3439), .B1(n_1_737_4889), .B2(n_1_737_3788), 
      .ZN(n_1_737_3369));
   OAI21_X1 i_1_737_3805 (.A(n_1_737_3371), .B1(n_1_737_5236), .B2(n_1_737_3372), 
      .ZN(n_1_737_3370));
   OAI22_X1 i_1_737_3806 (.A1(\out_bs[2] [6]), .A2(n_1_737_3375), .B1(
      n_1_737_5235), .B2(n_1_737_3373), .ZN(n_1_737_3371));
   INV_X1 i_1_737_3807 (.A(n_1_737_3373), .ZN(n_1_737_3372));
   NOR2_X1 i_1_737_3808 (.A1(\out_as[2] [6]), .A2(n_1_737_464), .ZN(n_1_737_3373));
   INV_X1 i_1_737_3809 (.A(n_1_737_3375), .ZN(n_1_737_3374));
   NOR2_X1 i_1_737_3810 (.A1(n_1_737_5650), .A2(n_1_737_4360), .ZN(n_1_737_3375));
   INV_X1 i_1_737_3811 (.A(n_1_737_3377), .ZN(n_1_737_3376));
   OAI21_X1 i_1_737_3812 (.A(n_1_737_3378), .B1(n_1_737_5366), .B2(n_1_737_3379), 
      .ZN(n_1_737_3377));
   OAI22_X1 i_1_737_3813 (.A1(\out_bs[4] [6]), .A2(n_1_737_3381), .B1(
      n_1_737_5365), .B2(n_1_737_3380), .ZN(n_1_737_3378));
   INV_X1 i_1_737_3814 (.A(n_1_737_3380), .ZN(n_1_737_3379));
   NOR2_X1 i_1_737_3815 (.A1(\out_as[4] [6]), .A2(n_1_737_466), .ZN(n_1_737_3380));
   INV_X1 i_1_737_3816 (.A(n_1_737_3382), .ZN(n_1_737_3381));
   AOI21_X1 i_1_737_3817 (.A(n_1_737_3456), .B1(n_1_737_4912), .B2(n_1_737_3810), 
      .ZN(n_1_737_3382));
   NOR3_X1 i_1_737_3818 (.A1(\out_as[6] [6]), .A2(n_1_737_461), .A3(n_1_737_3383), 
      .ZN(n_435));
   OAI21_X1 i_1_737_3819 (.A(n_1_737_3383), .B1(\out_as[6] [6]), .B2(n_1_737_461), 
      .ZN(n_436));
   INV_X1 i_1_737_3820 (.A(n_1_737_3384), .ZN(n_1_737_3383));
   OAI21_X1 i_1_737_3821 (.A(n_1_737_5607), .B1(n_1_737_4920), .B2(n_1_737_3546), 
      .ZN(n_1_737_3384));
   NOR3_X1 i_1_737_3822 (.A1(\out_as[5] [6]), .A2(n_1_737_460), .A3(n_1_737_3385), 
      .ZN(n_437));
   OAI21_X1 i_1_737_3823 (.A(n_1_737_3385), .B1(\out_as[5] [6]), .B2(n_1_737_460), 
      .ZN(n_438));
   NOR2_X1 i_1_737_3824 (.A1(n_1_737_3420), .A2(n_1_737_3386), .ZN(n_1_737_3385));
   NOR2_X1 i_1_737_3825 (.A1(n_1_737_4925), .A2(n_1_737_3756), .ZN(n_1_737_3386));
   OR4_X1 i_1_737_3826 (.A1(n_1_737_3393), .A2(n_1_737_3388), .A3(n_1_737_3398), 
      .A4(n_1_737_3412), .ZN(n_439));
   INV_X1 i_1_737_3827 (.A(n_1_737_3388), .ZN(n_1_737_3387));
   OAI21_X1 i_1_737_3828 (.A(n_1_737_3389), .B1(n_1_737_5236), .B2(n_1_737_3390), 
      .ZN(n_1_737_3388));
   OAI22_X1 i_1_737_3829 (.A1(\out_bs[2] [6]), .A2(n_1_737_3392), .B1(
      n_1_737_5235), .B2(n_1_737_3391), .ZN(n_1_737_3389));
   INV_X1 i_1_737_3830 (.A(n_1_737_3391), .ZN(n_1_737_3390));
   NOR2_X1 i_1_737_3831 (.A1(\out_as[2] [6]), .A2(n_1_737_457), .ZN(n_1_737_3391));
   INV_X1 i_1_737_3832 (.A(n_1_737_5680), .ZN(n_1_737_3392));
   INV_X1 i_1_737_3833 (.A(n_1_737_3394), .ZN(n_1_737_3393));
   OAI21_X1 i_1_737_3834 (.A(n_1_737_3395), .B1(n_1_737_5189), .B2(n_1_737_3397), 
      .ZN(n_1_737_3394));
   OAI22_X1 i_1_737_3835 (.A1(\out_as[3] [6]), .A2(n_1_737_458), .B1(
      n_1_737_5190), .B2(n_1_737_3396), .ZN(n_1_737_3395));
   INV_X1 i_1_737_3836 (.A(n_1_737_3397), .ZN(n_1_737_3396));
   NAND2_X1 i_1_737_3837 (.A1(n_1_737_5638), .A2(n_1_737_5679), .ZN(n_1_737_3397));
   OAI211_X1 i_1_737_3838 (.A(n_1_737_3399), .B(n_1_737_3404), .C1(n_1_737_5337), 
      .C2(n_1_737_3400), .ZN(n_1_737_3398));
   OAI22_X1 i_1_737_3839 (.A1(\out_bs[0] [6]), .A2(n_1_737_3402), .B1(
      n_1_737_5336), .B2(n_1_737_3401), .ZN(n_1_737_3399));
   INV_X1 i_1_737_3840 (.A(n_1_737_3401), .ZN(n_1_737_3400));
   NOR2_X1 i_1_737_3841 (.A1(\out_as[0] [6]), .A2(n_1_737_455), .ZN(n_1_737_3401));
   INV_X1 i_1_737_3842 (.A(n_1_737_3403), .ZN(n_1_737_3402));
   AOI21_X1 i_1_737_3843 (.A(n_1_737_3427), .B1(\out_bs[0] [5]), .B2(
      n_1_737_4392), .ZN(n_1_737_3403));
   INV_X1 i_1_737_3844 (.A(n_1_737_3405), .ZN(n_1_737_3404));
   OAI21_X1 i_1_737_3845 (.A(n_1_737_3406), .B1(n_1_737_5298), .B2(n_1_737_3407), 
      .ZN(n_1_737_3405));
   OAI22_X1 i_1_737_3846 (.A1(\out_bs[1] [6]), .A2(n_1_737_3409), .B1(
      n_1_737_5297), .B2(n_1_737_3408), .ZN(n_1_737_3406));
   INV_X1 i_1_737_3847 (.A(n_1_737_3408), .ZN(n_1_737_3407));
   NOR2_X1 i_1_737_3848 (.A1(\out_as[1] [6]), .A2(n_1_737_456), .ZN(n_1_737_3408));
   INV_X1 i_1_737_3849 (.A(n_1_737_3410), .ZN(n_1_737_3409));
   AOI21_X1 i_1_737_3850 (.A(n_1_737_3440), .B1(n_1_737_4933), .B2(n_1_737_3789), 
      .ZN(n_1_737_3410));
   INV_X1 i_1_737_3851 (.A(n_1_737_3412), .ZN(n_1_737_3411));
   OAI21_X1 i_1_737_3852 (.A(n_1_737_3413), .B1(n_1_737_5366), .B2(n_1_737_3414), 
      .ZN(n_1_737_3412));
   OAI22_X1 i_1_737_3853 (.A1(\out_bs[4] [6]), .A2(n_1_737_3416), .B1(
      n_1_737_5365), .B2(n_1_737_3415), .ZN(n_1_737_3413));
   INV_X1 i_1_737_3854 (.A(n_1_737_3415), .ZN(n_1_737_3414));
   NOR2_X1 i_1_737_3855 (.A1(\out_as[4] [6]), .A2(n_1_737_459), .ZN(n_1_737_3415));
   INV_X1 i_1_737_3856 (.A(n_1_737_3417), .ZN(n_1_737_3416));
   AOI21_X1 i_1_737_3857 (.A(n_1_737_3456), .B1(\out_bs[4] [5]), .B2(
      n_1_737_4398), .ZN(n_1_737_3417));
   OR2_X1 i_1_737_3858 (.A1(n_1271), .A2(n_441), .ZN(n_440));
   NOR2_X1 i_1_737_3859 (.A1(\out_as[6] [6]), .A2(n_1_737_454), .ZN(n_441));
   NOR3_X1 i_1_737_3860 (.A1(\out_as[5] [6]), .A2(n_1_737_453), .A3(n_1_737_3418), 
      .ZN(n_442));
   OAI21_X1 i_1_737_3861 (.A(n_1_737_3418), .B1(\out_as[5] [6]), .B2(n_1_737_453), 
      .ZN(n_443));
   AOI21_X1 i_1_737_3862 (.A(n_1_737_3420), .B1(n_1_737_4965), .B2(n_1_737_3757), 
      .ZN(n_1_737_3418));
   INV_X1 i_1_737_3863 (.A(n_1_737_3420), .ZN(n_1_737_3419));
   OAI21_X1 i_1_737_3864 (.A(n_1_737_5612), .B1(n_1_737_5611), .B2(n_1_737_4403), 
      .ZN(n_1_737_3420));
   OR3_X1 i_1_737_3865 (.A1(n_1_737_3441), .A2(n_1_737_3428), .A3(n_1_737_3421), 
      .ZN(n_444));
   OAI211_X1 i_1_737_3866 (.A(n_1_737_3447), .B(n_1_737_3434), .C1(n_1_737_3423), 
      .C2(n_1_737_3422), .ZN(n_1_737_3421));
   NOR2_X1 i_1_737_3867 (.A1(n_1_737_3425), .A2(n_1_737_3424), .ZN(n_1_737_3422));
   AOI21_X1 i_1_737_3868 (.A(n_1_737_5336), .B1(n_1_737_3425), .B2(n_1_737_3424), 
      .ZN(n_1_737_3423));
   NOR2_X1 i_1_737_3869 (.A1(\out_as[0] [6]), .A2(n_1_737_448), .ZN(n_1_737_3424));
   OAI21_X1 i_1_737_3870 (.A(n_1_737_3426), .B1(n_1_737_4992), .B2(n_1_737_3768), 
      .ZN(n_1_737_3425));
   NOR2_X1 i_1_737_3871 (.A1(\out_bs[0] [6]), .A2(n_1_737_3427), .ZN(
      n_1_737_3426));
   NOR2_X1 i_1_737_3872 (.A1(n_1_737_5670), .A2(n_1_737_4437), .ZN(n_1_737_3427));
   AOI21_X1 i_1_737_3873 (.A(n_1_737_3429), .B1(n_1_737_5190), .B2(n_1_737_3431), 
      .ZN(n_1_737_3428));
   INV_X1 i_1_737_3874 (.A(n_1_737_3430), .ZN(n_1_737_3429));
   OAI22_X1 i_1_737_3875 (.A1(\out_as[3] [6]), .A2(n_1_737_451), .B1(
      n_1_737_5190), .B2(n_1_737_3431), .ZN(n_1_737_3430));
   AOI21_X1 i_1_737_3876 (.A(n_1_737_3432), .B1(\out_bs[3] [5]), .B2(
      n_1_737_4428), .ZN(n_1_737_3431));
   OAI21_X1 i_1_737_3877 (.A(n_1_737_5638), .B1(n_1_737_5637), .B2(n_1_737_4426), 
      .ZN(n_1_737_3432));
   INV_X1 i_1_737_3878 (.A(n_1_737_3434), .ZN(n_1_737_3433));
   AOI21_X1 i_1_737_3879 (.A(n_1_737_3435), .B1(n_1_737_5297), .B2(n_1_737_3437), 
      .ZN(n_1_737_3434));
   AOI22_X1 i_1_737_3880 (.A1(n_1_737_3439), .A2(n_1_737_3438), .B1(n_1_737_5298), 
      .B2(n_1_737_3436), .ZN(n_1_737_3435));
   INV_X1 i_1_737_3881 (.A(n_1_737_3437), .ZN(n_1_737_3436));
   NOR2_X1 i_1_737_3882 (.A1(\out_as[1] [6]), .A2(n_1_737_449), .ZN(n_1_737_3437));
   NAND2_X1 i_1_737_3883 (.A1(\out_bs[1] [5]), .A2(n_1_737_4452), .ZN(
      n_1_737_3438));
   NOR2_X1 i_1_737_3884 (.A1(\out_bs[1] [6]), .A2(n_1_737_3440), .ZN(
      n_1_737_3439));
   NOR2_X1 i_1_737_3885 (.A1(n_1_737_5663), .A2(n_1_737_4450), .ZN(n_1_737_3440));
   OAI21_X1 i_1_737_3886 (.A(n_1_737_3442), .B1(n_1_737_5236), .B2(n_1_737_3443), 
      .ZN(n_1_737_3441));
   OAI22_X1 i_1_737_3887 (.A1(\out_bs[2] [6]), .A2(n_1_737_3445), .B1(
      n_1_737_5235), .B2(n_1_737_3444), .ZN(n_1_737_3442));
   INV_X1 i_1_737_3888 (.A(n_1_737_3444), .ZN(n_1_737_3443));
   NOR2_X1 i_1_737_3889 (.A1(\out_as[2] [6]), .A2(n_1_737_450), .ZN(n_1_737_3444));
   NOR3_X1 i_1_737_3890 (.A1(n_1_737_5649), .A2(n_1_737_4985), .A3(n_1_737_5650), 
      .ZN(n_1_737_3445));
   OAI21_X1 i_1_737_3891 (.A(n_1_737_5651), .B1(n_1_737_5650), .B2(n_1_737_4415), 
      .ZN(n_1_737_3446));
   INV_X1 i_1_737_3892 (.A(n_1_737_3448), .ZN(n_1_737_3447));
   OAI21_X1 i_1_737_3893 (.A(n_1_737_3449), .B1(n_1_737_5366), .B2(n_1_737_3450), 
      .ZN(n_1_737_3448));
   OAI22_X1 i_1_737_3894 (.A1(\out_bs[4] [6]), .A2(n_1_737_3455), .B1(
      n_1_737_5365), .B2(n_1_737_3451), .ZN(n_1_737_3449));
   INV_X1 i_1_737_3895 (.A(n_1_737_3451), .ZN(n_1_737_3450));
   NOR2_X1 i_1_737_3896 (.A1(\out_as[4] [6]), .A2(n_1_737_452), .ZN(n_1_737_3451));
   INV_X1 i_1_737_3897 (.A(n_1_737_3453), .ZN(n_1_737_3452));
   NOR2_X1 i_1_737_3898 (.A1(\out_bs[4] [6]), .A2(n_1_737_3456), .ZN(
      n_1_737_3453));
   INV_X1 i_1_737_3899 (.A(n_1_737_3455), .ZN(n_1_737_3454));
   NOR3_X1 i_1_737_3900 (.A1(n_1_737_5623), .A2(n_1_737_4999), .A3(n_1_737_5624), 
      .ZN(n_1_737_3455));
   INV_X1 i_1_737_3901 (.A(n_1_737_3457), .ZN(n_1_737_3456));
   NAND2_X1 i_1_737_3902 (.A1(\out_bs[4] [5]), .A2(n_1_737_4462), .ZN(
      n_1_737_3457));
   NOR3_X1 i_1_737_3903 (.A1(\out_as[6] [6]), .A2(n_1_737_447), .A3(n_1_737_3458), 
      .ZN(n_445));
   OAI21_X1 i_1_737_3904 (.A(n_1_737_3458), .B1(\out_as[6] [6]), .B2(n_1_737_447), 
      .ZN(n_446));
   INV_X1 i_1_737_3905 (.A(n_1_737_3459), .ZN(n_1_737_3458));
   OAI21_X1 i_1_737_3906 (.A(n_1_737_5607), .B1(n_1_737_4513), .B2(n_1_737_3546), 
      .ZN(n_1_737_3459));
   NOR3_X1 i_1_737_3907 (.A1(\out_as[5] [6]), .A2(n_1_737_446), .A3(n_1_737_3460), 
      .ZN(n_447));
   OAI21_X1 i_1_737_3908 (.A(n_1_737_3460), .B1(\out_as[5] [6]), .B2(n_1_737_446), 
      .ZN(n_448));
   AOI21_X1 i_1_737_3909 (.A(n_844), .B1(n_845), .B2(n_1_737_4519), .ZN(
      n_1_737_3460));
   OAI211_X1 i_1_737_3910 (.A(n_1_737_3461), .B(n_1_737_3476), .C1(n_1_737_3474), 
      .C2(n_1_737_3473), .ZN(n_449));
   AND3_X1 i_1_737_3911 (.A1(n_1_737_3466), .A2(n_1_737_3463), .A3(n_1_737_3469), 
      .ZN(n_1_737_3461));
   INV_X1 i_1_737_3912 (.A(n_1_737_3463), .ZN(n_1_737_3462));
   OAI22_X1 i_1_737_3913 (.A1(n_1_737_3530), .A2(n_1_737_3464), .B1(n_1_737_5297), 
      .B2(n_1_737_3465), .ZN(n_1_737_3463));
   AND2_X1 i_1_737_3914 (.A1(n_1_737_5297), .A2(n_1_737_3465), .ZN(n_1_737_3464));
   NOR2_X1 i_1_737_3915 (.A1(\out_as[1] [6]), .A2(n_1_737_442), .ZN(n_1_737_3465));
   AOI22_X1 i_1_737_3916 (.A1(n_1_737_3521), .A2(n_1_737_3468), .B1(n_1_737_5189), 
      .B2(n_1_737_3467), .ZN(n_1_737_3466));
   OAI21_X1 i_1_737_3917 (.A(n_1_737_3522), .B1(\out_as[3] [6]), .B2(n_1_737_444), 
      .ZN(n_1_737_3467));
   NOR2_X1 i_1_737_3918 (.A1(\out_as[3] [6]), .A2(n_1_737_444), .ZN(n_1_737_3468));
   OAI21_X1 i_1_737_3919 (.A(n_1_737_3470), .B1(n_1_737_5235), .B2(n_1_737_3472), 
      .ZN(n_1_737_3469));
   INV_X1 i_1_737_3920 (.A(n_1_737_3471), .ZN(n_1_737_3470));
   AOI221_X1 i_1_737_3921 (.A(\out_bs[2] [6]), .B1(\out_bs[2] [5]), .B2(
      n_1_737_4554), .C1(n_1_737_5235), .C2(n_1_737_3472), .ZN(n_1_737_3471));
   NOR2_X1 i_1_737_3922 (.A1(\out_as[2] [6]), .A2(n_1_737_443), .ZN(n_1_737_3472));
   NOR2_X1 i_1_737_3923 (.A1(n_1_737_3514), .A2(n_1_737_3475), .ZN(n_1_737_3473));
   AOI21_X1 i_1_737_3924 (.A(n_1_737_5336), .B1(n_1_737_3514), .B2(n_1_737_3475), 
      .ZN(n_1_737_3474));
   NOR2_X1 i_1_737_3925 (.A1(\out_as[0] [6]), .A2(n_1_737_441), .ZN(n_1_737_3475));
   OAI21_X1 i_1_737_3926 (.A(n_1_737_3477), .B1(n_1_737_5365), .B2(n_1_737_3479), 
      .ZN(n_1_737_3476));
   INV_X1 i_1_737_3927 (.A(n_1_737_3478), .ZN(n_1_737_3477));
   AOI221_X1 i_1_737_3928 (.A(\out_bs[4] [6]), .B1(\out_bs[4] [5]), .B2(
      n_1_737_4564), .C1(n_1_737_5365), .C2(n_1_737_3479), .ZN(n_1_737_3478));
   NOR2_X1 i_1_737_3929 (.A1(\out_as[4] [6]), .A2(n_1_737_445), .ZN(n_1_737_3479));
   NOR3_X1 i_1_737_3930 (.A1(\out_as[6] [6]), .A2(n_1_737_440), .A3(n_1_737_3480), 
      .ZN(n_450));
   OAI21_X1 i_1_737_3931 (.A(n_1_737_3480), .B1(\out_as[6] [6]), .B2(n_1_737_440), 
      .ZN(n_451));
   INV_X1 i_1_737_3932 (.A(n_1_737_3481), .ZN(n_1_737_3480));
   OAI21_X1 i_1_737_3933 (.A(n_1_737_5607), .B1(n_1_737_3941), .B2(n_1_737_3546), 
      .ZN(n_1_737_3481));
   NOR3_X1 i_1_737_3934 (.A1(\out_as[5] [6]), .A2(n_1_737_439), .A3(n_1_737_3482), 
      .ZN(n_452));
   OAI21_X1 i_1_737_3935 (.A(n_1_737_3482), .B1(\out_as[5] [6]), .B2(n_1_737_439), 
      .ZN(n_453));
   AOI21_X1 i_1_737_3936 (.A(n_844), .B1(n_1_737_5020), .B2(n_1_737_3757), 
      .ZN(n_1_737_3482));
   NAND3_X1 i_1_737_3937 (.A1(n_1_737_3499), .A2(n_1_737_3485), .A3(n_1_737_3483), 
      .ZN(n_454));
   AND4_X1 i_1_737_3938 (.A1(n_1_737_3505), .A2(n_1_737_3503), .A3(n_1_737_3495), 
      .A4(n_1_737_3490), .ZN(n_1_737_3483));
   INV_X1 i_1_737_3939 (.A(n_1_737_3485), .ZN(n_1_737_3484));
   AOI21_X1 i_1_737_3940 (.A(n_1_737_3486), .B1(n_1_737_5297), .B2(n_1_737_3488), 
      .ZN(n_1_737_3485));
   AOI21_X1 i_1_737_3941 (.A(n_1_737_3489), .B1(n_1_737_5298), .B2(n_1_737_3487), 
      .ZN(n_1_737_3486));
   INV_X1 i_1_737_3942 (.A(n_1_737_3488), .ZN(n_1_737_3487));
   NOR2_X1 i_1_737_3943 (.A1(\out_as[1] [6]), .A2(n_1_737_435), .ZN(n_1_737_3488));
   AOI21_X1 i_1_737_3944 (.A(\out_bs[1] [6]), .B1(\out_bs[1] [5]), .B2(
      n_1_737_4498), .ZN(n_1_737_3489));
   AOI22_X1 i_1_737_3945 (.A1(n_1_737_3494), .A2(n_1_737_3492), .B1(n_1_737_5189), 
      .B2(n_1_737_3491), .ZN(n_1_737_3490));
   OAI21_X1 i_1_737_3946 (.A(n_1_737_3493), .B1(\out_as[3] [6]), .B2(n_1_737_437), 
      .ZN(n_1_737_3491));
   INV_X1 i_1_737_3947 (.A(n_1_737_3493), .ZN(n_1_737_3492));
   AOI21_X1 i_1_737_3948 (.A(\out_bs[3] [6]), .B1(\out_bs[3] [5]), .B2(
      n_1_737_4491), .ZN(n_1_737_3493));
   NOR2_X1 i_1_737_3949 (.A1(\out_as[3] [6]), .A2(n_1_737_437), .ZN(n_1_737_3494));
   OAI21_X1 i_1_737_3950 (.A(n_1_737_3496), .B1(n_1_737_5235), .B2(n_1_737_3497), 
      .ZN(n_1_737_3495));
   OAI22_X1 i_1_737_3951 (.A1(\out_as[2] [6]), .A2(n_1_737_436), .B1(
      n_1_737_5236), .B2(n_1_737_3498), .ZN(n_1_737_3496));
   INV_X1 i_1_737_3952 (.A(n_1_737_3498), .ZN(n_1_737_3497));
   AOI21_X1 i_1_737_3953 (.A(\out_bs[2] [6]), .B1(\out_bs[2] [5]), .B2(
      n_1_737_4504), .ZN(n_1_737_3498));
   OAI21_X1 i_1_737_3954 (.A(n_1_737_3500), .B1(n_1_737_5365), .B2(n_1_737_3501), 
      .ZN(n_1_737_3499));
   OAI22_X1 i_1_737_3955 (.A1(\out_as[4] [6]), .A2(n_1_737_438), .B1(
      n_1_737_5366), .B2(n_1_737_3502), .ZN(n_1_737_3500));
   INV_X1 i_1_737_3956 (.A(n_1_737_3502), .ZN(n_1_737_3501));
   AOI21_X1 i_1_737_3957 (.A(\out_bs[4] [6]), .B1(\out_bs[4] [5]), .B2(
      n_1_737_4510), .ZN(n_1_737_3502));
   OAI21_X1 i_1_737_3958 (.A(n_1_737_3504), .B1(n_1_737_5336), .B2(n_1_737_3506), 
      .ZN(n_1_737_3503));
   OAI21_X1 i_1_737_3959 (.A(n_1_737_5671), .B1(n_1_737_5028), .B2(n_1_737_3768), 
      .ZN(n_1_737_3504));
   NAND2_X1 i_1_737_3960 (.A1(n_1_737_5336), .A2(n_1_737_3506), .ZN(n_1_737_3505));
   NOR2_X1 i_1_737_3961 (.A1(\out_as[0] [6]), .A2(n_1_737_434), .ZN(n_1_737_3506));
   NOR3_X1 i_1_737_3962 (.A1(\out_as[6] [6]), .A2(n_1_737_433), .A3(n_1_737_3507), 
      .ZN(n_455));
   OAI21_X1 i_1_737_3963 (.A(n_1_737_3507), .B1(\out_as[6] [6]), .B2(n_1_737_433), 
      .ZN(n_456));
   AOI21_X1 i_1_737_3964 (.A(\out_bs[6] [6]), .B1(\out_bs[6] [5]), .B2(
      n_1_737_4512), .ZN(n_1_737_3507));
   NOR3_X1 i_1_737_3965 (.A1(\out_as[5] [6]), .A2(n_1_737_432), .A3(n_1_737_3508), 
      .ZN(n_457));
   OAI21_X1 i_1_737_3966 (.A(n_1_737_3508), .B1(\out_as[5] [6]), .B2(n_1_737_432), 
      .ZN(n_458));
   AOI21_X1 i_1_737_3967 (.A(n_844), .B1(n_845), .B2(n_1_737_4516), .ZN(
      n_1_737_3508));
   NAND4_X1 i_1_737_3968 (.A1(n_1_737_3537), .A2(n_1_737_3523), .A3(n_1_737_3515), 
      .A4(n_1_737_3509), .ZN(n_459));
   AOI211_X1 i_1_737_3969 (.A(n_1_737_3510), .B(n_1_737_3531), .C1(n_1_737_5336), 
      .C2(n_1_737_3512), .ZN(n_1_737_3509));
   INV_X1 i_1_737_3970 (.A(n_1_737_3511), .ZN(n_1_737_3510));
   OAI22_X1 i_1_737_3971 (.A1(\out_bs[0] [6]), .A2(n_1_737_3513), .B1(
      n_1_737_5336), .B2(n_1_737_3512), .ZN(n_1_737_3511));
   NOR2_X1 i_1_737_3972 (.A1(\out_as[0] [6]), .A2(n_1_737_427), .ZN(n_1_737_3512));
   NOR2_X1 i_1_737_3973 (.A1(n_1_737_5670), .A2(n_1_737_4542), .ZN(n_1_737_3513));
   OAI21_X1 i_1_737_3974 (.A(n_1_737_5671), .B1(n_1_737_5329), .B2(n_1_737_3768), 
      .ZN(n_1_737_3514));
   OAI21_X1 i_1_737_3975 (.A(n_1_737_3516), .B1(n_1_737_5189), .B2(n_1_737_3517), 
      .ZN(n_1_737_3515));
   OAI22_X1 i_1_737_3976 (.A1(\out_as[3] [6]), .A2(n_1_737_430), .B1(
      n_1_737_5190), .B2(n_1_737_3518), .ZN(n_1_737_3516));
   INV_X1 i_1_737_3977 (.A(n_1_737_3518), .ZN(n_1_737_3517));
   NOR2_X1 i_1_737_3978 (.A1(\out_bs[3] [6]), .A2(n_1_737_3520), .ZN(
      n_1_737_3518));
   INV_X1 i_1_737_3979 (.A(n_1_737_3520), .ZN(n_1_737_3519));
   NOR2_X1 i_1_737_3980 (.A1(n_1_737_5637), .A2(n_1_737_4532), .ZN(n_1_737_3520));
   INV_X1 i_1_737_3981 (.A(n_1_737_3522), .ZN(n_1_737_3521));
   AOI21_X1 i_1_737_3982 (.A(\out_bs[3] [6]), .B1(\out_bs[3] [5]), .B2(
      n_1_737_4535), .ZN(n_1_737_3522));
   INV_X1 i_1_737_3983 (.A(n_1_737_3524), .ZN(n_1_737_3523));
   OAI21_X1 i_1_737_3984 (.A(n_1_737_3525), .B1(n_1_737_5298), .B2(n_1_737_3526), 
      .ZN(n_1_737_3524));
   OAI22_X1 i_1_737_3985 (.A1(\out_bs[1] [6]), .A2(n_1_737_3529), .B1(
      n_1_737_5297), .B2(n_1_737_3527), .ZN(n_1_737_3525));
   INV_X1 i_1_737_3986 (.A(n_1_737_3527), .ZN(n_1_737_3526));
   NOR2_X1 i_1_737_3987 (.A1(\out_as[1] [6]), .A2(n_1_737_428), .ZN(n_1_737_3527));
   INV_X1 i_1_737_3988 (.A(n_1_737_3529), .ZN(n_1_737_3528));
   NOR2_X1 i_1_737_3989 (.A1(n_1_737_5663), .A2(n_1_737_4527), .ZN(n_1_737_3529));
   OAI21_X1 i_1_737_3990 (.A(n_1_737_5664), .B1(n_1_737_5663), .B2(n_1_737_4528), 
      .ZN(n_1_737_3530));
   OAI21_X1 i_1_737_3991 (.A(n_1_737_3532), .B1(n_1_737_5236), .B2(n_1_737_3533), 
      .ZN(n_1_737_3531));
   OAI22_X1 i_1_737_3992 (.A1(\out_bs[2] [6]), .A2(n_1_737_3536), .B1(
      n_1_737_5235), .B2(n_1_737_3534), .ZN(n_1_737_3532));
   INV_X1 i_1_737_3993 (.A(n_1_737_3534), .ZN(n_1_737_3533));
   NOR2_X1 i_1_737_3994 (.A1(\out_as[2] [6]), .A2(n_1_737_429), .ZN(n_1_737_3534));
   INV_X1 i_1_737_3995 (.A(n_1_737_3536), .ZN(n_1_737_3535));
   NOR2_X1 i_1_737_3996 (.A1(n_1_737_5650), .A2(n_1_737_4551), .ZN(n_1_737_3536));
   INV_X1 i_1_737_3997 (.A(n_1_737_3538), .ZN(n_1_737_3537));
   OAI21_X1 i_1_737_3998 (.A(n_1_737_3539), .B1(n_1_737_5366), .B2(n_1_737_3540), 
      .ZN(n_1_737_3538));
   OAI22_X1 i_1_737_3999 (.A1(\out_bs[4] [6]), .A2(n_1_737_3543), .B1(
      n_1_737_5365), .B2(n_1_737_3541), .ZN(n_1_737_3539));
   INV_X1 i_1_737_4000 (.A(n_1_737_3541), .ZN(n_1_737_3540));
   NOR2_X1 i_1_737_4001 (.A1(\out_as[4] [6]), .A2(n_1_737_431), .ZN(n_1_737_3541));
   INV_X1 i_1_737_4002 (.A(n_1_737_3543), .ZN(n_1_737_3542));
   NOR2_X1 i_1_737_4003 (.A1(n_1_737_5624), .A2(n_1_737_4561), .ZN(n_1_737_3543));
   NOR3_X1 i_1_737_4004 (.A1(\out_as[6] [6]), .A2(n_1_737_426), .A3(n_1_737_3544), 
      .ZN(n_460));
   OAI21_X1 i_1_737_4005 (.A(n_1_737_3544), .B1(\out_as[6] [6]), .B2(n_1_737_426), 
      .ZN(n_461));
   INV_X1 i_1_737_4006 (.A(n_1_737_3545), .ZN(n_1_737_3544));
   OAI21_X1 i_1_737_4007 (.A(n_1_737_5607), .B1(n_1_737_4014), .B2(n_1_737_3546), 
      .ZN(n_1_737_3545));
   NAND2_X1 i_1_737_4008 (.A1(\out_bs[6] [5]), .A2(\out_bs[6] [4]), .ZN(
      n_1_737_3546));
   NOR3_X1 i_1_737_4009 (.A1(\out_as[5] [6]), .A2(n_1_737_425), .A3(n_1_737_3547), 
      .ZN(n_462));
   OAI21_X1 i_1_737_4010 (.A(n_1_737_3547), .B1(\out_as[5] [6]), .B2(n_1_737_425), 
      .ZN(n_463));
   AOI21_X1 i_1_737_4011 (.A(n_844), .B1(n_1_737_5172), .B2(n_1_737_3757), 
      .ZN(n_1_737_3547));
   NAND3_X1 i_1_737_4012 (.A1(n_1_737_3559), .A2(n_1_737_3554), .A3(n_1_737_3548), 
      .ZN(n_464));
   AND4_X1 i_1_737_4013 (.A1(n_1_737_3564), .A2(n_1_737_3563), .A3(n_1_737_3567), 
      .A4(n_1_737_3549), .ZN(n_1_737_3548));
   AOI21_X1 i_1_737_4014 (.A(n_1_737_3550), .B1(n_1_737_5297), .B2(n_1_737_3552), 
      .ZN(n_1_737_3549));
   AOI21_X1 i_1_737_4015 (.A(n_1_737_3553), .B1(n_1_737_5298), .B2(n_1_737_3551), 
      .ZN(n_1_737_3550));
   INV_X1 i_1_737_4016 (.A(n_1_737_3552), .ZN(n_1_737_3551));
   NOR2_X1 i_1_737_4017 (.A1(\out_as[1] [6]), .A2(n_1_737_421), .ZN(n_1_737_3552));
   AOI21_X1 i_1_737_4018 (.A(\out_bs[1] [6]), .B1(\out_bs[1] [5]), .B2(
      n_1_737_4583), .ZN(n_1_737_3553));
   AOI22_X1 i_1_737_4019 (.A1(n_1_737_3558), .A2(n_1_737_3556), .B1(n_1_737_5189), 
      .B2(n_1_737_3555), .ZN(n_1_737_3554));
   OAI21_X1 i_1_737_4020 (.A(n_1_737_3557), .B1(\out_as[3] [6]), .B2(n_1_737_423), 
      .ZN(n_1_737_3555));
   INV_X1 i_1_737_4021 (.A(n_1_737_3557), .ZN(n_1_737_3556));
   AOI21_X1 i_1_737_4022 (.A(\out_bs[3] [6]), .B1(\out_bs[3] [5]), .B2(
      n_1_737_4576), .ZN(n_1_737_3557));
   NOR2_X1 i_1_737_4023 (.A1(\out_as[3] [6]), .A2(n_1_737_423), .ZN(n_1_737_3558));
   OAI21_X1 i_1_737_4024 (.A(n_1_737_3560), .B1(n_1_737_5235), .B2(n_1_737_3561), 
      .ZN(n_1_737_3559));
   OAI22_X1 i_1_737_4025 (.A1(\out_as[2] [6]), .A2(n_1_737_422), .B1(
      n_1_737_5236), .B2(n_1_737_3562), .ZN(n_1_737_3560));
   INV_X1 i_1_737_4026 (.A(n_1_737_3562), .ZN(n_1_737_3561));
   AOI21_X1 i_1_737_4027 (.A(\out_bs[2] [6]), .B1(\out_bs[2] [5]), .B2(
      n_1_737_4588), .ZN(n_1_737_3562));
   NAND2_X1 i_1_737_4028 (.A1(n_1_737_5336), .A2(n_1_737_3565), .ZN(n_1_737_3563));
   OAI21_X1 i_1_737_4029 (.A(n_1_737_3566), .B1(n_1_737_5336), .B2(n_1_737_3565), 
      .ZN(n_1_737_3564));
   NOR2_X1 i_1_737_4030 (.A1(\out_as[0] [6]), .A2(n_1_737_420), .ZN(n_1_737_3565));
   OAI21_X1 i_1_737_4031 (.A(n_1_737_5671), .B1(n_1_737_5325), .B2(n_1_737_3768), 
      .ZN(n_1_737_3566));
   OAI21_X1 i_1_737_4032 (.A(n_1_737_3568), .B1(n_1_737_5365), .B2(n_1_737_3569), 
      .ZN(n_1_737_3567));
   OAI22_X1 i_1_737_4033 (.A1(\out_as[4] [6]), .A2(n_1_737_424), .B1(
      n_1_737_5366), .B2(n_1_737_3570), .ZN(n_1_737_3568));
   INV_X1 i_1_737_4034 (.A(n_1_737_3570), .ZN(n_1_737_3569));
   AOI21_X1 i_1_737_4035 (.A(\out_bs[4] [6]), .B1(\out_bs[4] [5]), .B2(
      n_1_737_4594), .ZN(n_1_737_3570));
   OR2_X1 i_1_737_4036 (.A1(n_1270), .A2(n_466), .ZN(n_465));
   NOR2_X1 i_1_737_4037 (.A1(\out_as[6] [6]), .A2(n_1_737_419), .ZN(n_466));
   NOR3_X1 i_1_737_4038 (.A1(\out_as[5] [6]), .A2(n_1_737_418), .A3(n_1_737_3754), 
      .ZN(n_467));
   OAI21_X1 i_1_737_4039 (.A(n_1_737_3754), .B1(\out_as[5] [6]), .B2(n_1_737_418), 
      .ZN(n_468));
   NAND3_X1 i_1_737_4040 (.A1(n_1_737_3583), .A2(n_1_737_3580), .A3(n_1_737_3571), 
      .ZN(n_469));
   NOR3_X1 i_1_737_4041 (.A1(n_1_737_3586), .A2(n_1_737_3576), .A3(n_1_737_3572), 
      .ZN(n_1_737_3571));
   OAI21_X1 i_1_737_4042 (.A(n_1_737_3573), .B1(n_1_737_5337), .B2(n_1_737_3574), 
      .ZN(n_1_737_3572));
   OAI21_X1 i_1_737_4043 (.A(n_1_737_3764), .B1(n_1_737_5336), .B2(n_1_737_3575), 
      .ZN(n_1_737_3573));
   INV_X1 i_1_737_4044 (.A(n_1_737_3575), .ZN(n_1_737_3574));
   NOR2_X1 i_1_737_4045 (.A1(\out_as[0] [6]), .A2(n_1_737_413), .ZN(n_1_737_3575));
   OAI21_X1 i_1_737_4046 (.A(n_1_737_3577), .B1(n_1_737_3806), .B2(n_1_737_3578), 
      .ZN(n_1_737_3576));
   OAI21_X1 i_1_737_4047 (.A(n_1_737_5365), .B1(n_1_737_3805), .B2(n_1_737_3579), 
      .ZN(n_1_737_3577));
   INV_X1 i_1_737_4048 (.A(n_1_737_3579), .ZN(n_1_737_3578));
   NOR2_X1 i_1_737_4049 (.A1(\out_as[4] [6]), .A2(n_1_737_417), .ZN(n_1_737_3579));
   AOI22_X1 i_1_737_4050 (.A1(n_1_737_3775), .A2(n_1_737_3582), .B1(n_1_737_5235), 
      .B2(n_1_737_3581), .ZN(n_1_737_3580));
   OAI21_X1 i_1_737_4051 (.A(n_1_737_3776), .B1(\out_as[2] [6]), .B2(n_1_737_415), 
      .ZN(n_1_737_3581));
   NOR2_X1 i_1_737_4052 (.A1(\out_as[2] [6]), .A2(n_1_737_415), .ZN(n_1_737_3582));
   AOI22_X1 i_1_737_4053 (.A1(n_1_737_3796), .A2(n_1_737_3585), .B1(n_1_737_5189), 
      .B2(n_1_737_3584), .ZN(n_1_737_3583));
   OAI21_X1 i_1_737_4054 (.A(n_1_737_3797), .B1(\out_as[3] [6]), .B2(n_1_737_416), 
      .ZN(n_1_737_3584));
   NOR2_X1 i_1_737_4055 (.A1(\out_as[3] [6]), .A2(n_1_737_416), .ZN(n_1_737_3585));
   INV_X1 i_1_737_4056 (.A(n_1_737_3587), .ZN(n_1_737_3586));
   OAI21_X1 i_1_737_4057 (.A(n_1_737_3588), .B1(n_1_737_5297), .B2(n_1_737_3590), 
      .ZN(n_1_737_3587));
   OAI21_X1 i_1_737_4058 (.A(n_1_737_3783), .B1(n_1_737_5298), .B2(n_1_737_3589), 
      .ZN(n_1_737_3588));
   INV_X1 i_1_737_4059 (.A(n_1_737_3590), .ZN(n_1_737_3589));
   NOR2_X1 i_1_737_4060 (.A1(\out_as[1] [6]), .A2(n_1_737_414), .ZN(n_1_737_3590));
   NOR2_X1 i_1_737_4061 (.A1(\out_as[6] [6]), .A2(n_1_737_412), .ZN(n_470));
   NOR3_X1 i_1_737_4062 (.A1(\out_as[5] [6]), .A2(n_1_737_411), .A3(n_1_737_3591), 
      .ZN(n_471));
   OAI21_X1 i_1_737_4063 (.A(n_1_737_3591), .B1(\out_as[5] [6]), .B2(n_1_737_411), 
      .ZN(n_472));
   AOI21_X1 i_1_737_4064 (.A(n_1_737_3753), .B1(n_845), .B2(n_1_737_4615), 
      .ZN(n_1_737_3591));
   OAI211_X1 i_1_737_4065 (.A(n_1_737_3592), .B(n_1_737_3612), .C1(n_1_737_3608), 
      .C2(n_1_737_3607), .ZN(n_473));
   AND3_X1 i_1_737_4066 (.A1(n_1_737_3599), .A2(n_1_737_3593), .A3(n_1_737_3603), 
      .ZN(n_1_737_3592));
   INV_X1 i_1_737_4067 (.A(n_1_737_3594), .ZN(n_1_737_3593));
   OAI21_X1 i_1_737_4068 (.A(n_1_737_3595), .B1(n_1_737_5298), .B2(n_1_737_3596), 
      .ZN(n_1_737_3594));
   OAI21_X1 i_1_737_4069 (.A(n_1_737_3598), .B1(n_1_737_5297), .B2(n_1_737_3597), 
      .ZN(n_1_737_3595));
   INV_X1 i_1_737_4070 (.A(n_1_737_3597), .ZN(n_1_737_3596));
   NOR2_X1 i_1_737_4071 (.A1(\out_as[1] [6]), .A2(n_1_737_407), .ZN(n_1_737_3597));
   OAI21_X1 i_1_737_4072 (.A(n_1_737_3783), .B1(n_1_737_5663), .B2(n_1_737_4631), 
      .ZN(n_1_737_3598));
   AOI22_X1 i_1_737_4073 (.A1(n_1_737_3602), .A2(n_1_737_3601), .B1(n_1_737_5189), 
      .B2(n_1_737_3600), .ZN(n_1_737_3599));
   OR2_X1 i_1_737_4074 (.A1(n_1_737_3602), .A2(n_1_737_3601), .ZN(n_1_737_3600));
   OAI21_X1 i_1_737_4075 (.A(n_1_737_3797), .B1(n_1_737_5637), .B2(n_1_737_4622), 
      .ZN(n_1_737_3601));
   NOR2_X1 i_1_737_4076 (.A1(\out_as[3] [6]), .A2(n_1_737_409), .ZN(n_1_737_3602));
   OAI21_X1 i_1_737_4077 (.A(n_1_737_3604), .B1(n_1_737_5235), .B2(n_1_737_3606), 
      .ZN(n_1_737_3603));
   OAI22_X1 i_1_737_4078 (.A1(\out_as[2] [6]), .A2(n_1_737_408), .B1(
      n_1_737_5236), .B2(n_1_737_3605), .ZN(n_1_737_3604));
   INV_X1 i_1_737_4079 (.A(n_1_737_3606), .ZN(n_1_737_3605));
   OAI21_X1 i_1_737_4080 (.A(n_1_737_3776), .B1(n_1_737_5650), .B2(n_1_737_4638), 
      .ZN(n_1_737_3606));
   NOR2_X1 i_1_737_4081 (.A1(n_1_737_3610), .A2(n_1_737_3609), .ZN(n_1_737_3607));
   AOI21_X1 i_1_737_4082 (.A(n_1_737_5336), .B1(n_1_737_3610), .B2(n_1_737_3609), 
      .ZN(n_1_737_3608));
   NOR2_X1 i_1_737_4083 (.A1(\out_as[0] [6]), .A2(n_1_737_406), .ZN(n_1_737_3609));
   OAI21_X1 i_1_737_4084 (.A(n_1_737_3765), .B1(n_1_737_5670), .B2(n_1_737_4626), 
      .ZN(n_1_737_3610));
   INV_X1 i_1_737_4085 (.A(n_1_737_3612), .ZN(n_1_737_3611));
   OAI21_X1 i_1_737_4086 (.A(n_1_737_3613), .B1(n_1_737_5365), .B2(n_1_737_3615), 
      .ZN(n_1_737_3612));
   OAI22_X1 i_1_737_4087 (.A1(\out_as[4] [6]), .A2(n_1_737_410), .B1(
      n_1_737_5366), .B2(n_1_737_3614), .ZN(n_1_737_3613));
   INV_X1 i_1_737_4088 (.A(n_1_737_3615), .ZN(n_1_737_3614));
   OAI21_X1 i_1_737_4089 (.A(n_1_737_3806), .B1(n_1_737_5624), .B2(n_1_737_4643), 
      .ZN(n_1_737_3615));
   NOR2_X1 i_1_737_4090 (.A1(\out_as[6] [6]), .A2(n_1_737_405), .ZN(n_474));
   NOR3_X1 i_1_737_4091 (.A1(\out_as[5] [6]), .A2(n_1_737_404), .A3(n_1_737_3616), 
      .ZN(n_475));
   OAI21_X1 i_1_737_4092 (.A(n_1_737_3616), .B1(\out_as[5] [6]), .B2(n_1_737_404), 
      .ZN(n_476));
   AOI21_X1 i_1_737_4093 (.A(n_1_737_3753), .B1(n_845), .B2(n_1_737_4646), 
      .ZN(n_1_737_3616));
   NAND3_X1 i_1_737_4094 (.A1(n_1_737_3632), .A2(n_1_737_3624), .A3(n_1_737_3617), 
      .ZN(n_477));
   AND4_X1 i_1_737_4095 (.A1(n_1_737_3629), .A2(n_1_737_3628), .A3(n_1_737_3637), 
      .A4(n_1_737_3618), .ZN(n_1_737_3617));
   INV_X1 i_1_737_4096 (.A(n_1_737_3619), .ZN(n_1_737_3618));
   OAI21_X1 i_1_737_4097 (.A(n_1_737_3620), .B1(n_1_737_5298), .B2(n_1_737_3621), 
      .ZN(n_1_737_3619));
   OAI21_X1 i_1_737_4098 (.A(n_1_737_3623), .B1(n_1_737_5297), .B2(n_1_737_3622), 
      .ZN(n_1_737_3620));
   INV_X1 i_1_737_4099 (.A(n_1_737_3622), .ZN(n_1_737_3621));
   NOR2_X1 i_1_737_4100 (.A1(\out_as[1] [6]), .A2(n_1_737_400), .ZN(n_1_737_3622));
   OAI21_X1 i_1_737_4101 (.A(n_1_737_3783), .B1(n_1_737_5663), .B2(n_1_737_4653), 
      .ZN(n_1_737_3623));
   AOI22_X1 i_1_737_4102 (.A1(n_1_737_3627), .A2(n_1_737_3626), .B1(n_1_737_5189), 
      .B2(n_1_737_3625), .ZN(n_1_737_3624));
   OR2_X1 i_1_737_4103 (.A1(n_1_737_3627), .A2(n_1_737_3626), .ZN(n_1_737_3625));
   OAI21_X1 i_1_737_4104 (.A(n_1_737_3797), .B1(n_1_737_5637), .B2(n_1_737_4658), 
      .ZN(n_1_737_3626));
   NOR2_X1 i_1_737_4105 (.A1(\out_as[3] [6]), .A2(n_1_737_402), .ZN(n_1_737_3627));
   NAND2_X1 i_1_737_4106 (.A1(n_1_737_5336), .A2(n_1_737_3630), .ZN(n_1_737_3628));
   OAI21_X1 i_1_737_4107 (.A(n_1_737_3631), .B1(n_1_737_5336), .B2(n_1_737_3630), 
      .ZN(n_1_737_3629));
   NOR2_X1 i_1_737_4108 (.A1(\out_as[0] [6]), .A2(n_1_737_399), .ZN(n_1_737_3630));
   OAI21_X1 i_1_737_4109 (.A(n_1_737_3765), .B1(n_1_737_5670), .B2(n_1_737_4669), 
      .ZN(n_1_737_3631));
   OAI21_X1 i_1_737_4110 (.A(n_1_737_3633), .B1(n_1_737_5235), .B2(n_1_737_3635), 
      .ZN(n_1_737_3632));
   OAI22_X1 i_1_737_4111 (.A1(\out_as[2] [6]), .A2(n_1_737_401), .B1(
      n_1_737_5236), .B2(n_1_737_3634), .ZN(n_1_737_3633));
   INV_X1 i_1_737_4112 (.A(n_1_737_3635), .ZN(n_1_737_3634));
   OAI21_X1 i_1_737_4113 (.A(n_1_737_3776), .B1(n_1_737_5650), .B2(n_1_737_4664), 
      .ZN(n_1_737_3635));
   INV_X1 i_1_737_4114 (.A(n_1_737_3637), .ZN(n_1_737_3636));
   OAI21_X1 i_1_737_4115 (.A(n_1_737_3638), .B1(n_1_737_5365), .B2(n_1_737_3640), 
      .ZN(n_1_737_3637));
   OAI22_X1 i_1_737_4116 (.A1(\out_as[4] [6]), .A2(n_1_737_403), .B1(
      n_1_737_5366), .B2(n_1_737_3639), .ZN(n_1_737_3638));
   INV_X1 i_1_737_4117 (.A(n_1_737_3640), .ZN(n_1_737_3639));
   OAI21_X1 i_1_737_4118 (.A(n_1_737_3806), .B1(n_1_737_5624), .B2(n_1_737_4676), 
      .ZN(n_1_737_3640));
   NOR2_X1 i_1_737_4119 (.A1(\out_as[6] [6]), .A2(n_1_737_398), .ZN(n_478));
   NOR3_X1 i_1_737_4120 (.A1(\out_as[5] [6]), .A2(n_1_737_397), .A3(n_1_737_3641), 
      .ZN(n_479));
   OAI21_X1 i_1_737_4121 (.A(n_1_737_3641), .B1(\out_as[5] [6]), .B2(n_1_737_397), 
      .ZN(n_480));
   AOI21_X1 i_1_737_4122 (.A(n_1_737_3753), .B1(n_845), .B2(n_1_737_4679), 
      .ZN(n_1_737_3641));
   OAI211_X1 i_1_737_4123 (.A(n_1_737_3657), .B(n_1_737_3642), .C1(n_1_737_3644), 
      .C2(n_1_737_3643), .ZN(n_481));
   AND3_X1 i_1_737_4124 (.A1(n_1_737_3662), .A2(n_1_737_3651), .A3(n_1_737_3647), 
      .ZN(n_1_737_3642));
   NOR2_X1 i_1_737_4125 (.A1(n_1_737_3646), .A2(n_1_737_3645), .ZN(n_1_737_3643));
   AOI21_X1 i_1_737_4126 (.A(n_1_737_5336), .B1(n_1_737_3646), .B2(n_1_737_3645), 
      .ZN(n_1_737_3644));
   NOR2_X1 i_1_737_4127 (.A1(\out_as[0] [6]), .A2(n_1_737_392), .ZN(n_1_737_3645));
   OAI21_X1 i_1_737_4128 (.A(n_1_737_5671), .B1(n_1_737_5670), .B2(n_1_737_4684), 
      .ZN(n_1_737_3646));
   OAI21_X1 i_1_737_4129 (.A(n_1_737_3648), .B1(n_1_737_5189), .B2(n_1_737_3650), 
      .ZN(n_1_737_3647));
   OAI22_X1 i_1_737_4130 (.A1(\out_as[3] [6]), .A2(n_1_737_395), .B1(
      n_1_737_5190), .B2(n_1_737_3649), .ZN(n_1_737_3648));
   INV_X1 i_1_737_4131 (.A(n_1_737_3650), .ZN(n_1_737_3649));
   OAI21_X1 i_1_737_4132 (.A(n_1_737_3797), .B1(n_1_737_5637), .B2(n_1_737_4691), 
      .ZN(n_1_737_3650));
   INV_X1 i_1_737_4133 (.A(n_1_737_3652), .ZN(n_1_737_3651));
   OAI21_X1 i_1_737_4134 (.A(n_1_737_3653), .B1(n_1_737_5298), .B2(n_1_737_3654), 
      .ZN(n_1_737_3652));
   OAI21_X1 i_1_737_4135 (.A(n_1_737_3656), .B1(n_1_737_5297), .B2(n_1_737_3655), 
      .ZN(n_1_737_3653));
   INV_X1 i_1_737_4136 (.A(n_1_737_3655), .ZN(n_1_737_3654));
   NOR2_X1 i_1_737_4137 (.A1(\out_as[1] [6]), .A2(n_1_737_393), .ZN(n_1_737_3655));
   OAI21_X1 i_1_737_4138 (.A(n_1_737_5664), .B1(n_1_737_5663), .B2(n_1_737_4697), 
      .ZN(n_1_737_3656));
   AOI21_X1 i_1_737_4139 (.A(n_1_737_3658), .B1(n_1_737_5235), .B2(n_1_737_3660), 
      .ZN(n_1_737_3657));
   INV_X1 i_1_737_4140 (.A(n_1_737_3659), .ZN(n_1_737_3658));
   OAI21_X1 i_1_737_4141 (.A(n_1_737_3661), .B1(n_1_737_5235), .B2(n_1_737_3660), 
      .ZN(n_1_737_3659));
   NOR2_X1 i_1_737_4142 (.A1(\out_as[2] [6]), .A2(n_1_737_394), .ZN(n_1_737_3660));
   OAI21_X1 i_1_737_4143 (.A(n_1_737_5651), .B1(n_1_737_5650), .B2(n_1_737_4705), 
      .ZN(n_1_737_3661));
   INV_X1 i_1_737_4144 (.A(n_1_737_3663), .ZN(n_1_737_3662));
   OAI21_X1 i_1_737_4145 (.A(n_1_737_3664), .B1(n_1_737_5366), .B2(n_1_737_3665), 
      .ZN(n_1_737_3663));
   OAI21_X1 i_1_737_4146 (.A(n_1_737_3667), .B1(n_1_737_5365), .B2(n_1_737_3666), 
      .ZN(n_1_737_3664));
   INV_X1 i_1_737_4147 (.A(n_1_737_3666), .ZN(n_1_737_3665));
   NOR2_X1 i_1_737_4148 (.A1(\out_as[4] [6]), .A2(n_1_737_396), .ZN(n_1_737_3666));
   OAI21_X1 i_1_737_4149 (.A(n_1_737_5625), .B1(n_1_737_5624), .B2(n_1_737_4713), 
      .ZN(n_1_737_3667));
   NOR3_X1 i_1_737_4150 (.A1(\out_as[6] [6]), .A2(n_1_737_391), .A3(n_1_737_3668), 
      .ZN(n_482));
   OAI21_X1 i_1_737_4151 (.A(n_1_737_3668), .B1(\out_as[6] [6]), .B2(n_1_737_391), 
      .ZN(n_483));
   AOI21_X1 i_1_737_4152 (.A(\out_bs[6] [6]), .B1(\out_bs[6] [5]), .B2(
      n_1_737_3697), .ZN(n_1_737_3668));
   NOR3_X1 i_1_737_4153 (.A1(\out_as[5] [6]), .A2(n_1_737_390), .A3(n_1_737_3669), 
      .ZN(n_484));
   OAI21_X1 i_1_737_4154 (.A(n_1_737_3669), .B1(\out_as[5] [6]), .B2(n_1_737_390), 
      .ZN(n_485));
   AOI21_X1 i_1_737_4155 (.A(n_844), .B1(n_845), .B2(n_1_737_4741), .ZN(
      n_1_737_3669));
   OAI211_X1 i_1_737_4156 (.A(n_1_737_3670), .B(n_1_737_3690), .C1(n_1_737_3686), 
      .C2(n_1_737_3685), .ZN(n_486));
   AND3_X1 i_1_737_4157 (.A1(n_1_737_3677), .A2(n_1_737_3671), .A3(n_1_737_3681), 
      .ZN(n_1_737_3670));
   INV_X1 i_1_737_4158 (.A(n_1_737_3672), .ZN(n_1_737_3671));
   OAI21_X1 i_1_737_4159 (.A(n_1_737_3673), .B1(n_1_737_5298), .B2(n_1_737_3674), 
      .ZN(n_1_737_3672));
   OAI21_X1 i_1_737_4160 (.A(n_1_737_3676), .B1(n_1_737_5297), .B2(n_1_737_3675), 
      .ZN(n_1_737_3673));
   INV_X1 i_1_737_4161 (.A(n_1_737_3675), .ZN(n_1_737_3674));
   NOR2_X1 i_1_737_4162 (.A1(\out_as[1] [6]), .A2(n_1_737_386), .ZN(n_1_737_3675));
   OAI21_X1 i_1_737_4163 (.A(n_1_737_5664), .B1(n_1_737_5663), .B2(n_1_737_4752), 
      .ZN(n_1_737_3676));
   AOI22_X1 i_1_737_4164 (.A1(n_1_737_3680), .A2(n_1_737_3679), .B1(n_1_737_5189), 
      .B2(n_1_737_3678), .ZN(n_1_737_3677));
   OR2_X1 i_1_737_4165 (.A1(n_1_737_3680), .A2(n_1_737_3679), .ZN(n_1_737_3678));
   OAI21_X1 i_1_737_4166 (.A(n_1_737_5638), .B1(n_1_737_5637), .B2(n_1_737_4762), 
      .ZN(n_1_737_3679));
   NOR2_X1 i_1_737_4167 (.A1(\out_as[3] [6]), .A2(n_1_737_388), .ZN(n_1_737_3680));
   OAI21_X1 i_1_737_4168 (.A(n_1_737_3682), .B1(n_1_737_5235), .B2(n_1_737_3684), 
      .ZN(n_1_737_3681));
   OAI22_X1 i_1_737_4169 (.A1(\out_as[2] [6]), .A2(n_1_737_387), .B1(
      n_1_737_5236), .B2(n_1_737_3683), .ZN(n_1_737_3682));
   INV_X1 i_1_737_4170 (.A(n_1_737_3684), .ZN(n_1_737_3683));
   OAI21_X1 i_1_737_4171 (.A(n_1_737_5651), .B1(n_1_737_5650), .B2(n_1_737_4771), 
      .ZN(n_1_737_3684));
   NOR2_X1 i_1_737_4172 (.A1(n_1_737_3688), .A2(n_1_737_3687), .ZN(n_1_737_3685));
   AOI21_X1 i_1_737_4173 (.A(n_1_737_5336), .B1(n_1_737_3688), .B2(n_1_737_3687), 
      .ZN(n_1_737_3686));
   NOR2_X1 i_1_737_4174 (.A1(\out_as[0] [6]), .A2(n_1_737_385), .ZN(n_1_737_3687));
   OAI21_X1 i_1_737_4175 (.A(n_1_737_5671), .B1(n_1_737_5670), .B2(n_1_737_4779), 
      .ZN(n_1_737_3688));
   INV_X1 i_1_737_4176 (.A(n_1_737_3690), .ZN(n_1_737_3689));
   OAI21_X1 i_1_737_4177 (.A(n_1_737_3691), .B1(n_1_737_5365), .B2(n_1_737_3693), 
      .ZN(n_1_737_3690));
   OAI22_X1 i_1_737_4178 (.A1(\out_as[4] [6]), .A2(n_1_737_389), .B1(
      n_1_737_5366), .B2(n_1_737_3692), .ZN(n_1_737_3691));
   INV_X1 i_1_737_4179 (.A(n_1_737_3693), .ZN(n_1_737_3692));
   OAI21_X1 i_1_737_4180 (.A(n_1_737_5625), .B1(n_1_737_5624), .B2(n_1_737_4789), 
      .ZN(n_1_737_3693));
   NOR3_X1 i_1_737_4181 (.A1(\out_as[6] [6]), .A2(n_1_737_384), .A3(n_1_737_3694), 
      .ZN(n_487));
   OAI21_X1 i_1_737_4182 (.A(n_1_737_3694), .B1(\out_as[6] [6]), .B2(n_1_737_384), 
      .ZN(n_488));
   AOI21_X1 i_1_737_4183 (.A(\out_bs[6] [6]), .B1(\out_bs[6] [5]), .B2(
      n_1_737_3695), .ZN(n_1_737_3694));
   OAI21_X1 i_1_737_4184 (.A(n_1_737_3696), .B1(n_1_737_5604), .B2(n_1_737_3943), 
      .ZN(n_1_737_3695));
   INV_X1 i_1_737_4185 (.A(n_1_737_3697), .ZN(n_1_737_3696));
   OAI21_X1 i_1_737_4186 (.A(n_1_737_5605), .B1(n_1_737_5604), .B2(n_1_737_5603), 
      .ZN(n_1_737_3697));
   NOR3_X1 i_1_737_4187 (.A1(\out_as[5] [6]), .A2(n_1_737_383), .A3(n_1_737_3698), 
      .ZN(n_489));
   OAI21_X1 i_1_737_4188 (.A(n_1_737_3698), .B1(\out_as[5] [6]), .B2(n_1_737_383), 
      .ZN(n_490));
   AOI21_X1 i_1_737_4189 (.A(n_844), .B1(n_845), .B2(n_1_737_4738), .ZN(
      n_1_737_3698));
   OR4_X1 i_1_737_4190 (.A1(n_1_737_3715), .A2(n_1_737_3710), .A3(n_1_737_3699), 
      .A4(n_1_737_3721), .ZN(n_491));
   OAI211_X1 i_1_737_4191 (.A(n_1_737_3700), .B(n_1_737_3705), .C1(n_1_737_5337), 
      .C2(n_1_737_3701), .ZN(n_1_737_3699));
   OAI21_X1 i_1_737_4192 (.A(n_1_737_3703), .B1(n_1_737_5336), .B2(n_1_737_3702), 
      .ZN(n_1_737_3700));
   INV_X1 i_1_737_4193 (.A(n_1_737_3702), .ZN(n_1_737_3701));
   NOR2_X1 i_1_737_4194 (.A1(\out_as[0] [6]), .A2(n_1_737_378), .ZN(n_1_737_3702));
   OAI21_X1 i_1_737_4195 (.A(n_1_737_5671), .B1(n_1_737_5670), .B2(n_1_737_4777), 
      .ZN(n_1_737_3703));
   INV_X1 i_1_737_4196 (.A(n_1_737_3705), .ZN(n_1_737_3704));
   OAI21_X1 i_1_737_4197 (.A(n_1_737_3706), .B1(n_1_737_5189), .B2(n_1_737_3708), 
      .ZN(n_1_737_3705));
   OAI22_X1 i_1_737_4198 (.A1(\out_as[3] [6]), .A2(n_1_737_381), .B1(
      n_1_737_5190), .B2(n_1_737_3707), .ZN(n_1_737_3706));
   INV_X1 i_1_737_4199 (.A(n_1_737_3708), .ZN(n_1_737_3707));
   OAI21_X1 i_1_737_4200 (.A(n_1_737_5638), .B1(n_1_737_5637), .B2(n_1_737_4760), 
      .ZN(n_1_737_3708));
   INV_X1 i_1_737_4201 (.A(n_1_737_3710), .ZN(n_1_737_3709));
   OAI21_X1 i_1_737_4202 (.A(n_1_737_3711), .B1(n_1_737_5298), .B2(n_1_737_3712), 
      .ZN(n_1_737_3710));
   OAI21_X1 i_1_737_4203 (.A(n_1_737_3714), .B1(n_1_737_5297), .B2(n_1_737_3713), 
      .ZN(n_1_737_3711));
   INV_X1 i_1_737_4204 (.A(n_1_737_3713), .ZN(n_1_737_3712));
   NOR2_X1 i_1_737_4205 (.A1(\out_as[1] [6]), .A2(n_1_737_379), .ZN(n_1_737_3713));
   OAI21_X1 i_1_737_4206 (.A(n_1_737_5664), .B1(n_1_737_5663), .B2(n_1_737_4750), 
      .ZN(n_1_737_3714));
   OAI21_X1 i_1_737_4207 (.A(n_1_737_3716), .B1(n_1_737_5236), .B2(n_1_737_3717), 
      .ZN(n_1_737_3715));
   OAI21_X1 i_1_737_4208 (.A(n_1_737_3719), .B1(n_1_737_5235), .B2(n_1_737_3718), 
      .ZN(n_1_737_3716));
   INV_X1 i_1_737_4209 (.A(n_1_737_3718), .ZN(n_1_737_3717));
   NOR2_X1 i_1_737_4210 (.A1(\out_as[2] [6]), .A2(n_1_737_380), .ZN(n_1_737_3718));
   OAI21_X1 i_1_737_4211 (.A(n_1_737_5651), .B1(n_1_737_5650), .B2(n_1_737_4769), 
      .ZN(n_1_737_3719));
   INV_X1 i_1_737_4212 (.A(n_1_737_3721), .ZN(n_1_737_3720));
   OAI21_X1 i_1_737_4213 (.A(n_1_737_3722), .B1(n_1_737_5366), .B2(n_1_737_3723), 
      .ZN(n_1_737_3721));
   OAI21_X1 i_1_737_4214 (.A(n_1_737_3725), .B1(n_1_737_5365), .B2(n_1_737_3724), 
      .ZN(n_1_737_3722));
   INV_X1 i_1_737_4215 (.A(n_1_737_3724), .ZN(n_1_737_3723));
   NOR2_X1 i_1_737_4216 (.A1(\out_as[4] [6]), .A2(n_1_737_382), .ZN(n_1_737_3724));
   OAI21_X1 i_1_737_4217 (.A(n_1_737_5625), .B1(n_1_737_5624), .B2(n_1_737_4787), 
      .ZN(n_1_737_3725));
   NOR3_X1 i_1_737_4218 (.A1(\out_as[6] [6]), .A2(n_1_737_377), .A3(n_1_737_3748), 
      .ZN(n_492));
   OAI21_X1 i_1_737_4219 (.A(n_1_737_3748), .B1(\out_as[6] [6]), .B2(n_1_737_377), 
      .ZN(n_493));
   NOR3_X1 i_1_737_4220 (.A1(\out_as[5] [6]), .A2(n_1_737_376), .A3(n_1_737_3752), 
      .ZN(n_494));
   OAI21_X1 i_1_737_4221 (.A(n_1_737_3752), .B1(\out_as[5] [6]), .B2(n_1_737_376), 
      .ZN(n_495));
   NAND4_X1 i_1_737_4222 (.A1(n_1_737_3738), .A2(n_1_737_3733), .A3(n_1_737_3726), 
      .A4(n_1_737_3742), .ZN(n_496));
   AND3_X1 i_1_737_4223 (.A1(n_1_737_3728), .A2(n_1_737_3727), .A3(n_1_737_3730), 
      .ZN(n_1_737_3726));
   NAND2_X1 i_1_737_4224 (.A1(n_1_737_5336), .A2(n_1_737_3729), .ZN(n_1_737_3727));
   OAI21_X1 i_1_737_4225 (.A(n_1_737_3763), .B1(n_1_737_5336), .B2(n_1_737_3729), 
      .ZN(n_1_737_3728));
   NOR2_X1 i_1_737_4226 (.A1(\out_as[0] [6]), .A2(n_1_737_371), .ZN(n_1_737_3729));
   OAI22_X1 i_1_737_4227 (.A1(n_1_737_3795), .A2(n_1_737_3731), .B1(n_1_737_5189), 
      .B2(n_1_737_3732), .ZN(n_1_737_3730));
   AND2_X1 i_1_737_4228 (.A1(n_1_737_5189), .A2(n_1_737_3732), .ZN(n_1_737_3731));
   NOR2_X1 i_1_737_4229 (.A1(\out_as[3] [6]), .A2(n_1_737_374), .ZN(n_1_737_3732));
   INV_X1 i_1_737_4230 (.A(n_1_737_3734), .ZN(n_1_737_3733));
   OAI21_X1 i_1_737_4231 (.A(n_1_737_3735), .B1(n_1_737_5298), .B2(n_1_737_3736), 
      .ZN(n_1_737_3734));
   OAI22_X1 i_1_737_4232 (.A1(\out_bs[1] [6]), .A2(n_1_737_3786), .B1(
      n_1_737_5297), .B2(n_1_737_3737), .ZN(n_1_737_3735));
   INV_X1 i_1_737_4233 (.A(n_1_737_3737), .ZN(n_1_737_3736));
   NOR2_X1 i_1_737_4234 (.A1(\out_as[1] [6]), .A2(n_1_737_372), .ZN(n_1_737_3737));
   AOI21_X1 i_1_737_4235 (.A(n_1_737_3739), .B1(n_1_737_5235), .B2(n_1_737_3741), 
      .ZN(n_1_737_3738));
   AOI22_X1 i_1_737_4236 (.A1(n_1_737_5651), .A2(n_1_737_3777), .B1(n_1_737_5236), 
      .B2(n_1_737_3740), .ZN(n_1_737_3739));
   INV_X1 i_1_737_4237 (.A(n_1_737_3741), .ZN(n_1_737_3740));
   NOR2_X1 i_1_737_4238 (.A1(\out_as[2] [6]), .A2(n_1_737_373), .ZN(n_1_737_3741));
   AOI21_X1 i_1_737_4239 (.A(n_1_737_3743), .B1(n_1_737_5365), .B2(n_1_737_3745), 
      .ZN(n_1_737_3742));
   AOI22_X1 i_1_737_4240 (.A1(n_1_737_5625), .A2(n_1_737_3809), .B1(n_1_737_5366), 
      .B2(n_1_737_3744), .ZN(n_1_737_3743));
   INV_X1 i_1_737_4241 (.A(n_1_737_3745), .ZN(n_1_737_3744));
   NOR2_X1 i_1_737_4242 (.A1(\out_as[4] [6]), .A2(n_1_737_375), .ZN(n_1_737_3745));
   NOR3_X1 i_1_737_4243 (.A1(\out_as[6] [6]), .A2(n_1_737_370), .A3(n_1_737_3746), 
      .ZN(n_497));
   OAI21_X1 i_1_737_4244 (.A(n_1_737_3746), .B1(\out_as[6] [6]), .B2(n_1_737_370), 
      .ZN(n_498));
   INV_X1 i_1_737_4245 (.A(n_1_737_3747), .ZN(n_1_737_3746));
   OAI21_X1 i_1_737_4246 (.A(n_1_737_5607), .B1(n_1_737_5606), .B2(n_1_737_3749), 
      .ZN(n_1_737_3747));
   AOI21_X1 i_1_737_4247 (.A(\out_bs[6] [6]), .B1(\out_bs[6] [5]), .B2(
      n_1_737_3750), .ZN(n_1_737_3748));
   AOI21_X1 i_1_737_4248 (.A(\out_bs[6] [4]), .B1(n_847), .B2(n_1_737_4015), 
      .ZN(n_1_737_3749));
   OAI21_X1 i_1_737_4249 (.A(n_1_737_5605), .B1(n_1_737_5604), .B2(n_1_737_4515), 
      .ZN(n_1_737_3750));
   NOR3_X1 i_1_737_4250 (.A1(\out_as[5] [6]), .A2(n_1_737_369), .A3(n_1_737_3751), 
      .ZN(n_499));
   OAI21_X1 i_1_737_4251 (.A(n_1_737_3751), .B1(\out_as[5] [6]), .B2(n_1_737_369), 
      .ZN(n_500));
   AND2_X1 i_1_737_4252 (.A1(n_1_737_5612), .A2(n_1_737_3755), .ZN(n_1_737_3751));
   AOI21_X1 i_1_737_4253 (.A(n_844), .B1(n_845), .B2(n_1_737_4812), .ZN(
      n_1_737_3752));
   INV_X1 i_1_737_4254 (.A(n_1_737_3754), .ZN(n_1_737_3753));
   NOR2_X1 i_1_737_4255 (.A1(n_844), .A2(n_1_737_3757), .ZN(n_1_737_3754));
   OAI21_X1 i_1_737_4256 (.A(n_845), .B1(n_848), .B2(n_1_737_4810), .ZN(
      n_1_737_3755));
   INV_X1 i_1_737_4257 (.A(n_1_737_3757), .ZN(n_1_737_3756));
   NOR2_X1 i_1_737_4258 (.A1(n_1_737_5611), .A2(n_1_737_5610), .ZN(n_1_737_3757));
   NAND3_X1 i_1_737_4259 (.A1(n_1_737_3790), .A2(n_1_737_3770), .A3(n_1_737_3758), 
      .ZN(n_501));
   NOR3_X1 i_1_737_4260 (.A1(n_1_737_3801), .A2(n_1_737_3779), .A3(n_1_737_3759), 
      .ZN(n_1_737_3758));
   OAI21_X1 i_1_737_4261 (.A(n_1_737_3760), .B1(n_1_737_5337), .B2(n_1_737_3761), 
      .ZN(n_1_737_3759));
   OAI22_X1 i_1_737_4262 (.A1(n_1_737_3766), .A2(n_1_737_3763), .B1(n_1_737_5336), 
      .B2(n_1_737_3762), .ZN(n_1_737_3760));
   INV_X1 i_1_737_4263 (.A(n_1_737_3762), .ZN(n_1_737_3761));
   NOR2_X1 i_1_737_4264 (.A1(\out_as[0] [6]), .A2(n_1_737_364), .ZN(n_1_737_3762));
   NAND2_X1 i_1_737_4265 (.A1(n_1_737_5671), .A2(n_1_737_3767), .ZN(n_1_737_3763));
   INV_X1 i_1_737_4266 (.A(n_1_737_3765), .ZN(n_1_737_3764));
   NOR2_X1 i_1_737_4267 (.A1(\out_bs[0] [6]), .A2(n_1_737_3769), .ZN(
      n_1_737_3765));
   AND2_X1 i_1_737_4268 (.A1(\out_bs[0] [5]), .A2(n_1_737_4824), .ZN(
      n_1_737_3766));
   OAI21_X1 i_1_737_4269 (.A(\out_bs[0] [5]), .B1(\out_bs[0] [4]), .B2(
      n_1_737_4823), .ZN(n_1_737_3767));
   INV_X1 i_1_737_4270 (.A(n_1_737_3769), .ZN(n_1_737_3768));
   NOR2_X1 i_1_737_4271 (.A1(n_1_737_5670), .A2(n_1_737_5669), .ZN(n_1_737_3769));
   AOI21_X1 i_1_737_4272 (.A(n_1_737_3771), .B1(n_1_737_5235), .B2(n_1_737_3773), 
      .ZN(n_1_737_3770));
   INV_X1 i_1_737_4273 (.A(n_1_737_3772), .ZN(n_1_737_3771));
   OAI21_X1 i_1_737_4274 (.A(n_1_737_3774), .B1(n_1_737_5235), .B2(n_1_737_3773), 
      .ZN(n_1_737_3772));
   NOR2_X1 i_1_737_4275 (.A1(\out_as[2] [6]), .A2(n_1_737_366), .ZN(n_1_737_3773));
   OAI21_X1 i_1_737_4276 (.A(n_1_737_5651), .B1(n_1_737_5650), .B2(n_1_737_4850), 
      .ZN(n_1_737_3774));
   INV_X1 i_1_737_4277 (.A(n_1_737_3776), .ZN(n_1_737_3775));
   NOR2_X1 i_1_737_4278 (.A1(\out_bs[2] [6]), .A2(n_1_737_3778), .ZN(
      n_1_737_3776));
   OAI21_X1 i_1_737_4279 (.A(\out_bs[2] [5]), .B1(\out_bs[2] [4]), .B2(
      n_1_737_4854), .ZN(n_1_737_3777));
   NOR2_X1 i_1_737_4280 (.A1(n_1_737_5650), .A2(n_1_737_5649), .ZN(n_1_737_3778));
   OAI21_X1 i_1_737_4281 (.A(n_1_737_3780), .B1(n_1_737_5298), .B2(n_1_737_3781), 
      .ZN(n_1_737_3779));
   OAI22_X1 i_1_737_4282 (.A1(\out_bs[1] [6]), .A2(n_1_737_3784), .B1(
      n_1_737_5297), .B2(n_1_737_3782), .ZN(n_1_737_3780));
   INV_X1 i_1_737_4283 (.A(n_1_737_3782), .ZN(n_1_737_3781));
   NOR2_X1 i_1_737_4284 (.A1(\out_as[1] [6]), .A2(n_1_737_365), .ZN(n_1_737_3782));
   NOR2_X1 i_1_737_4285 (.A1(\out_bs[1] [6]), .A2(n_1_737_3789), .ZN(
      n_1_737_3783));
   INV_X1 i_1_737_4286 (.A(n_1_737_3785), .ZN(n_1_737_3784));
   OAI21_X1 i_1_737_4287 (.A(\out_bs[1] [5]), .B1(\out_bs[1] [4]), .B2(
      n_1_737_4841), .ZN(n_1_737_3785));
   INV_X1 i_1_737_4288 (.A(n_1_737_3787), .ZN(n_1_737_3786));
   OAI21_X1 i_1_737_4289 (.A(\out_bs[1] [5]), .B1(\out_bs[1] [4]), .B2(
      n_1_737_4845), .ZN(n_1_737_3787));
   INV_X1 i_1_737_4290 (.A(n_1_737_3789), .ZN(n_1_737_3788));
   NOR2_X1 i_1_737_4291 (.A1(n_1_737_5663), .A2(n_1_737_5662), .ZN(n_1_737_3789));
   AOI21_X1 i_1_737_4292 (.A(n_1_737_3791), .B1(n_1_737_5189), .B2(n_1_737_3793), 
      .ZN(n_1_737_3790));
   INV_X1 i_1_737_4293 (.A(n_1_737_3792), .ZN(n_1_737_3791));
   OAI21_X1 i_1_737_4294 (.A(n_1_737_3794), .B1(n_1_737_5189), .B2(n_1_737_3793), 
      .ZN(n_1_737_3792));
   NOR2_X1 i_1_737_4295 (.A1(\out_as[3] [6]), .A2(n_1_737_367), .ZN(n_1_737_3793));
   OAI21_X1 i_1_737_4296 (.A(n_1_737_5638), .B1(n_1_737_5637), .B2(n_1_737_4829), 
      .ZN(n_1_737_3794));
   NAND2_X1 i_1_737_4297 (.A1(n_1_737_5638), .A2(n_1_737_3798), .ZN(n_1_737_3795));
   INV_X1 i_1_737_4298 (.A(n_1_737_3797), .ZN(n_1_737_3796));
   NOR2_X1 i_1_737_4299 (.A1(\out_bs[3] [6]), .A2(n_1_737_3799), .ZN(
      n_1_737_3797));
   OAI21_X1 i_1_737_4300 (.A(\out_bs[3] [5]), .B1(\out_bs[3] [4]), .B2(
      n_1_737_4835), .ZN(n_1_737_3798));
   NOR2_X1 i_1_737_4301 (.A1(n_1_737_5637), .A2(n_1_737_5636), .ZN(n_1_737_3799));
   INV_X1 i_1_737_4302 (.A(n_1_737_3801), .ZN(n_1_737_3800));
   OAI21_X1 i_1_737_4303 (.A(n_1_737_3802), .B1(n_1_737_5366), .B2(n_1_737_3803), 
      .ZN(n_1_737_3801));
   OAI22_X1 i_1_737_4304 (.A1(\out_bs[4] [6]), .A2(n_1_737_3807), .B1(
      n_1_737_5365), .B2(n_1_737_3804), .ZN(n_1_737_3802));
   INV_X1 i_1_737_4305 (.A(n_1_737_3804), .ZN(n_1_737_3803));
   NOR2_X1 i_1_737_4306 (.A1(\out_as[4] [6]), .A2(n_1_737_368), .ZN(n_1_737_3804));
   INV_X1 i_1_737_4307 (.A(n_1_737_3806), .ZN(n_1_737_3805));
   NOR2_X1 i_1_737_4308 (.A1(\out_bs[4] [6]), .A2(n_1_737_3810), .ZN(
      n_1_737_3806));
   INV_X1 i_1_737_4309 (.A(n_1_737_3808), .ZN(n_1_737_3807));
   OAI21_X1 i_1_737_4310 (.A(\out_bs[4] [5]), .B1(\out_bs[4] [4]), .B2(
      n_1_737_4860), .ZN(n_1_737_3808));
   OAI21_X1 i_1_737_4311 (.A(\out_bs[4] [5]), .B1(\out_bs[4] [4]), .B2(
      n_1_737_4863), .ZN(n_1_737_3809));
   NOR2_X1 i_1_737_4312 (.A1(n_1_737_5624), .A2(n_1_737_5623), .ZN(n_1_737_3810));
   NOR3_X1 i_1_737_4313 (.A1(\out_as[6] [6]), .A2(n_1_737_363), .A3(n_1_737_4010), 
      .ZN(n_502));
   OAI21_X1 i_1_737_4314 (.A(n_1_737_4010), .B1(\out_as[6] [6]), .B2(n_1_737_363), 
      .ZN(n_503));
   NOR3_X1 i_1_737_4315 (.A1(\out_as[5] [6]), .A2(n_1_737_362), .A3(n_1_737_4019), 
      .ZN(n_504));
   OAI21_X1 i_1_737_4316 (.A(n_1_737_4019), .B1(\out_as[5] [6]), .B2(n_1_737_362), 
      .ZN(n_505));
   NAND4_X1 i_1_737_4317 (.A1(n_1_737_3822), .A2(n_1_737_3820), .A3(n_1_737_3826), 
      .A4(n_1_737_3811), .ZN(n_506));
   AOI211_X1 i_1_737_4318 (.A(n_1_737_3812), .B(n_1_737_3816), .C1(n_1_737_4027), 
      .C2(n_1_737_3821), .ZN(n_1_737_3811));
   INV_X1 i_1_737_4319 (.A(n_1_737_3813), .ZN(n_1_737_3812));
   AOI22_X1 i_1_737_4320 (.A1(n_1_737_4035), .A2(n_1_737_3815), .B1(n_1_737_5189), 
      .B2(n_1_737_3814), .ZN(n_1_737_3813));
   OAI21_X1 i_1_737_4321 (.A(n_1_737_4036), .B1(\out_as[3] [6]), .B2(n_1_737_360), 
      .ZN(n_1_737_3814));
   NOR2_X1 i_1_737_4322 (.A1(\out_as[3] [6]), .A2(n_1_737_360), .ZN(n_1_737_3815));
   INV_X1 i_1_737_4323 (.A(n_1_737_3817), .ZN(n_1_737_3816));
   AOI22_X1 i_1_737_4324 (.A1(n_1_737_4068), .A2(n_1_737_3819), .B1(n_1_737_5365), 
      .B2(n_1_737_3818), .ZN(n_1_737_3817));
   OAI21_X1 i_1_737_4325 (.A(n_1_737_4069), .B1(\out_as[4] [6]), .B2(n_1_737_361), 
      .ZN(n_1_737_3818));
   NOR2_X1 i_1_737_4326 (.A1(\out_as[4] [6]), .A2(n_1_737_361), .ZN(n_1_737_3819));
   OAI21_X1 i_1_737_4327 (.A(n_1_737_5336), .B1(n_1_737_4027), .B2(n_1_737_3821), 
      .ZN(n_1_737_3820));
   NOR2_X1 i_1_737_4328 (.A1(\out_as[0] [6]), .A2(n_1_737_357), .ZN(n_1_737_3821));
   AOI22_X1 i_1_737_4329 (.A1(n_1_737_4057), .A2(n_1_737_3824), .B1(n_1_737_5235), 
      .B2(n_1_737_3823), .ZN(n_1_737_3822));
   OAI21_X1 i_1_737_4330 (.A(n_1_737_4058), .B1(\out_as[2] [6]), .B2(n_1_737_359), 
      .ZN(n_1_737_3823));
   NOR2_X1 i_1_737_4331 (.A1(\out_as[2] [6]), .A2(n_1_737_359), .ZN(n_1_737_3824));
   INV_X1 i_1_737_4332 (.A(n_1_737_3826), .ZN(n_1_737_3825));
   OAI21_X1 i_1_737_4333 (.A(n_1_737_3827), .B1(n_1_737_5297), .B2(n_1_737_3829), 
      .ZN(n_1_737_3826));
   OAI21_X1 i_1_737_4334 (.A(n_1_737_4045), .B1(n_1_737_5298), .B2(n_1_737_3828), 
      .ZN(n_1_737_3827));
   INV_X1 i_1_737_4335 (.A(n_1_737_3829), .ZN(n_1_737_3828));
   NOR2_X1 i_1_737_4336 (.A1(\out_as[1] [6]), .A2(n_1_737_358), .ZN(n_1_737_3829));
   NOR3_X1 i_1_737_4337 (.A1(\out_as[6] [6]), .A2(n_1_737_356), .A3(n_1_737_3830), 
      .ZN(n_507));
   OAI21_X1 i_1_737_4338 (.A(n_1_737_3830), .B1(\out_as[6] [6]), .B2(n_1_737_356), 
      .ZN(n_508));
   AOI21_X1 i_1_737_4339 (.A(\out_bs[6] [6]), .B1(\out_bs[6] [5]), .B2(
      n_1_737_3831), .ZN(n_1_737_3830));
   OAI21_X1 i_1_737_4340 (.A(n_1_737_4919), .B1(n_1_737_5603), .B2(n_1_737_3943), 
      .ZN(n_1_737_3831));
   NOR3_X1 i_1_737_4341 (.A1(\out_as[5] [6]), .A2(n_1_737_355), .A3(n_1_737_3832), 
      .ZN(n_509));
   OAI21_X1 i_1_737_4342 (.A(n_1_737_3832), .B1(\out_as[5] [6]), .B2(n_1_737_355), 
      .ZN(n_510));
   AOI21_X1 i_1_737_4343 (.A(n_844), .B1(n_845), .B2(n_1_737_4881), .ZN(
      n_1_737_3832));
   NAND4_X1 i_1_737_4344 (.A1(n_1_737_3848), .A2(n_1_737_3836), .A3(n_1_737_3852), 
      .A4(n_1_737_3833), .ZN(n_511));
   AOI211_X1 i_1_737_4345 (.A(n_1_737_3834), .B(n_1_737_3843), .C1(n_1_737_5336), 
      .C2(n_1_737_3840), .ZN(n_1_737_3833));
   INV_X1 i_1_737_4346 (.A(n_1_737_3835), .ZN(n_1_737_3834));
   OAI21_X1 i_1_737_4347 (.A(n_1_737_3841), .B1(n_1_737_5336), .B2(n_1_737_3840), 
      .ZN(n_1_737_3835));
   AOI22_X1 i_1_737_4348 (.A1(n_1_737_3839), .A2(n_1_737_3838), .B1(n_1_737_5189), 
      .B2(n_1_737_3837), .ZN(n_1_737_3836));
   OR2_X1 i_1_737_4349 (.A1(n_1_737_3839), .A2(n_1_737_3838), .ZN(n_1_737_3837));
   OAI21_X1 i_1_737_4350 (.A(n_1_737_4036), .B1(n_1_737_5637), .B2(n_1_737_4895), 
      .ZN(n_1_737_3838));
   NOR2_X1 i_1_737_4351 (.A1(\out_as[3] [6]), .A2(n_1_737_353), .ZN(n_1_737_3839));
   NOR2_X1 i_1_737_4352 (.A1(\out_as[0] [6]), .A2(n_1_737_350), .ZN(n_1_737_3840));
   OAI21_X1 i_1_737_4353 (.A(n_1_737_5671), .B1(n_1_737_5670), .B2(n_1_737_4904), 
      .ZN(n_1_737_3841));
   INV_X1 i_1_737_4354 (.A(n_1_737_3843), .ZN(n_1_737_3842));
   OAI21_X1 i_1_737_4355 (.A(n_1_737_3844), .B1(n_1_737_5298), .B2(n_1_737_3845), 
      .ZN(n_1_737_3843));
   OAI21_X1 i_1_737_4356 (.A(n_1_737_3847), .B1(n_1_737_5297), .B2(n_1_737_3846), 
      .ZN(n_1_737_3844));
   INV_X1 i_1_737_4357 (.A(n_1_737_3846), .ZN(n_1_737_3845));
   NOR2_X1 i_1_737_4358 (.A1(\out_as[1] [6]), .A2(n_1_737_351), .ZN(n_1_737_3846));
   OAI21_X1 i_1_737_4359 (.A(n_1_737_4045), .B1(n_1_737_5663), .B2(n_1_737_4889), 
      .ZN(n_1_737_3847));
   OAI21_X1 i_1_737_4360 (.A(n_1_737_3849), .B1(n_1_737_5235), .B2(n_1_737_3850), 
      .ZN(n_1_737_3848));
   OAI22_X1 i_1_737_4361 (.A1(\out_as[2] [6]), .A2(n_1_737_352), .B1(
      n_1_737_5236), .B2(n_1_737_3851), .ZN(n_1_737_3849));
   INV_X1 i_1_737_4362 (.A(n_1_737_3851), .ZN(n_1_737_3850));
   AOI21_X1 i_1_737_4363 (.A(n_1_737_4057), .B1(\out_bs[2] [5]), .B2(
      n_1_737_4901), .ZN(n_1_737_3851));
   OAI21_X1 i_1_737_4364 (.A(n_1_737_3853), .B1(n_1_737_5365), .B2(n_1_737_3855), 
      .ZN(n_1_737_3852));
   OAI22_X1 i_1_737_4365 (.A1(\out_as[4] [6]), .A2(n_1_737_354), .B1(
      n_1_737_5366), .B2(n_1_737_3854), .ZN(n_1_737_3853));
   INV_X1 i_1_737_4366 (.A(n_1_737_3855), .ZN(n_1_737_3854));
   OAI21_X1 i_1_737_4367 (.A(n_1_737_4069), .B1(n_1_737_5624), .B2(n_1_737_4911), 
      .ZN(n_1_737_3855));
   NOR3_X1 i_1_737_4368 (.A1(\out_as[6] [6]), .A2(n_1_737_349), .A3(n_1_737_3856), 
      .ZN(n_512));
   OAI21_X1 i_1_737_4369 (.A(n_1_737_3856), .B1(\out_as[6] [6]), .B2(n_1_737_349), 
      .ZN(n_513));
   AOI21_X1 i_1_737_4370 (.A(\out_bs[6] [6]), .B1(\out_bs[6] [5]), .B2(
      n_1_737_4917), .ZN(n_1_737_3856));
   NOR3_X1 i_1_737_4371 (.A1(\out_as[5] [6]), .A2(n_1_737_348), .A3(n_1_737_3857), 
      .ZN(n_514));
   OAI21_X1 i_1_737_4372 (.A(n_1_737_3857), .B1(\out_as[5] [6]), .B2(n_1_737_348), 
      .ZN(n_515));
   AOI21_X1 i_1_737_4373 (.A(n_844), .B1(n_845), .B2(n_1_737_4922), .ZN(
      n_1_737_3857));
   NAND4_X1 i_1_737_4374 (.A1(n_1_737_3877), .A2(n_1_737_3859), .A3(n_1_737_3865), 
      .A4(n_1_737_3858), .ZN(n_516));
   AND3_X1 i_1_737_4375 (.A1(n_1_737_3874), .A2(n_1_737_3873), .A3(n_1_737_3869), 
      .ZN(n_1_737_3858));
   INV_X1 i_1_737_4376 (.A(n_1_737_3860), .ZN(n_1_737_3859));
   OAI21_X1 i_1_737_4377 (.A(n_1_737_3861), .B1(n_1_737_5298), .B2(n_1_737_3862), 
      .ZN(n_1_737_3860));
   OAI21_X1 i_1_737_4378 (.A(n_1_737_3864), .B1(n_1_737_5297), .B2(n_1_737_3863), 
      .ZN(n_1_737_3861));
   INV_X1 i_1_737_4379 (.A(n_1_737_3863), .ZN(n_1_737_3862));
   NOR2_X1 i_1_737_4380 (.A1(\out_as[1] [6]), .A2(n_1_737_344), .ZN(n_1_737_3863));
   OAI21_X1 i_1_737_4381 (.A(n_1_737_5664), .B1(n_1_737_5663), .B2(n_1_737_4932), 
      .ZN(n_1_737_3864));
   AOI22_X1 i_1_737_4382 (.A1(n_1_737_3868), .A2(n_1_737_3867), .B1(n_1_737_5189), 
      .B2(n_1_737_3866), .ZN(n_1_737_3865));
   OR2_X1 i_1_737_4383 (.A1(n_1_737_3868), .A2(n_1_737_3867), .ZN(n_1_737_3866));
   OAI21_X1 i_1_737_4384 (.A(n_1_737_5638), .B1(n_1_737_5637), .B2(n_1_737_4939), 
      .ZN(n_1_737_3867));
   NOR2_X1 i_1_737_4385 (.A1(\out_as[3] [6]), .A2(n_1_737_346), .ZN(n_1_737_3868));
   OAI21_X1 i_1_737_4386 (.A(n_1_737_3870), .B1(n_1_737_5235), .B2(n_1_737_3872), 
      .ZN(n_1_737_3869));
   OAI22_X1 i_1_737_4387 (.A1(\out_as[2] [6]), .A2(n_1_737_345), .B1(
      n_1_737_5236), .B2(n_1_737_3871), .ZN(n_1_737_3870));
   INV_X1 i_1_737_4388 (.A(n_1_737_3872), .ZN(n_1_737_3871));
   OAI21_X1 i_1_737_4389 (.A(n_1_737_5651), .B1(n_1_737_5650), .B2(n_1_737_4953), 
      .ZN(n_1_737_3872));
   NAND2_X1 i_1_737_4390 (.A1(n_1_737_5336), .A2(n_1_737_3875), .ZN(n_1_737_3873));
   OAI21_X1 i_1_737_4391 (.A(n_1_737_3876), .B1(n_1_737_5336), .B2(n_1_737_3875), 
      .ZN(n_1_737_3874));
   NOR2_X1 i_1_737_4392 (.A1(\out_as[0] [6]), .A2(n_1_737_343), .ZN(n_1_737_3875));
   OAI21_X1 i_1_737_4393 (.A(n_1_737_5671), .B1(n_1_737_5670), .B2(n_1_737_4946), 
      .ZN(n_1_737_3876));
   OAI21_X1 i_1_737_4394 (.A(n_1_737_3878), .B1(n_1_737_5365), .B2(n_1_737_3880), 
      .ZN(n_1_737_3877));
   OAI22_X1 i_1_737_4395 (.A1(\out_as[4] [6]), .A2(n_1_737_347), .B1(
      n_1_737_5366), .B2(n_1_737_3879), .ZN(n_1_737_3878));
   INV_X1 i_1_737_4396 (.A(n_1_737_3880), .ZN(n_1_737_3879));
   OAI21_X1 i_1_737_4397 (.A(n_1_737_5625), .B1(n_1_737_5624), .B2(n_1_737_4960), 
      .ZN(n_1_737_3880));
   NOR3_X1 i_1_737_4398 (.A1(\out_as[6] [6]), .A2(n_1_737_342), .A3(n_1_737_3881), 
      .ZN(n_517));
   OAI21_X1 i_1_737_4399 (.A(n_1_737_3881), .B1(\out_as[6] [6]), .B2(n_1_737_342), 
      .ZN(n_518));
   AOI21_X1 i_1_737_4400 (.A(\out_bs[6] [6]), .B1(\out_bs[6] [5]), .B2(
      n_1_737_3882), .ZN(n_1_737_3881));
   NAND2_X1 i_1_737_4401 (.A1(n_1_737_4919), .A2(n_1_737_3884), .ZN(n_1_737_3882));
   INV_X1 i_1_737_4402 (.A(n_1_737_3884), .ZN(n_1_737_3883));
   OAI21_X1 i_1_737_4403 (.A(n_851), .B1(n_1311), .B2(\out_bs[6] [0]), .ZN(
      n_1_737_3884));
   NOR3_X1 i_1_737_4404 (.A1(\out_as[5] [6]), .A2(n_1_737_341), .A3(n_1_737_3885), 
      .ZN(n_519));
   OAI21_X1 i_1_737_4405 (.A(n_1_737_3885), .B1(\out_as[5] [6]), .B2(n_1_737_341), 
      .ZN(n_520));
   AOI21_X1 i_1_737_4406 (.A(n_844), .B1(n_845), .B2(n_1_737_4963), .ZN(
      n_1_737_3885));
   NAND4_X1 i_1_737_4407 (.A1(n_1_737_3909), .A2(n_1_737_3897), .A3(n_1_737_3892), 
      .A4(n_1_737_3886), .ZN(n_521));
   AOI211_X1 i_1_737_4408 (.A(n_1_737_3887), .B(n_1_737_3904), .C1(n_1_737_5336), 
      .C2(n_1_737_3889), .ZN(n_1_737_3886));
   AOI22_X1 i_1_737_4409 (.A1(n_1_737_5671), .A2(n_1_737_3890), .B1(n_1_737_5337), 
      .B2(n_1_737_3888), .ZN(n_1_737_3887));
   INV_X1 i_1_737_4410 (.A(n_1_737_3889), .ZN(n_1_737_3888));
   NOR2_X1 i_1_737_4411 (.A1(\out_as[0] [6]), .A2(n_1_737_336), .ZN(n_1_737_3889));
   AOI22_X1 i_1_737_4412 (.A1(\out_bs[0] [5]), .A2(n_1_737_5333), .B1(
      \out_bs[0] [2]), .B2(n_1_737_4029), .ZN(n_1_737_3890));
   INV_X1 i_1_737_4413 (.A(n_1_737_3892), .ZN(n_1_737_3891));
   OAI21_X1 i_1_737_4414 (.A(n_1_737_3893), .B1(n_1_737_5189), .B2(n_1_737_3894), 
      .ZN(n_1_737_3892));
   OAI22_X1 i_1_737_4415 (.A1(\out_as[3] [6]), .A2(n_1_737_339), .B1(
      n_1_737_5190), .B2(n_1_737_3895), .ZN(n_1_737_3893));
   INV_X1 i_1_737_4416 (.A(n_1_737_3895), .ZN(n_1_737_3894));
   NOR2_X1 i_1_737_4417 (.A1(n_1_737_4035), .A2(n_1_737_3896), .ZN(n_1_737_3895));
   NOR3_X1 i_1_737_4418 (.A1(n_1_737_5637), .A2(n_1_737_5634), .A3(n_1_737_5232), 
      .ZN(n_1_737_3896));
   INV_X1 i_1_737_4419 (.A(n_1_737_3898), .ZN(n_1_737_3897));
   OAI21_X1 i_1_737_4420 (.A(n_1_737_3899), .B1(n_1_737_5298), .B2(n_1_737_3900), 
      .ZN(n_1_737_3898));
   OAI22_X1 i_1_737_4421 (.A1(\out_bs[1] [6]), .A2(n_1_737_3902), .B1(
      n_1_737_5297), .B2(n_1_737_3901), .ZN(n_1_737_3899));
   INV_X1 i_1_737_4422 (.A(n_1_737_3901), .ZN(n_1_737_3900));
   NOR2_X1 i_1_737_4423 (.A1(\out_as[1] [6]), .A2(n_1_737_337), .ZN(n_1_737_3901));
   INV_X1 i_1_737_4424 (.A(n_1_737_3903), .ZN(n_1_737_3902));
   AOI21_X1 i_1_737_4425 (.A(n_1_737_4050), .B1(\out_bs[1] [2]), .B2(
      n_1_737_4051), .ZN(n_1_737_3903));
   OAI21_X1 i_1_737_4426 (.A(n_1_737_3905), .B1(n_1_737_5236), .B2(n_1_737_3906), 
      .ZN(n_1_737_3904));
   OAI22_X1 i_1_737_4427 (.A1(\out_bs[2] [6]), .A2(n_1_737_3908), .B1(
      n_1_737_5235), .B2(n_1_737_3907), .ZN(n_1_737_3905));
   INV_X1 i_1_737_4428 (.A(n_1_737_3907), .ZN(n_1_737_3906));
   NOR2_X1 i_1_737_4429 (.A1(\out_as[2] [6]), .A2(n_1_737_338), .ZN(n_1_737_3907));
   AOI21_X1 i_1_737_4430 (.A(n_1_737_5650), .B1(n_1_737_5649), .B2(n_1_737_4985), 
      .ZN(n_1_737_3908));
   INV_X1 i_1_737_4431 (.A(n_1_737_3910), .ZN(n_1_737_3909));
   OAI21_X1 i_1_737_4432 (.A(n_1_737_3911), .B1(n_1_737_5366), .B2(n_1_737_3912), 
      .ZN(n_1_737_3910));
   OAI22_X1 i_1_737_4433 (.A1(\out_bs[4] [6]), .A2(n_1_737_3915), .B1(
      n_1_737_5365), .B2(n_1_737_3913), .ZN(n_1_737_3911));
   INV_X1 i_1_737_4434 (.A(n_1_737_3913), .ZN(n_1_737_3912));
   NOR2_X1 i_1_737_4435 (.A1(\out_as[4] [6]), .A2(n_1_737_340), .ZN(n_1_737_3913));
   INV_X1 i_1_737_4436 (.A(n_1_737_3915), .ZN(n_1_737_3914));
   AOI21_X1 i_1_737_4437 (.A(n_1_737_5624), .B1(n_1_737_5623), .B2(n_1_737_4999), 
      .ZN(n_1_737_3915));
   NOR3_X1 i_1_737_4438 (.A1(\out_as[6] [6]), .A2(n_1_737_335), .A3(n_1_737_4009), 
      .ZN(n_522));
   OAI21_X1 i_1_737_4439 (.A(n_1_737_4009), .B1(\out_as[6] [6]), .B2(n_1_737_335), 
      .ZN(n_523));
   NOR3_X1 i_1_737_4440 (.A1(\out_as[5] [6]), .A2(n_1_737_334), .A3(n_1_737_4018), 
      .ZN(n_524));
   OAI21_X1 i_1_737_4441 (.A(n_1_737_4018), .B1(\out_as[5] [6]), .B2(n_1_737_334), 
      .ZN(n_525));
   OAI211_X1 i_1_737_4442 (.A(n_1_737_3916), .B(n_1_737_3935), .C1(n_1_737_3932), 
      .C2(n_1_737_3931), .ZN(n_526));
   NOR3_X1 i_1_737_4443 (.A1(n_1_737_3922), .A2(n_1_737_3918), .A3(n_1_737_3926), 
      .ZN(n_1_737_3916));
   INV_X1 i_1_737_4444 (.A(n_1_737_3918), .ZN(n_1_737_3917));
   OAI21_X1 i_1_737_4445 (.A(n_1_737_3919), .B1(n_1_737_5298), .B2(n_1_737_3920), 
      .ZN(n_1_737_3918));
   OAI22_X1 i_1_737_4446 (.A1(\out_bs[1] [6]), .A2(n_1_737_4049), .B1(
      n_1_737_5297), .B2(n_1_737_3921), .ZN(n_1_737_3919));
   INV_X1 i_1_737_4447 (.A(n_1_737_3921), .ZN(n_1_737_3920));
   NOR2_X1 i_1_737_4448 (.A1(\out_as[1] [6]), .A2(n_1_737_330), .ZN(n_1_737_3921));
   INV_X1 i_1_737_4449 (.A(n_1_737_3923), .ZN(n_1_737_3922));
   AOI22_X1 i_1_737_4450 (.A1(n_1_737_4034), .A2(n_1_737_3925), .B1(n_1_737_5189), 
      .B2(n_1_737_3924), .ZN(n_1_737_3923));
   OR2_X1 i_1_737_4451 (.A1(n_1_737_4034), .A2(n_1_737_3925), .ZN(n_1_737_3924));
   NOR2_X1 i_1_737_4452 (.A1(\out_as[3] [6]), .A2(n_1_737_332), .ZN(n_1_737_3925));
   INV_X1 i_1_737_4453 (.A(n_1_737_3927), .ZN(n_1_737_3926));
   OAI21_X1 i_1_737_4454 (.A(n_1_737_3928), .B1(n_1_737_5235), .B2(n_1_737_3930), 
      .ZN(n_1_737_3927));
   OAI211_X1 i_1_737_4455 (.A(n_1_737_5651), .B(n_1_737_4061), .C1(n_1_737_5236), 
      .C2(n_1_737_3929), .ZN(n_1_737_3928));
   INV_X1 i_1_737_4456 (.A(n_1_737_3930), .ZN(n_1_737_3929));
   NOR2_X1 i_1_737_4457 (.A1(\out_as[2] [6]), .A2(n_1_737_331), .ZN(n_1_737_3930));
   NOR2_X1 i_1_737_4458 (.A1(n_1_737_4026), .A2(n_1_737_3933), .ZN(n_1_737_3931));
   AOI21_X1 i_1_737_4459 (.A(n_1_737_5336), .B1(n_1_737_4026), .B2(n_1_737_3933), 
      .ZN(n_1_737_3932));
   NOR2_X1 i_1_737_4460 (.A1(\out_as[0] [6]), .A2(n_1_737_329), .ZN(n_1_737_3933));
   INV_X1 i_1_737_4461 (.A(n_1_737_3935), .ZN(n_1_737_3934));
   OAI21_X1 i_1_737_4462 (.A(n_1_737_3936), .B1(n_1_737_5365), .B2(n_1_737_3938), 
      .ZN(n_1_737_3935));
   OAI211_X1 i_1_737_4463 (.A(n_1_737_5625), .B(n_1_737_4072), .C1(n_1_737_5366), 
      .C2(n_1_737_3937), .ZN(n_1_737_3936));
   INV_X1 i_1_737_4464 (.A(n_1_737_3938), .ZN(n_1_737_3937));
   NOR2_X1 i_1_737_4465 (.A1(\out_as[4] [6]), .A2(n_1_737_333), .ZN(n_1_737_3938));
   NOR3_X1 i_1_737_4466 (.A1(\out_as[6] [6]), .A2(n_1_737_328), .A3(n_1_737_3939), 
      .ZN(n_527));
   OAI21_X1 i_1_737_4467 (.A(n_1_737_3939), .B1(\out_as[6] [6]), .B2(n_1_737_328), 
      .ZN(n_528));
   NOR3_X1 i_1_737_4468 (.A1(\out_bs[6] [6]), .A2(n_1_737_4012), .A3(
      n_1_737_3940), .ZN(n_1_737_3939));
   NOR2_X1 i_1_737_4469 (.A1(n_1_737_5606), .A2(n_1_737_3943), .ZN(n_1_737_3940));
   NOR2_X1 i_1_737_4470 (.A1(n_847), .A2(n_1_737_3942), .ZN(n_1_737_3941));
   NAND2_X1 i_1_737_4471 (.A1(n_1_737_5603), .A2(n_1_737_3943), .ZN(n_1_737_3942));
   NAND2_X1 i_1_737_4472 (.A1(n_1311), .A2(\out_bs[6] [0]), .ZN(n_1_737_3943));
   NOR3_X1 i_1_737_4473 (.A1(\out_as[5] [6]), .A2(n_1_737_327), .A3(n_1_737_3944), 
      .ZN(n_529));
   OAI21_X1 i_1_737_4474 (.A(n_1_737_3944), .B1(\out_as[5] [6]), .B2(n_1_737_327), 
      .ZN(n_530));
   NOR2_X1 i_1_737_4475 (.A1(n_1_737_4017), .A2(n_1_737_3945), .ZN(n_1_737_3944));
   NOR2_X1 i_1_737_4476 (.A1(n_1_737_5611), .A2(n_1_737_5023), .ZN(n_1_737_3945));
   OR4_X1 i_1_737_4477 (.A1(n_1_737_3952), .A2(n_1_737_3946), .A3(n_1_737_3958), 
      .A4(n_1_737_3972), .ZN(n_531));
   OAI21_X1 i_1_737_4478 (.A(n_1_737_3947), .B1(n_1_737_5236), .B2(n_1_737_3948), 
      .ZN(n_1_737_3946));
   OAI22_X1 i_1_737_4479 (.A1(\out_bs[2] [6]), .A2(n_1_737_3950), .B1(
      n_1_737_5235), .B2(n_1_737_3949), .ZN(n_1_737_3947));
   INV_X1 i_1_737_4480 (.A(n_1_737_3949), .ZN(n_1_737_3948));
   NOR2_X1 i_1_737_4481 (.A1(\out_as[2] [6]), .A2(n_1_737_324), .ZN(n_1_737_3949));
   INV_X1 i_1_737_4482 (.A(n_1_737_3951), .ZN(n_1_737_3950));
   OAI21_X1 i_1_737_4483 (.A(\out_bs[2] [5]), .B1(\out_bs[2] [4]), .B2(
      n_1_737_5053), .ZN(n_1_737_3951));
   INV_X1 i_1_737_4484 (.A(n_1_737_3953), .ZN(n_1_737_3952));
   OAI21_X1 i_1_737_4485 (.A(n_1_737_3954), .B1(n_1_737_5189), .B2(n_1_737_3956), 
      .ZN(n_1_737_3953));
   OAI22_X1 i_1_737_4486 (.A1(\out_as[3] [6]), .A2(n_1_737_325), .B1(
      n_1_737_5190), .B2(n_1_737_3955), .ZN(n_1_737_3954));
   INV_X1 i_1_737_4487 (.A(n_1_737_3956), .ZN(n_1_737_3955));
   NAND2_X1 i_1_737_4488 (.A1(n_1_737_5638), .A2(n_1_737_3957), .ZN(n_1_737_3956));
   OAI21_X1 i_1_737_4489 (.A(\out_bs[3] [5]), .B1(\out_bs[3] [4]), .B2(
      n_1_737_5035), .ZN(n_1_737_3957));
   OAI211_X1 i_1_737_4490 (.A(n_1_737_3959), .B(n_1_737_3964), .C1(n_1_737_5337), 
      .C2(n_1_737_3960), .ZN(n_1_737_3958));
   OAI22_X1 i_1_737_4491 (.A1(\out_bs[0] [6]), .A2(n_1_737_3962), .B1(
      n_1_737_5336), .B2(n_1_737_3961), .ZN(n_1_737_3959));
   INV_X1 i_1_737_4492 (.A(n_1_737_3961), .ZN(n_1_737_3960));
   NOR2_X1 i_1_737_4493 (.A1(\out_as[0] [6]), .A2(n_1_737_322), .ZN(n_1_737_3961));
   INV_X1 i_1_737_4494 (.A(n_1_737_3963), .ZN(n_1_737_3962));
   OAI21_X1 i_1_737_4495 (.A(\out_bs[0] [5]), .B1(\out_bs[0] [4]), .B2(
      n_1_737_5027), .ZN(n_1_737_3963));
   INV_X1 i_1_737_4496 (.A(n_1_737_3965), .ZN(n_1_737_3964));
   OAI21_X1 i_1_737_4497 (.A(n_1_737_3966), .B1(n_1_737_5298), .B2(n_1_737_3967), 
      .ZN(n_1_737_3965));
   OAI22_X1 i_1_737_4498 (.A1(\out_bs[1] [6]), .A2(n_1_737_3969), .B1(
      n_1_737_5297), .B2(n_1_737_3968), .ZN(n_1_737_3966));
   INV_X1 i_1_737_4499 (.A(n_1_737_3968), .ZN(n_1_737_3967));
   NOR2_X1 i_1_737_4500 (.A1(\out_as[1] [6]), .A2(n_1_737_323), .ZN(n_1_737_3968));
   INV_X1 i_1_737_4501 (.A(n_1_737_3970), .ZN(n_1_737_3969));
   OAI21_X1 i_1_737_4502 (.A(\out_bs[1] [5]), .B1(\out_bs[1] [4]), .B2(
      n_1_737_5046), .ZN(n_1_737_3970));
   INV_X1 i_1_737_4503 (.A(n_1_737_3972), .ZN(n_1_737_3971));
   OAI21_X1 i_1_737_4504 (.A(n_1_737_3973), .B1(n_1_737_5366), .B2(n_1_737_3974), 
      .ZN(n_1_737_3972));
   OAI22_X1 i_1_737_4505 (.A1(\out_bs[4] [6]), .A2(n_1_737_3976), .B1(
      n_1_737_5365), .B2(n_1_737_3975), .ZN(n_1_737_3973));
   INV_X1 i_1_737_4506 (.A(n_1_737_3975), .ZN(n_1_737_3974));
   NOR2_X1 i_1_737_4507 (.A1(\out_as[4] [6]), .A2(n_1_737_326), .ZN(n_1_737_3975));
   INV_X1 i_1_737_4508 (.A(n_1_737_3977), .ZN(n_1_737_3976));
   OAI21_X1 i_1_737_4509 (.A(\out_bs[4] [5]), .B1(\out_bs[4] [4]), .B2(
      n_1_737_5062), .ZN(n_1_737_3977));
   NOR3_X1 i_1_737_4510 (.A1(\out_as[6] [6]), .A2(n_1_737_321), .A3(n_1_737_3978), 
      .ZN(n_532));
   OAI21_X1 i_1_737_4511 (.A(n_1_737_3978), .B1(\out_as[6] [6]), .B2(n_1_737_321), 
      .ZN(n_533));
   INV_X1 i_1_737_4512 (.A(n_1_737_3979), .ZN(n_1_737_3978));
   OAI21_X1 i_1_737_4513 (.A(n_1_737_4010), .B1(n_1_737_4915), .B2(n_1_737_4515), 
      .ZN(n_1_737_3979));
   NOR3_X1 i_1_737_4514 (.A1(\out_as[5] [6]), .A2(n_1_737_320), .A3(n_1_737_3980), 
      .ZN(n_534));
   OAI21_X1 i_1_737_4515 (.A(n_1_737_3980), .B1(\out_as[5] [6]), .B2(n_1_737_320), 
      .ZN(n_535));
   AOI21_X1 i_1_737_4516 (.A(n_844), .B1(n_845), .B2(n_1_737_5071), .ZN(
      n_1_737_3980));
   OAI211_X1 i_1_737_4517 (.A(n_1_737_4003), .B(n_1_737_3981), .C1(n_1_737_5337), 
      .C2(n_1_737_4005), .ZN(n_536));
   NOR4_X1 i_1_737_4518 (.A1(n_1_737_3988), .A2(n_1_737_3983), .A3(n_1_737_3993), 
      .A4(n_1_737_3998), .ZN(n_1_737_3981));
   INV_X1 i_1_737_4519 (.A(n_1_737_3983), .ZN(n_1_737_3982));
   OAI21_X1 i_1_737_4520 (.A(n_1_737_3984), .B1(n_1_737_5298), .B2(n_1_737_3985), 
      .ZN(n_1_737_3983));
   OAI21_X1 i_1_737_4521 (.A(n_1_737_3987), .B1(n_1_737_5297), .B2(n_1_737_3986), 
      .ZN(n_1_737_3984));
   INV_X1 i_1_737_4522 (.A(n_1_737_3986), .ZN(n_1_737_3985));
   NOR2_X1 i_1_737_4523 (.A1(\out_as[1] [6]), .A2(n_1_737_316), .ZN(n_1_737_3986));
   OAI21_X1 i_1_737_4524 (.A(n_1_737_5664), .B1(n_1_737_5663), .B2(n_1_737_5109), 
      .ZN(n_1_737_3987));
   INV_X1 i_1_737_4525 (.A(n_1_737_3989), .ZN(n_1_737_3988));
   AOI22_X1 i_1_737_4526 (.A1(n_1_737_3992), .A2(n_1_737_3991), .B1(n_1_737_5189), 
      .B2(n_1_737_3990), .ZN(n_1_737_3989));
   OR2_X1 i_1_737_4527 (.A1(n_1_737_3992), .A2(n_1_737_3991), .ZN(n_1_737_3990));
   OAI21_X1 i_1_737_4528 (.A(n_1_737_5638), .B1(n_1_737_5637), .B2(n_1_737_5120), 
      .ZN(n_1_737_3991));
   NOR2_X1 i_1_737_4529 (.A1(\out_as[3] [6]), .A2(n_1_737_318), .ZN(n_1_737_3992));
   INV_X1 i_1_737_4530 (.A(n_1_737_3994), .ZN(n_1_737_3993));
   OAI21_X1 i_1_737_4531 (.A(n_1_737_3995), .B1(n_1_737_5235), .B2(n_1_737_3997), 
      .ZN(n_1_737_3994));
   OAI22_X1 i_1_737_4532 (.A1(\out_as[2] [6]), .A2(n_1_737_317), .B1(
      n_1_737_5236), .B2(n_1_737_3996), .ZN(n_1_737_3995));
   INV_X1 i_1_737_4533 (.A(n_1_737_3997), .ZN(n_1_737_3996));
   OAI21_X1 i_1_737_4534 (.A(n_1_737_5651), .B1(n_1_737_5650), .B2(n_1_737_5093), 
      .ZN(n_1_737_3997));
   INV_X1 i_1_737_4535 (.A(n_1_737_3999), .ZN(n_1_737_3998));
   OAI21_X1 i_1_737_4536 (.A(n_1_737_4000), .B1(n_1_737_5365), .B2(n_1_737_4002), 
      .ZN(n_1_737_3999));
   OAI22_X1 i_1_737_4537 (.A1(\out_as[4] [6]), .A2(n_1_737_319), .B1(
      n_1_737_5366), .B2(n_1_737_4001), .ZN(n_1_737_4000));
   INV_X1 i_1_737_4538 (.A(n_1_737_4002), .ZN(n_1_737_4001));
   OAI21_X1 i_1_737_4539 (.A(n_1_737_5625), .B1(n_1_737_5624), .B2(n_1_737_5128), 
      .ZN(n_1_737_4002));
   OAI21_X1 i_1_737_4540 (.A(n_1_737_4004), .B1(n_1_737_5336), .B2(n_1_737_4006), 
      .ZN(n_1_737_4003));
   OAI21_X1 i_1_737_4541 (.A(n_1_737_5671), .B1(n_1_737_5670), .B2(n_1_737_5079), 
      .ZN(n_1_737_4004));
   INV_X1 i_1_737_4542 (.A(n_1_737_4006), .ZN(n_1_737_4005));
   NOR2_X1 i_1_737_4543 (.A1(\out_as[0] [6]), .A2(n_1_737_315), .ZN(n_1_737_4006));
   NOR3_X1 i_1_737_4544 (.A1(\out_as[6] [6]), .A2(n_1_737_314), .A3(n_1_737_4007), 
      .ZN(n_537));
   OAI21_X1 i_1_737_4545 (.A(n_1_737_4007), .B1(\out_as[6] [6]), .B2(n_1_737_314), 
      .ZN(n_538));
   INV_X1 i_1_737_4546 (.A(n_1_737_4008), .ZN(n_1_737_4007));
   OAI21_X1 i_1_737_4547 (.A(n_1_737_5607), .B1(n_1_737_5606), .B2(n_1_737_4013), 
      .ZN(n_1_737_4008));
   NOR2_X1 i_1_737_4548 (.A1(\out_bs[6] [6]), .A2(n_1_737_4012), .ZN(
      n_1_737_4009));
   AOI21_X1 i_1_737_4549 (.A(\out_bs[6] [6]), .B1(\out_bs[6] [5]), .B2(
      n_1_737_4918), .ZN(n_1_737_4010));
   INV_X1 i_1_737_4550 (.A(n_1_737_4012), .ZN(n_1_737_4011));
   AOI21_X1 i_1_737_4551 (.A(n_1_737_5606), .B1(n_1_737_5605), .B2(n_1_737_4513), 
      .ZN(n_1_737_4012));
   NOR3_X1 i_1_737_4552 (.A1(n_847), .A2(n_1_737_4015), .A3(\out_bs[6] [4]), 
      .ZN(n_1_737_4013));
   NOR2_X1 i_1_737_4553 (.A1(n_847), .A2(n_1_737_4015), .ZN(n_1_737_4014));
   OR2_X1 i_1_737_4554 (.A1(\out_bs[6] [0]), .A2(n_1_737_4514), .ZN(n_1_737_4015));
   NOR3_X1 i_1_737_4555 (.A1(\out_as[5] [6]), .A2(n_1_737_313), .A3(n_1_737_4016), 
      .ZN(n_539));
   OAI21_X1 i_1_737_4556 (.A(n_1_737_4016), .B1(\out_as[5] [6]), .B2(n_1_737_313), 
      .ZN(n_540));
   NOR2_X1 i_1_737_4557 (.A1(n_1_737_4021), .A2(n_1_737_4017), .ZN(n_1_737_4016));
   INV_X1 i_1_737_4558 (.A(n_1_737_4018), .ZN(n_1_737_4017));
   NOR2_X1 i_1_737_4559 (.A1(n_844), .A2(n_1_737_4020), .ZN(n_1_737_4018));
   AOI21_X1 i_1_737_4560 (.A(n_844), .B1(n_845), .B2(n_1_737_5177), .ZN(
      n_1_737_4019));
   AOI21_X1 i_1_737_4561 (.A(n_1_737_5611), .B1(n_1_737_5610), .B2(n_1_737_5175), 
      .ZN(n_1_737_4020));
   NOR2_X1 i_1_737_4562 (.A1(n_1_737_5611), .A2(n_1_737_5183), .ZN(n_1_737_4021));
   OR4_X1 i_1_737_4563 (.A1(n_1_737_4053), .A2(n_1_737_4041), .A3(n_1_737_4022), 
      .A4(n_1_737_4064), .ZN(n_541));
   OAI211_X1 i_1_737_4564 (.A(n_1_737_4023), .B(n_1_737_4030), .C1(n_1_737_5337), 
      .C2(n_1_737_4024), .ZN(n_1_737_4022));
   OAI22_X1 i_1_737_4565 (.A1(n_1_737_4029), .A2(n_1_737_4026), .B1(n_1_737_5336), 
      .B2(n_1_737_4025), .ZN(n_1_737_4023));
   INV_X1 i_1_737_4566 (.A(n_1_737_4025), .ZN(n_1_737_4024));
   NOR2_X1 i_1_737_4567 (.A1(\out_as[0] [6]), .A2(n_1_737_308), .ZN(n_1_737_4025));
   NAND2_X1 i_1_737_4568 (.A1(n_1_737_5671), .A2(n_1_737_4028), .ZN(n_1_737_4026));
   OAI21_X1 i_1_737_4569 (.A(n_1_737_5671), .B1(n_1_737_5670), .B2(n_1_737_5334), 
      .ZN(n_1_737_4027));
   OAI21_X1 i_1_737_4570 (.A(\out_bs[0] [5]), .B1(\out_bs[0] [4]), .B2(
      n_1_737_5328), .ZN(n_1_737_4028));
   NOR2_X1 i_1_737_4571 (.A1(n_1_737_5670), .A2(n_1_737_5335), .ZN(n_1_737_4029));
   OAI21_X1 i_1_737_4572 (.A(n_1_737_4031), .B1(n_1_737_5189), .B2(n_1_737_4033), 
      .ZN(n_1_737_4030));
   OAI22_X1 i_1_737_4573 (.A1(\out_as[3] [6]), .A2(n_1_737_311), .B1(
      n_1_737_5190), .B2(n_1_737_4032), .ZN(n_1_737_4031));
   INV_X1 i_1_737_4574 (.A(n_1_737_4033), .ZN(n_1_737_4032));
   NAND2_X1 i_1_737_4575 (.A1(n_1_737_5638), .A2(n_1_737_4037), .ZN(n_1_737_4033));
   NAND2_X1 i_1_737_4576 (.A1(n_1_737_5638), .A2(n_1_737_4038), .ZN(n_1_737_4034));
   INV_X1 i_1_737_4577 (.A(n_1_737_4036), .ZN(n_1_737_4035));
   NOR2_X1 i_1_737_4578 (.A1(\out_bs[3] [6]), .A2(n_1_737_4039), .ZN(
      n_1_737_4036));
   OAI21_X1 i_1_737_4579 (.A(\out_bs[3] [5]), .B1(\out_bs[3] [4]), .B2(
      n_1_737_5223), .ZN(n_1_737_4037));
   OAI21_X1 i_1_737_4580 (.A(\out_bs[3] [5]), .B1(\out_bs[3] [4]), .B2(
      n_1_737_5224), .ZN(n_1_737_4038));
   NOR2_X1 i_1_737_4581 (.A1(n_1_737_5637), .A2(n_1_737_5231), .ZN(n_1_737_4039));
   INV_X1 i_1_737_4582 (.A(n_1_737_4041), .ZN(n_1_737_4040));
   OAI21_X1 i_1_737_4583 (.A(n_1_737_4042), .B1(n_1_737_5298), .B2(n_1_737_4043), 
      .ZN(n_1_737_4041));
   OAI22_X1 i_1_737_4584 (.A1(\out_bs[1] [6]), .A2(n_1_737_4046), .B1(
      n_1_737_5297), .B2(n_1_737_4044), .ZN(n_1_737_4042));
   INV_X1 i_1_737_4585 (.A(n_1_737_4044), .ZN(n_1_737_4043));
   NOR2_X1 i_1_737_4586 (.A1(\out_as[1] [6]), .A2(n_1_737_309), .ZN(n_1_737_4044));
   NOR2_X1 i_1_737_4587 (.A1(\out_bs[1] [6]), .A2(n_1_737_4050), .ZN(
      n_1_737_4045));
   INV_X1 i_1_737_4588 (.A(n_1_737_4047), .ZN(n_1_737_4046));
   NOR2_X1 i_1_737_4589 (.A1(n_1_737_4051), .A2(n_1_737_4049), .ZN(n_1_737_4047));
   INV_X1 i_1_737_4590 (.A(n_1_737_4049), .ZN(n_1_737_4048));
   AOI21_X1 i_1_737_4591 (.A(n_1_737_5663), .B1(n_1_737_5662), .B2(n_1_737_5289), 
      .ZN(n_1_737_4049));
   NOR2_X1 i_1_737_4592 (.A1(n_1_737_5663), .A2(n_1_737_5295), .ZN(n_1_737_4050));
   NOR2_X1 i_1_737_4593 (.A1(n_1_737_5663), .A2(n_1_737_5296), .ZN(n_1_737_4051));
   INV_X1 i_1_737_4594 (.A(n_1_737_4053), .ZN(n_1_737_4052));
   OAI21_X1 i_1_737_4595 (.A(n_1_737_4054), .B1(n_1_737_5236), .B2(n_1_737_4055), 
      .ZN(n_1_737_4053));
   OAI22_X1 i_1_737_4596 (.A1(\out_bs[2] [6]), .A2(n_1_737_4059), .B1(
      n_1_737_5235), .B2(n_1_737_4056), .ZN(n_1_737_4054));
   INV_X1 i_1_737_4597 (.A(n_1_737_4056), .ZN(n_1_737_4055));
   NOR2_X1 i_1_737_4598 (.A1(\out_as[2] [6]), .A2(n_1_737_310), .ZN(n_1_737_4056));
   INV_X1 i_1_737_4599 (.A(n_1_737_4058), .ZN(n_1_737_4057));
   NOR2_X1 i_1_737_4600 (.A1(\out_bs[2] [6]), .A2(n_1_737_4062), .ZN(
      n_1_737_4058));
   INV_X1 i_1_737_4601 (.A(n_1_737_4060), .ZN(n_1_737_4059));
   OAI21_X1 i_1_737_4602 (.A(\out_bs[2] [5]), .B1(\out_bs[2] [4]), .B2(
      n_1_737_5254), .ZN(n_1_737_4060));
   OAI21_X1 i_1_737_4603 (.A(\out_bs[2] [5]), .B1(\out_bs[2] [4]), .B2(
      n_1_737_5256), .ZN(n_1_737_4061));
   NOR2_X1 i_1_737_4604 (.A1(n_1_737_5650), .A2(n_1_737_5262), .ZN(n_1_737_4062));
   INV_X1 i_1_737_4605 (.A(n_1_737_4064), .ZN(n_1_737_4063));
   OAI21_X1 i_1_737_4606 (.A(n_1_737_4065), .B1(n_1_737_5366), .B2(n_1_737_4066), 
      .ZN(n_1_737_4064));
   OAI22_X1 i_1_737_4607 (.A1(\out_bs[4] [6]), .A2(n_1_737_4070), .B1(
      n_1_737_5365), .B2(n_1_737_4067), .ZN(n_1_737_4065));
   INV_X1 i_1_737_4608 (.A(n_1_737_4067), .ZN(n_1_737_4066));
   NOR2_X1 i_1_737_4609 (.A1(\out_as[4] [6]), .A2(n_1_737_312), .ZN(n_1_737_4067));
   INV_X1 i_1_737_4610 (.A(n_1_737_4069), .ZN(n_1_737_4068));
   NOR2_X1 i_1_737_4611 (.A1(\out_bs[4] [6]), .A2(n_1_737_4073), .ZN(
      n_1_737_4069));
   INV_X1 i_1_737_4612 (.A(n_1_737_4071), .ZN(n_1_737_4070));
   OAI21_X1 i_1_737_4613 (.A(\out_bs[4] [5]), .B1(\out_bs[4] [4]), .B2(
      n_1_737_5394), .ZN(n_1_737_4071));
   OAI21_X1 i_1_737_4614 (.A(\out_bs[4] [5]), .B1(\out_bs[4] [4]), .B2(
      n_1_737_5397), .ZN(n_1_737_4072));
   NOR2_X1 i_1_737_4615 (.A1(n_1_737_5624), .A2(n_1_737_5403), .ZN(n_1_737_4073));
   NOR3_X1 i_1_737_4616 (.A1(\out_as[6] [6]), .A2(n_1_737_307), .A3(n_1_737_4915), 
      .ZN(n_542));
   OAI21_X1 i_1_737_4617 (.A(n_1_737_4915), .B1(\out_as[6] [6]), .B2(n_1_737_307), 
      .ZN(n_543));
   NOR3_X1 i_1_737_4618 (.A1(\out_as[5] [6]), .A2(n_1_737_306), .A3(n_1_737_5182), 
      .ZN(n_544));
   OAI21_X1 i_1_737_4619 (.A(n_1_737_5182), .B1(\out_as[5] [6]), .B2(n_1_737_306), 
      .ZN(n_545));
   NAND4_X1 i_1_737_4620 (.A1(n_1_737_4088), .A2(n_1_737_4074), .A3(n_1_737_4085), 
      .A4(n_1_737_4078), .ZN(n_546));
   AOI211_X1 i_1_737_4621 (.A(n_1_737_4075), .B(n_1_737_4081), .C1(n_1_737_5336), 
      .C2(n_1_737_4077), .ZN(n_1_737_4074));
   INV_X1 i_1_737_4622 (.A(n_1_737_4076), .ZN(n_1_737_4075));
   OAI21_X1 i_1_737_4623 (.A(n_1_737_5083), .B1(n_1_737_5336), .B2(n_1_737_4077), 
      .ZN(n_1_737_4076));
   NOR2_X1 i_1_737_4624 (.A1(\out_as[0] [6]), .A2(n_1_737_301), .ZN(n_1_737_4077));
   AOI21_X1 i_1_737_4625 (.A(n_1_737_4079), .B1(n_1_737_5365), .B2(n_1_737_4080), 
      .ZN(n_1_737_4078));
   NOR3_X1 i_1_737_4626 (.A1(\out_as[4] [6]), .A2(n_1_737_305), .A3(n_1_737_5393), 
      .ZN(n_1_737_4079));
   OAI21_X1 i_1_737_4627 (.A(n_1_737_5393), .B1(\out_as[4] [6]), .B2(n_1_737_305), 
      .ZN(n_1_737_4080));
   INV_X1 i_1_737_4628 (.A(n_1_737_4082), .ZN(n_1_737_4081));
   AOI21_X1 i_1_737_4629 (.A(n_1_737_4083), .B1(n_1_737_5297), .B2(n_1_737_4084), 
      .ZN(n_1_737_4082));
   NOR3_X1 i_1_737_4630 (.A1(\out_as[1] [6]), .A2(n_1_737_302), .A3(n_1_737_5285), 
      .ZN(n_1_737_4083));
   OAI21_X1 i_1_737_4631 (.A(n_1_737_5285), .B1(\out_as[1] [6]), .B2(n_1_737_302), 
      .ZN(n_1_737_4084));
   AOI21_X1 i_1_737_4632 (.A(n_1_737_4086), .B1(n_1_737_5189), .B2(n_1_737_4087), 
      .ZN(n_1_737_4085));
   NOR3_X1 i_1_737_4633 (.A1(\out_as[3] [6]), .A2(n_1_737_304), .A3(n_1_737_5222), 
      .ZN(n_1_737_4086));
   OAI21_X1 i_1_737_4634 (.A(n_1_737_5222), .B1(\out_as[3] [6]), .B2(n_1_737_304), 
      .ZN(n_1_737_4087));
   AOI21_X1 i_1_737_4635 (.A(n_1_737_4089), .B1(n_1_737_5235), .B2(n_1_737_4090), 
      .ZN(n_1_737_4088));
   NOR3_X1 i_1_737_4636 (.A1(\out_as[2] [6]), .A2(n_1_737_303), .A3(n_1_737_5253), 
      .ZN(n_1_737_4089));
   OAI21_X1 i_1_737_4637 (.A(n_1_737_5253), .B1(\out_as[2] [6]), .B2(n_1_737_303), 
      .ZN(n_1_737_4090));
   INV_X1 i_1_737_4638 (.A(n_1_737_4091), .ZN(n_547));
   OAI21_X1 i_1_737_4639 (.A(n_1_737_5168), .B1(n_1_737_5181), .B2(n_1_737_4092), 
      .ZN(n_1_737_4091));
   OAI211_X1 i_1_737_4640 (.A(n_1_737_5182), .B(n_1_737_5167), .C1(n_1_737_5610), 
      .C2(n_1_737_4614), .ZN(n_548));
   NAND4_X1 i_1_737_4642 (.A1(n_1_737_4109), .A2(n_1_737_4102), .A3(n_1_737_4114), 
      .A4(n_1_737_4093), .ZN(n_549));
   INV_X1 i_1_737_4643 (.A(n_1_737_4094), .ZN(n_1_737_4093));
   OAI211_X1 i_1_737_4644 (.A(n_1_737_4095), .B(n_1_737_4097), .C1(n_1_737_5358), 
      .C2(n_1_737_5337), .ZN(n_1_737_4094));
   OAI22_X1 i_1_737_4645 (.A1(n_1_737_5083), .A2(n_1_737_4096), .B1(n_1_737_5359), 
      .B2(n_1_737_5336), .ZN(n_1_737_4095));
   NOR2_X1 i_1_737_4646 (.A1(n_1_737_5669), .A2(n_1_737_4626), .ZN(n_1_737_4096));
   AOI22_X1 i_1_737_4647 (.A1(n_1_737_5387), .A2(n_1_737_4099), .B1(n_1_737_5365), 
      .B2(n_1_737_4098), .ZN(n_1_737_4097));
   NAND3_X1 i_1_737_4648 (.A1(n_1_737_5625), .A2(n_1_737_4100), .A3(n_1_737_5386), 
      .ZN(n_1_737_4098));
   NAND2_X1 i_1_737_4649 (.A1(n_1_737_5625), .A2(n_1_737_4100), .ZN(n_1_737_4099));
   NOR2_X1 i_1_737_4650 (.A1(\out_bs[4] [5]), .A2(n_1_737_4101), .ZN(
      n_1_737_4100));
   NOR2_X1 i_1_737_4651 (.A1(n_1_737_5623), .A2(n_1_737_4643), .ZN(n_1_737_4101));
   INV_X1 i_1_737_4652 (.A(n_1_737_4103), .ZN(n_1_737_4102));
   OAI21_X1 i_1_737_4653 (.A(n_1_737_4105), .B1(n_1_737_5236), .B2(n_1_737_4104), 
      .ZN(n_1_737_4103));
   NOR2_X1 i_1_737_4654 (.A1(n_1_737_5275), .A2(n_1_737_4106), .ZN(n_1_737_4104));
   NAND2_X1 i_1_737_4655 (.A1(n_1_737_5275), .A2(n_1_737_4106), .ZN(n_1_737_4105));
   NAND2_X1 i_1_737_4656 (.A1(n_1_737_5651), .A2(n_1_737_4107), .ZN(n_1_737_4106));
   NOR2_X1 i_1_737_4657 (.A1(\out_bs[2] [5]), .A2(n_1_737_4108), .ZN(
      n_1_737_4107));
   NOR2_X1 i_1_737_4658 (.A1(n_1_737_5649), .A2(n_1_737_4638), .ZN(n_1_737_4108));
   AOI22_X1 i_1_737_4659 (.A1(n_1_737_5216), .A2(n_1_737_4111), .B1(n_1_737_5189), 
      .B2(n_1_737_4110), .ZN(n_1_737_4109));
   NAND3_X1 i_1_737_4660 (.A1(n_1_737_5638), .A2(n_1_737_4112), .A3(n_1_737_5215), 
      .ZN(n_1_737_4110));
   NAND2_X1 i_1_737_4661 (.A1(n_1_737_5638), .A2(n_1_737_4112), .ZN(n_1_737_4111));
   NOR2_X1 i_1_737_4662 (.A1(\out_bs[3] [5]), .A2(n_1_737_4113), .ZN(
      n_1_737_4112));
   NOR2_X1 i_1_737_4663 (.A1(n_1_737_5636), .A2(n_1_737_4622), .ZN(n_1_737_4113));
   INV_X1 i_1_737_4664 (.A(n_1_737_4115), .ZN(n_1_737_4114));
   OAI21_X1 i_1_737_4665 (.A(n_1_737_4116), .B1(n_1_737_5320), .B2(n_1_737_5298), 
      .ZN(n_1_737_4115));
   OAI22_X1 i_1_737_4666 (.A1(n_1_737_5284), .A2(n_1_737_4118), .B1(n_1_737_5321), 
      .B2(n_1_737_5297), .ZN(n_1_737_4116));
   NOR2_X1 i_1_737_4667 (.A1(\out_bs[1] [5]), .A2(n_1_737_4118), .ZN(
      n_1_737_4117));
   NOR2_X1 i_1_737_4668 (.A1(n_1_737_5662), .A2(n_1_737_4631), .ZN(n_1_737_4118));
   NOR2_X1 i_1_737_4669 (.A1(n_1_737_300), .A2(n_1_737_5155), .ZN(n_550));
   AOI211_X1 i_1_737_4670 (.A(n_1_737_299), .B(n_1_737_5167), .C1(n_1_737_5182), 
      .C2(n_1_737_4119), .ZN(n_551));
   OAI211_X1 i_1_737_4671 (.A(n_1_737_5182), .B(n_1_737_4119), .C1(n_1_737_299), 
      .C2(n_1_737_5167), .ZN(n_552));
   INV_X1 i_1_737_4672 (.A(n_1_737_4120), .ZN(n_1_737_4119));
   NOR2_X1 i_1_737_4673 (.A1(n_1_737_5610), .A2(n_1_737_4645), .ZN(n_1_737_4120));
   NAND3_X1 i_1_737_4674 (.A1(n_1_737_4139), .A2(n_1_737_4128), .A3(n_1_737_4121), 
      .ZN(n_553));
   NOR3_X1 i_1_737_4675 (.A1(n_1_737_4145), .A2(n_1_737_4123), .A3(n_1_737_4134), 
      .ZN(n_1_737_4121));
   INV_X1 i_1_737_4676 (.A(n_1_737_4123), .ZN(n_1_737_4122));
   OAI21_X1 i_1_737_4677 (.A(n_1_737_4124), .B1(n_1_737_5298), .B2(n_1_737_4125), 
      .ZN(n_1_737_4123));
   OAI21_X1 i_1_737_4678 (.A(n_1_737_4127), .B1(n_1_737_5297), .B2(n_1_737_4126), 
      .ZN(n_1_737_4124));
   INV_X1 i_1_737_4679 (.A(n_1_737_4126), .ZN(n_1_737_4125));
   NOR2_X1 i_1_737_4680 (.A1(n_1_737_295), .A2(n_1_737_5320), .ZN(n_1_737_4126));
   OAI21_X1 i_1_737_4681 (.A(n_1_737_5285), .B1(n_1_737_5662), .B2(n_1_737_4653), 
      .ZN(n_1_737_4127));
   AOI22_X1 i_1_737_4682 (.A1(n_1_737_4133), .A2(n_1_737_4130), .B1(n_1_737_5189), 
      .B2(n_1_737_4129), .ZN(n_1_737_4128));
   OAI21_X1 i_1_737_4683 (.A(n_1_737_4131), .B1(n_1_737_297), .B2(n_1_737_5215), 
      .ZN(n_1_737_4129));
   INV_X1 i_1_737_4684 (.A(n_1_737_4131), .ZN(n_1_737_4130));
   NOR2_X1 i_1_737_4685 (.A1(n_1_737_5221), .A2(n_1_737_4132), .ZN(n_1_737_4131));
   NOR2_X1 i_1_737_4686 (.A1(n_1_737_5636), .A2(n_1_737_4658), .ZN(n_1_737_4132));
   NOR2_X1 i_1_737_4687 (.A1(n_1_737_297), .A2(n_1_737_5215), .ZN(n_1_737_4133));
   OAI21_X1 i_1_737_4688 (.A(n_1_737_4135), .B1(n_1_737_5337), .B2(n_1_737_4136), 
      .ZN(n_1_737_4134));
   OAI22_X1 i_1_737_4689 (.A1(n_1_737_5083), .A2(n_1_737_4138), .B1(n_1_737_5336), 
      .B2(n_1_737_4137), .ZN(n_1_737_4135));
   INV_X1 i_1_737_4690 (.A(n_1_737_4137), .ZN(n_1_737_4136));
   NOR2_X1 i_1_737_4691 (.A1(n_1_737_294), .A2(n_1_737_5358), .ZN(n_1_737_4137));
   NOR2_X1 i_1_737_4692 (.A1(n_1_737_5669), .A2(n_1_737_4669), .ZN(n_1_737_4138));
   OAI22_X1 i_1_737_4693 (.A1(n_1_737_4144), .A2(n_1_737_4140), .B1(n_1_737_5235), 
      .B2(n_1_737_4141), .ZN(n_1_737_4139));
   AND2_X1 i_1_737_4694 (.A1(n_1_737_5235), .A2(n_1_737_4141), .ZN(n_1_737_4140));
   NAND2_X1 i_1_737_4695 (.A1(n_1_737_5651), .A2(n_1_737_4142), .ZN(n_1_737_4141));
   NOR2_X1 i_1_737_4696 (.A1(\out_bs[2] [5]), .A2(n_1_737_4143), .ZN(
      n_1_737_4142));
   NOR2_X1 i_1_737_4697 (.A1(n_1_737_5649), .A2(n_1_737_4664), .ZN(n_1_737_4143));
   NOR2_X1 i_1_737_4698 (.A1(n_1_737_296), .A2(n_1_737_5274), .ZN(n_1_737_4144));
   INV_X1 i_1_737_4699 (.A(n_1_737_4146), .ZN(n_1_737_4145));
   OAI22_X1 i_1_737_4700 (.A1(n_1_737_4151), .A2(n_1_737_4147), .B1(n_1_737_5365), 
      .B2(n_1_737_4148), .ZN(n_1_737_4146));
   AND2_X1 i_1_737_4701 (.A1(n_1_737_5365), .A2(n_1_737_4148), .ZN(n_1_737_4147));
   NAND2_X1 i_1_737_4702 (.A1(n_1_737_5625), .A2(n_1_737_4149), .ZN(n_1_737_4148));
   NOR2_X1 i_1_737_4703 (.A1(\out_bs[4] [5]), .A2(n_1_737_4150), .ZN(
      n_1_737_4149));
   NOR2_X1 i_1_737_4704 (.A1(n_1_737_5623), .A2(n_1_737_4676), .ZN(n_1_737_4150));
   NOR2_X1 i_1_737_4705 (.A1(n_1_737_298), .A2(n_1_737_5386), .ZN(n_1_737_4151));
   NOR2_X1 i_1_737_4706 (.A1(n_1_737_293), .A2(n_1_737_5155), .ZN(n_554));
   NOR3_X1 i_1_737_4707 (.A1(n_1_737_292), .A2(n_1_737_5167), .A3(n_1_737_4152), 
      .ZN(n_555));
   OAI21_X1 i_1_737_4708 (.A(n_1_737_4152), .B1(n_1_737_292), .B2(n_1_737_5167), 
      .ZN(n_556));
   NOR2_X1 i_1_737_4709 (.A1(n_1_737_5181), .A2(n_1_737_4153), .ZN(n_1_737_4152));
   NOR2_X1 i_1_737_4710 (.A1(n_1_737_5610), .A2(n_1_737_4678), .ZN(n_1_737_4153));
   NAND3_X1 i_1_737_4711 (.A1(n_1_737_4173), .A2(n_1_737_4160), .A3(n_1_737_4154), 
      .ZN(n_557));
   NOR3_X1 i_1_737_4712 (.A1(n_1_737_4180), .A2(n_1_737_4167), .A3(n_1_737_4155), 
      .ZN(n_1_737_4154));
   OAI21_X1 i_1_737_4713 (.A(n_1_737_4156), .B1(n_1_737_5337), .B2(n_1_737_4157), 
      .ZN(n_1_737_4155));
   OAI22_X1 i_1_737_4714 (.A1(n_1_737_5083), .A2(n_1_737_4159), .B1(n_1_737_5336), 
      .B2(n_1_737_4158), .ZN(n_1_737_4156));
   INV_X1 i_1_737_4715 (.A(n_1_737_4158), .ZN(n_1_737_4157));
   NOR2_X1 i_1_737_4716 (.A1(n_1_737_287), .A2(n_1_737_5358), .ZN(n_1_737_4158));
   NOR2_X1 i_1_737_4717 (.A1(n_1_737_5669), .A2(n_1_737_4685), .ZN(n_1_737_4159));
   OAI22_X1 i_1_737_4718 (.A1(n_1_737_4165), .A2(n_1_737_4161), .B1(n_1_737_5189), 
      .B2(n_1_737_4162), .ZN(n_1_737_4160));
   AND2_X1 i_1_737_4719 (.A1(n_1_737_5189), .A2(n_1_737_4162), .ZN(n_1_737_4161));
   NAND2_X1 i_1_737_4720 (.A1(n_1_737_5638), .A2(n_1_737_4163), .ZN(n_1_737_4162));
   NOR2_X1 i_1_737_4721 (.A1(\out_bs[3] [5]), .A2(n_1_737_4164), .ZN(
      n_1_737_4163));
   NOR2_X1 i_1_737_4722 (.A1(n_1_737_5636), .A2(n_1_737_4691), .ZN(n_1_737_4164));
   NOR2_X1 i_1_737_4723 (.A1(n_1_737_290), .A2(n_1_737_5215), .ZN(n_1_737_4165));
   INV_X1 i_1_737_4724 (.A(n_1_737_4167), .ZN(n_1_737_4166));
   OAI21_X1 i_1_737_4725 (.A(n_1_737_4168), .B1(n_1_737_5298), .B2(n_1_737_4169), 
      .ZN(n_1_737_4167));
   OAI22_X1 i_1_737_4726 (.A1(n_1_737_5284), .A2(n_1_737_4172), .B1(n_1_737_5297), 
      .B2(n_1_737_4170), .ZN(n_1_737_4168));
   INV_X1 i_1_737_4727 (.A(n_1_737_4170), .ZN(n_1_737_4169));
   NOR2_X1 i_1_737_4728 (.A1(n_1_737_288), .A2(n_1_737_5320), .ZN(n_1_737_4170));
   NOR2_X1 i_1_737_4729 (.A1(\out_bs[1] [5]), .A2(n_1_737_4172), .ZN(
      n_1_737_4171));
   NOR2_X1 i_1_737_4730 (.A1(n_1_737_5662), .A2(n_1_737_4698), .ZN(n_1_737_4172));
   AOI21_X1 i_1_737_4731 (.A(n_1_737_4174), .B1(n_1_737_5235), .B2(n_1_737_4176), 
      .ZN(n_1_737_4173));
   AOI22_X1 i_1_737_4732 (.A1(n_1_737_5651), .A2(n_1_737_4177), .B1(n_1_737_5236), 
      .B2(n_1_737_4175), .ZN(n_1_737_4174));
   INV_X1 i_1_737_4733 (.A(n_1_737_4176), .ZN(n_1_737_4175));
   NOR2_X1 i_1_737_4734 (.A1(n_1_737_289), .A2(n_1_737_5274), .ZN(n_1_737_4176));
   NOR2_X1 i_1_737_4735 (.A1(\out_bs[2] [5]), .A2(n_1_737_4178), .ZN(
      n_1_737_4177));
   NOR2_X1 i_1_737_4736 (.A1(n_1_737_5649), .A2(n_1_737_4706), .ZN(n_1_737_4178));
   INV_X1 i_1_737_4737 (.A(n_1_737_4180), .ZN(n_1_737_4179));
   OAI21_X1 i_1_737_4738 (.A(n_1_737_4181), .B1(n_1_737_5366), .B2(n_1_737_4182), 
      .ZN(n_1_737_4180));
   OAI21_X1 i_1_737_4739 (.A(n_1_737_4184), .B1(n_1_737_5365), .B2(n_1_737_4183), 
      .ZN(n_1_737_4181));
   INV_X1 i_1_737_4740 (.A(n_1_737_4183), .ZN(n_1_737_4182));
   NOR2_X1 i_1_737_4741 (.A1(n_1_737_291), .A2(n_1_737_5386), .ZN(n_1_737_4183));
   OAI21_X1 i_1_737_4742 (.A(n_1_737_5393), .B1(n_1_737_5623), .B2(n_1_737_4714), 
      .ZN(n_1_737_4184));
   NOR2_X1 i_1_737_4743 (.A1(n_1_737_286), .A2(n_1_737_5155), .ZN(n_558));
   NOR3_X1 i_1_737_4744 (.A1(n_1_737_285), .A2(n_1_737_5167), .A3(n_1_737_4208), 
      .ZN(n_559));
   OAI21_X1 i_1_737_4745 (.A(n_1_737_4208), .B1(n_1_737_285), .B2(n_1_737_5167), 
      .ZN(n_560));
   NAND4_X1 i_1_737_4746 (.A1(n_1_737_4200), .A2(n_1_737_4199), .A3(n_1_737_4185), 
      .A4(n_1_737_4202), .ZN(n_561));
   NOR3_X1 i_1_737_4747 (.A1(n_1_737_4191), .A2(n_1_737_4186), .A3(n_1_737_4195), 
      .ZN(n_1_737_4185));
   INV_X1 i_1_737_4748 (.A(n_1_737_4187), .ZN(n_1_737_4186));
   OAI21_X1 i_1_737_4749 (.A(n_1_737_4188), .B1(n_1_737_5297), .B2(n_1_737_4190), 
      .ZN(n_1_737_4187));
   OAI211_X1 i_1_737_4750 (.A(n_1_737_5285), .B(n_1_737_4218), .C1(n_1_737_5298), 
      .C2(n_1_737_4189), .ZN(n_1_737_4188));
   INV_X1 i_1_737_4751 (.A(n_1_737_4190), .ZN(n_1_737_4189));
   NOR2_X1 i_1_737_4752 (.A1(n_1_737_281), .A2(n_1_737_5320), .ZN(n_1_737_4190));
   OAI21_X1 i_1_737_4753 (.A(n_1_737_4193), .B1(n_1_737_5190), .B2(n_1_737_4192), 
      .ZN(n_1_737_4191));
   NOR2_X1 i_1_737_4754 (.A1(n_1_737_4224), .A2(n_1_737_4194), .ZN(n_1_737_4192));
   NAND2_X1 i_1_737_4755 (.A1(n_1_737_4224), .A2(n_1_737_4194), .ZN(n_1_737_4193));
   NOR2_X1 i_1_737_4756 (.A1(n_1_737_283), .A2(n_1_737_5215), .ZN(n_1_737_4194));
   INV_X1 i_1_737_4757 (.A(n_1_737_4196), .ZN(n_1_737_4195));
   AOI22_X1 i_1_737_4758 (.A1(n_1_737_4233), .A2(n_1_737_4198), .B1(n_1_737_5235), 
      .B2(n_1_737_4197), .ZN(n_1_737_4196));
   OR2_X1 i_1_737_4759 (.A1(n_1_737_4233), .A2(n_1_737_4198), .ZN(n_1_737_4197));
   NOR2_X1 i_1_737_4760 (.A1(n_1_737_282), .A2(n_1_737_5274), .ZN(n_1_737_4198));
   NAND2_X1 i_1_737_4761 (.A1(n_1_737_5336), .A2(n_1_737_4201), .ZN(n_1_737_4199));
   OAI22_X1 i_1_737_4762 (.A1(n_1_737_5083), .A2(n_1_737_4243), .B1(n_1_737_5336), 
      .B2(n_1_737_4201), .ZN(n_1_737_4200));
   NOR2_X1 i_1_737_4763 (.A1(n_1_737_280), .A2(n_1_737_5358), .ZN(n_1_737_4201));
   OAI22_X1 i_1_737_4764 (.A1(n_1_737_4251), .A2(n_1_737_4203), .B1(n_1_737_5365), 
      .B2(n_1_737_4204), .ZN(n_1_737_4202));
   AND2_X1 i_1_737_4765 (.A1(n_1_737_5365), .A2(n_1_737_4204), .ZN(n_1_737_4203));
   NOR2_X1 i_1_737_4766 (.A1(n_1_737_284), .A2(n_1_737_5386), .ZN(n_1_737_4204));
   NOR2_X1 i_1_737_4767 (.A1(n_1_737_279), .A2(n_1_737_5155), .ZN(n_562));
   NOR3_X1 i_1_737_4768 (.A1(n_1_737_278), .A2(n_1_737_5167), .A3(n_1_737_4205), 
      .ZN(n_563));
   OAI21_X1 i_1_737_4769 (.A(n_1_737_4205), .B1(n_1_737_278), .B2(n_1_737_5167), 
      .ZN(n_564));
   NOR2_X1 i_1_737_4770 (.A1(n_1_737_5181), .A2(n_1_737_4206), .ZN(n_1_737_4205));
   INV_X1 i_1_737_4771 (.A(n_1_737_4207), .ZN(n_1_737_4206));
   AOI21_X1 i_1_737_4772 (.A(n_1_737_4209), .B1(n_1_737_5022), .B2(n_1_737_4404), 
      .ZN(n_1_737_4207));
   NOR2_X1 i_1_737_4773 (.A1(n_1_737_5181), .A2(n_1_737_4209), .ZN(n_1_737_4208));
   NOR2_X1 i_1_737_4774 (.A1(n_1_737_5608), .A2(n_1_737_4403), .ZN(n_1_737_4209));
   NAND3_X1 i_1_737_4775 (.A1(n_1_737_4227), .A2(n_1_737_4219), .A3(n_1_737_4210), 
      .ZN(n_565));
   NOR3_X1 i_1_737_4776 (.A1(n_1_737_4245), .A2(n_1_737_4212), .A3(n_1_737_4236), 
      .ZN(n_1_737_4210));
   INV_X1 i_1_737_4777 (.A(n_1_737_4212), .ZN(n_1_737_4211));
   OAI21_X1 i_1_737_4778 (.A(n_1_737_4213), .B1(n_1_737_5298), .B2(n_1_737_4214), 
      .ZN(n_1_737_4212));
   OAI22_X1 i_1_737_4779 (.A1(n_1_737_5284), .A2(n_1_737_4217), .B1(n_1_737_5297), 
      .B2(n_1_737_4215), .ZN(n_1_737_4213));
   INV_X1 i_1_737_4780 (.A(n_1_737_4215), .ZN(n_1_737_4214));
   NOR2_X1 i_1_737_4781 (.A1(n_1_737_274), .A2(n_1_737_5320), .ZN(n_1_737_4215));
   INV_X1 i_1_737_4782 (.A(n_1_737_4217), .ZN(n_1_737_4216));
   OAI21_X1 i_1_737_4783 (.A(n_1_737_4218), .B1(n_1_737_5048), .B2(n_1_737_4450), 
      .ZN(n_1_737_4217));
   NAND2_X1 i_1_737_4784 (.A1(\out_bs[1] [4]), .A2(n_1_737_4753), .ZN(
      n_1_737_4218));
   AOI22_X1 i_1_737_4785 (.A1(n_1_737_4226), .A2(n_1_737_4221), .B1(n_1_737_5189), 
      .B2(n_1_737_4220), .ZN(n_1_737_4219));
   OAI21_X1 i_1_737_4786 (.A(n_1_737_4222), .B1(n_1_737_276), .B2(n_1_737_5215), 
      .ZN(n_1_737_4220));
   INV_X1 i_1_737_4787 (.A(n_1_737_4222), .ZN(n_1_737_4221));
   NOR2_X1 i_1_737_4788 (.A1(n_1_737_5221), .A2(n_1_737_4223), .ZN(n_1_737_4222));
   OAI21_X1 i_1_737_4789 (.A(n_1_737_4225), .B1(n_1_737_5039), .B2(n_1_737_4426), 
      .ZN(n_1_737_4223));
   NAND2_X1 i_1_737_4790 (.A1(n_1_737_5222), .A2(n_1_737_4225), .ZN(n_1_737_4224));
   NAND2_X1 i_1_737_4791 (.A1(\out_bs[3] [4]), .A2(n_1_737_4763), .ZN(
      n_1_737_4225));
   NOR2_X1 i_1_737_4792 (.A1(n_1_737_276), .A2(n_1_737_5215), .ZN(n_1_737_4226));
   OAI22_X1 i_1_737_4793 (.A1(n_1_737_4235), .A2(n_1_737_4228), .B1(n_1_737_5235), 
      .B2(n_1_737_4229), .ZN(n_1_737_4227));
   NOR2_X1 i_1_737_4794 (.A1(n_1_737_5236), .A2(n_1_737_4230), .ZN(n_1_737_4228));
   INV_X1 i_1_737_4795 (.A(n_1_737_4230), .ZN(n_1_737_4229));
   NOR2_X1 i_1_737_4796 (.A1(n_1_737_5252), .A2(n_1_737_4232), .ZN(n_1_737_4230));
   INV_X1 i_1_737_4797 (.A(n_1_737_4232), .ZN(n_1_737_4231));
   OAI21_X1 i_1_737_4798 (.A(n_1_737_4234), .B1(n_1_737_5056), .B2(n_1_737_4415), 
      .ZN(n_1_737_4232));
   NAND2_X1 i_1_737_4799 (.A1(n_1_737_5253), .A2(n_1_737_4234), .ZN(n_1_737_4233));
   NAND2_X1 i_1_737_4800 (.A1(\out_bs[2] [4]), .A2(n_1_737_4772), .ZN(
      n_1_737_4234));
   NOR2_X1 i_1_737_4801 (.A1(n_1_737_275), .A2(n_1_737_5274), .ZN(n_1_737_4235));
   OAI21_X1 i_1_737_4802 (.A(n_1_737_4237), .B1(n_1_737_5337), .B2(n_1_737_4238), 
      .ZN(n_1_737_4236));
   OAI22_X1 i_1_737_4803 (.A1(n_1_737_5083), .A2(n_1_737_4241), .B1(n_1_737_5336), 
      .B2(n_1_737_4239), .ZN(n_1_737_4237));
   INV_X1 i_1_737_4804 (.A(n_1_737_4239), .ZN(n_1_737_4238));
   NOR2_X1 i_1_737_4805 (.A1(n_1_737_273), .A2(n_1_737_5358), .ZN(n_1_737_4239));
   NOR2_X1 i_1_737_4806 (.A1(\out_bs[0] [5]), .A2(n_1_737_4241), .ZN(
      n_1_737_4240));
   INV_X1 i_1_737_4807 (.A(n_1_737_4242), .ZN(n_1_737_4241));
   AOI21_X1 i_1_737_4808 (.A(n_1_737_4243), .B1(n_1_737_5030), .B2(n_1_737_4438), 
      .ZN(n_1_737_4242));
   NOR2_X1 i_1_737_4809 (.A1(n_1_737_5667), .A2(n_1_737_4437), .ZN(n_1_737_4243));
   INV_X1 i_1_737_4810 (.A(n_1_737_4245), .ZN(n_1_737_4244));
   OAI21_X1 i_1_737_4811 (.A(n_1_737_4246), .B1(n_1_737_5366), .B2(n_1_737_4247), 
      .ZN(n_1_737_4245));
   OAI22_X1 i_1_737_4812 (.A1(n_1_737_5392), .A2(n_1_737_4249), .B1(n_1_737_5365), 
      .B2(n_1_737_4248), .ZN(n_1_737_4246));
   INV_X1 i_1_737_4813 (.A(n_1_737_4248), .ZN(n_1_737_4247));
   NOR2_X1 i_1_737_4814 (.A1(n_1_737_277), .A2(n_1_737_5386), .ZN(n_1_737_4248));
   INV_X1 i_1_737_4815 (.A(n_1_737_4250), .ZN(n_1_737_4249));
   AOI21_X1 i_1_737_4816 (.A(n_1_737_4253), .B1(n_1_737_5065), .B2(n_1_737_4462), 
      .ZN(n_1_737_4250));
   NAND2_X1 i_1_737_4817 (.A1(n_1_737_5625), .A2(n_1_737_4252), .ZN(n_1_737_4251));
   NOR2_X1 i_1_737_4818 (.A1(\out_bs[4] [5]), .A2(n_1_737_4253), .ZN(
      n_1_737_4252));
   NOR3_X1 i_1_737_4819 (.A1(n_1_737_5623), .A2(n_1_737_5622), .A3(n_1_737_5621), 
      .ZN(n_1_737_4253));
   NOR2_X1 i_1_737_4820 (.A1(n_1_737_272), .A2(n_1_737_5155), .ZN(n_566));
   AOI211_X1 i_1_737_4821 (.A(n_1_737_271), .B(n_1_737_5167), .C1(n_1_737_5182), 
      .C2(n_1_737_4254), .ZN(n_567));
   OAI211_X1 i_1_737_4822 (.A(n_1_737_5182), .B(n_1_737_4254), .C1(n_1_737_271), 
      .C2(n_1_737_5167), .ZN(n_568));
   INV_X1 i_1_737_4823 (.A(n_1_737_4255), .ZN(n_1_737_4254));
   NOR2_X1 i_1_737_4824 (.A1(n_1_737_5610), .A2(n_1_737_4813), .ZN(n_1_737_4255));
   NAND4_X1 i_1_737_4825 (.A1(n_1_737_4259), .A2(n_1_737_4256), .A3(n_1_737_4274), 
      .A4(n_1_737_4281), .ZN(n_569));
   AOI211_X1 i_1_737_4826 (.A(n_1_737_4257), .B(n_1_737_4268), .C1(n_1_737_5336), 
      .C2(n_1_737_4265), .ZN(n_1_737_4256));
   INV_X1 i_1_737_4827 (.A(n_1_737_4258), .ZN(n_1_737_4257));
   OAI22_X1 i_1_737_4828 (.A1(n_1_737_5083), .A2(n_1_737_4266), .B1(n_1_737_5336), 
      .B2(n_1_737_4265), .ZN(n_1_737_4258));
   AOI22_X1 i_1_737_4829 (.A1(n_1_737_4264), .A2(n_1_737_4261), .B1(n_1_737_5189), 
      .B2(n_1_737_4260), .ZN(n_1_737_4259));
   OAI21_X1 i_1_737_4830 (.A(n_1_737_4262), .B1(n_1_737_269), .B2(n_1_737_5215), 
      .ZN(n_1_737_4260));
   INV_X1 i_1_737_4831 (.A(n_1_737_4262), .ZN(n_1_737_4261));
   NOR2_X1 i_1_737_4832 (.A1(n_1_737_5221), .A2(n_1_737_4263), .ZN(n_1_737_4262));
   NOR2_X1 i_1_737_4833 (.A1(n_1_737_5636), .A2(n_1_737_4834), .ZN(n_1_737_4263));
   NOR2_X1 i_1_737_4834 (.A1(n_1_737_269), .A2(n_1_737_5215), .ZN(n_1_737_4264));
   NOR2_X1 i_1_737_4835 (.A1(n_1_737_266), .A2(n_1_737_5358), .ZN(n_1_737_4265));
   NOR2_X1 i_1_737_4836 (.A1(n_1_737_5669), .A2(n_1_737_4822), .ZN(n_1_737_4266));
   INV_X1 i_1_737_4837 (.A(n_1_737_4268), .ZN(n_1_737_4267));
   OAI21_X1 i_1_737_4838 (.A(n_1_737_4269), .B1(n_1_737_5298), .B2(n_1_737_4270), 
      .ZN(n_1_737_4268));
   OAI22_X1 i_1_737_4839 (.A1(n_1_737_5284), .A2(n_1_737_4273), .B1(n_1_737_5297), 
      .B2(n_1_737_4271), .ZN(n_1_737_4269));
   INV_X1 i_1_737_4840 (.A(n_1_737_4271), .ZN(n_1_737_4270));
   NOR2_X1 i_1_737_4841 (.A1(n_1_737_267), .A2(n_1_737_5320), .ZN(n_1_737_4271));
   NOR2_X1 i_1_737_4842 (.A1(\out_bs[1] [5]), .A2(n_1_737_4273), .ZN(
      n_1_737_4272));
   NOR2_X1 i_1_737_4843 (.A1(n_1_737_5662), .A2(n_1_737_4844), .ZN(n_1_737_4273));
   OAI22_X1 i_1_737_4844 (.A1(n_1_737_4279), .A2(n_1_737_4275), .B1(n_1_737_5235), 
      .B2(n_1_737_4276), .ZN(n_1_737_4274));
   AND2_X1 i_1_737_4845 (.A1(n_1_737_5235), .A2(n_1_737_4276), .ZN(n_1_737_4275));
   NAND2_X1 i_1_737_4846 (.A1(n_1_737_5651), .A2(n_1_737_4277), .ZN(n_1_737_4276));
   NOR2_X1 i_1_737_4847 (.A1(\out_bs[2] [5]), .A2(n_1_737_4278), .ZN(
      n_1_737_4277));
   NOR2_X1 i_1_737_4848 (.A1(n_1_737_5649), .A2(n_1_737_4853), .ZN(n_1_737_4278));
   NOR2_X1 i_1_737_4849 (.A1(n_1_737_268), .A2(n_1_737_5274), .ZN(n_1_737_4279));
   INV_X1 i_1_737_4850 (.A(n_1_737_4281), .ZN(n_1_737_4280));
   OAI21_X1 i_1_737_4851 (.A(n_1_737_4282), .B1(n_1_737_5365), .B2(n_1_737_4283), 
      .ZN(n_1_737_4281));
   OAI22_X1 i_1_737_4852 (.A1(n_1_737_270), .A2(n_1_737_5386), .B1(n_1_737_5366), 
      .B2(n_1_737_4284), .ZN(n_1_737_4282));
   INV_X1 i_1_737_4853 (.A(n_1_737_4284), .ZN(n_1_737_4283));
   NOR2_X1 i_1_737_4854 (.A1(n_1_737_5392), .A2(n_1_737_4285), .ZN(n_1_737_4284));
   NOR2_X1 i_1_737_4855 (.A1(n_1_737_5623), .A2(n_1_737_4862), .ZN(n_1_737_4285));
   NOR2_X1 i_1_737_4856 (.A1(n_1_737_265), .A2(n_1_737_5155), .ZN(n_570));
   NOR3_X1 i_1_737_4857 (.A1(n_1_737_264), .A2(n_1_737_5167), .A3(n_1_737_4286), 
      .ZN(n_571));
   OAI21_X1 i_1_737_4858 (.A(n_1_737_4286), .B1(n_1_737_264), .B2(n_1_737_5167), 
      .ZN(n_572));
   AOI21_X1 i_1_737_4859 (.A(n_1_737_5181), .B1(n_848), .B2(n_1_737_4810), 
      .ZN(n_1_737_4286));
   NAND3_X1 i_1_737_4860 (.A1(n_1_737_4304), .A2(n_1_737_4293), .A3(n_1_737_4287), 
      .ZN(n_573));
   NOR3_X1 i_1_737_4861 (.A1(n_1_737_4310), .A2(n_1_737_4299), .A3(n_1_737_4288), 
      .ZN(n_1_737_4287));
   OAI21_X1 i_1_737_4862 (.A(n_1_737_4289), .B1(n_1_737_5337), .B2(n_1_737_4290), 
      .ZN(n_1_737_4288));
   OAI22_X1 i_1_737_4863 (.A1(n_1_737_5083), .A2(n_1_737_4292), .B1(n_1_737_5336), 
      .B2(n_1_737_4291), .ZN(n_1_737_4289));
   INV_X1 i_1_737_4864 (.A(n_1_737_4291), .ZN(n_1_737_4290));
   NOR2_X1 i_1_737_4865 (.A1(n_1_737_259), .A2(n_1_737_5358), .ZN(n_1_737_4291));
   NOR2_X1 i_1_737_4866 (.A1(n_1_737_5669), .A2(n_1_737_4820), .ZN(n_1_737_4292));
   AOI21_X1 i_1_737_4867 (.A(n_1_737_4294), .B1(n_1_737_5235), .B2(n_1_737_4296), 
      .ZN(n_1_737_4293));
   INV_X1 i_1_737_4868 (.A(n_1_737_4295), .ZN(n_1_737_4294));
   OAI22_X1 i_1_737_4869 (.A1(n_1_737_5252), .A2(n_1_737_4297), .B1(n_1_737_5235), 
      .B2(n_1_737_4296), .ZN(n_1_737_4295));
   NOR2_X1 i_1_737_4870 (.A1(n_1_737_261), .A2(n_1_737_5274), .ZN(n_1_737_4296));
   NOR2_X1 i_1_737_4871 (.A1(n_1_737_5649), .A2(n_1_737_4851), .ZN(n_1_737_4297));
   INV_X1 i_1_737_4872 (.A(n_1_737_4299), .ZN(n_1_737_4298));
   OAI21_X1 i_1_737_4873 (.A(n_1_737_4300), .B1(n_1_737_5298), .B2(n_1_737_4301), 
      .ZN(n_1_737_4299));
   OAI22_X1 i_1_737_4874 (.A1(n_1_737_5284), .A2(n_1_737_4303), .B1(n_1_737_5297), 
      .B2(n_1_737_4302), .ZN(n_1_737_4300));
   INV_X1 i_1_737_4875 (.A(n_1_737_4302), .ZN(n_1_737_4301));
   NOR2_X1 i_1_737_4876 (.A1(n_1_737_260), .A2(n_1_737_5320), .ZN(n_1_737_4302));
   NOR2_X1 i_1_737_4877 (.A1(n_1_737_5662), .A2(n_1_737_4840), .ZN(n_1_737_4303));
   AOI21_X1 i_1_737_4878 (.A(n_1_737_4305), .B1(n_1_737_5189), .B2(n_1_737_4307), 
      .ZN(n_1_737_4304));
   INV_X1 i_1_737_4879 (.A(n_1_737_4306), .ZN(n_1_737_4305));
   OAI22_X1 i_1_737_4880 (.A1(n_1_737_5221), .A2(n_1_737_4308), .B1(n_1_737_5189), 
      .B2(n_1_737_4307), .ZN(n_1_737_4306));
   NOR2_X1 i_1_737_4881 (.A1(n_1_737_262), .A2(n_1_737_5215), .ZN(n_1_737_4307));
   NOR2_X1 i_1_737_4882 (.A1(n_1_737_5636), .A2(n_1_737_4830), .ZN(n_1_737_4308));
   INV_X1 i_1_737_4883 (.A(n_1_737_4310), .ZN(n_1_737_4309));
   OAI21_X1 i_1_737_4884 (.A(n_1_737_4311), .B1(n_1_737_5366), .B2(n_1_737_4312), 
      .ZN(n_1_737_4310));
   OAI22_X1 i_1_737_4885 (.A1(n_1_737_5392), .A2(n_1_737_4314), .B1(n_1_737_5365), 
      .B2(n_1_737_4313), .ZN(n_1_737_4311));
   INV_X1 i_1_737_4886 (.A(n_1_737_4313), .ZN(n_1_737_4312));
   NOR2_X1 i_1_737_4887 (.A1(n_1_737_263), .A2(n_1_737_5386), .ZN(n_1_737_4313));
   NOR2_X1 i_1_737_4888 (.A1(n_1_737_5623), .A2(n_1_737_4861), .ZN(n_1_737_4314));
   NOR2_X1 i_1_737_4889 (.A1(n_1_737_258), .A2(n_1_737_5155), .ZN(n_574));
   NOR3_X1 i_1_737_4890 (.A1(n_1_737_257), .A2(n_1_737_5167), .A3(n_1_737_4402), 
      .ZN(n_575));
   OAI21_X1 i_1_737_4891 (.A(n_1_737_4402), .B1(n_1_737_257), .B2(n_1_737_5167), 
      .ZN(n_576));
   NAND3_X1 i_1_737_4892 (.A1(n_1_737_4327), .A2(n_1_737_4324), .A3(n_1_737_4315), 
      .ZN(n_577));
   NOR3_X1 i_1_737_4893 (.A1(n_1_737_4330), .A2(n_1_737_4320), .A3(n_1_737_4316), 
      .ZN(n_1_737_4315));
   OAI21_X1 i_1_737_4894 (.A(n_1_737_4317), .B1(n_1_737_5337), .B2(n_1_737_4318), 
      .ZN(n_1_737_4316));
   OAI21_X1 i_1_737_4895 (.A(n_1_737_4434), .B1(n_1_737_5336), .B2(n_1_737_4319), 
      .ZN(n_1_737_4317));
   INV_X1 i_1_737_4896 (.A(n_1_737_4319), .ZN(n_1_737_4318));
   NOR2_X1 i_1_737_4897 (.A1(n_1_737_252), .A2(n_1_737_5358), .ZN(n_1_737_4319));
   INV_X1 i_1_737_4898 (.A(n_1_737_4321), .ZN(n_1_737_4320));
   AOI22_X1 i_1_737_4899 (.A1(n_1_737_4457), .A2(n_1_737_4323), .B1(n_1_737_5365), 
      .B2(n_1_737_4322), .ZN(n_1_737_4321));
   OAI21_X1 i_1_737_4900 (.A(n_1_737_4458), .B1(n_1_737_256), .B2(n_1_737_5386), 
      .ZN(n_1_737_4322));
   NOR2_X1 i_1_737_4901 (.A1(n_1_737_256), .A2(n_1_737_5386), .ZN(n_1_737_4323));
   AOI22_X1 i_1_737_4902 (.A1(n_1_737_4409), .A2(n_1_737_4326), .B1(n_1_737_5235), 
      .B2(n_1_737_4325), .ZN(n_1_737_4324));
   OAI21_X1 i_1_737_4903 (.A(n_1_737_4410), .B1(n_1_737_254), .B2(n_1_737_5274), 
      .ZN(n_1_737_4325));
   NOR2_X1 i_1_737_4904 (.A1(n_1_737_254), .A2(n_1_737_5274), .ZN(n_1_737_4326));
   AOI22_X1 i_1_737_4905 (.A1(n_1_737_4421), .A2(n_1_737_4329), .B1(n_1_737_5189), 
      .B2(n_1_737_4328), .ZN(n_1_737_4327));
   OAI21_X1 i_1_737_4906 (.A(n_1_737_4422), .B1(n_1_737_255), .B2(n_1_737_5215), 
      .ZN(n_1_737_4328));
   NOR2_X1 i_1_737_4907 (.A1(n_1_737_255), .A2(n_1_737_5215), .ZN(n_1_737_4329));
   OAI22_X1 i_1_737_4908 (.A1(n_1_737_4445), .A2(n_1_737_4331), .B1(n_1_737_5298), 
      .B2(n_1_737_4332), .ZN(n_1_737_4330));
   NOR2_X1 i_1_737_4909 (.A1(n_1_737_5297), .A2(n_1_737_4333), .ZN(n_1_737_4331));
   INV_X1 i_1_737_4910 (.A(n_1_737_4333), .ZN(n_1_737_4332));
   NOR2_X1 i_1_737_4911 (.A1(n_1_737_253), .A2(n_1_737_5320), .ZN(n_1_737_4333));
   NOR2_X1 i_1_737_4912 (.A1(n_1_737_251), .A2(n_1_737_5155), .ZN(n_578));
   NOR3_X1 i_1_737_4913 (.A1(n_1_737_250), .A2(n_1_737_5167), .A3(n_1_737_4334), 
      .ZN(n_579));
   OAI21_X1 i_1_737_4914 (.A(n_1_737_4334), .B1(n_1_737_250), .B2(n_1_737_5167), 
      .ZN(n_580));
   AOI21_X1 i_1_737_4915 (.A(n_1_737_4401), .B1(n_848), .B2(n_1_737_4883), 
      .ZN(n_1_737_4334));
   OR3_X1 i_1_737_4916 (.A1(n_1_737_4355), .A2(n_1_737_4342), .A3(n_1_737_4335), 
      .ZN(n_581));
   OAI211_X1 i_1_737_4917 (.A(n_1_737_4361), .B(n_1_737_4349), .C1(n_1_737_4337), 
      .C2(n_1_737_4336), .ZN(n_1_737_4335));
   NOR2_X1 i_1_737_4918 (.A1(n_1_737_4339), .A2(n_1_737_4338), .ZN(n_1_737_4336));
   AOI21_X1 i_1_737_4919 (.A(n_1_737_5336), .B1(n_1_737_4339), .B2(n_1_737_4338), 
      .ZN(n_1_737_4337));
   NOR2_X1 i_1_737_4920 (.A1(n_1_737_245), .A2(n_1_737_5358), .ZN(n_1_737_4338));
   NAND3_X1 i_1_737_4921 (.A1(n_1_737_5670), .A2(n_1_737_4340), .A3(n_1_737_5671), 
      .ZN(n_1_737_4339));
   OAI21_X1 i_1_737_4922 (.A(\out_bs[0] [4]), .B1(\out_bs[0] [3]), .B2(
      n_1_737_4905), .ZN(n_1_737_4340));
   NOR2_X1 i_1_737_4923 (.A1(\out_bs[0] [0]), .A2(n_1_737_4435), .ZN(
      n_1_737_4341));
   AOI21_X1 i_1_737_4924 (.A(n_1_737_4343), .B1(n_1_737_5190), .B2(n_1_737_4344), 
      .ZN(n_1_737_4342));
   AOI21_X1 i_1_737_4925 (.A(n_1_737_4348), .B1(n_1_737_5189), .B2(n_1_737_4345), 
      .ZN(n_1_737_4343));
   INV_X1 i_1_737_4926 (.A(n_1_737_4345), .ZN(n_1_737_4344));
   NAND2_X1 i_1_737_4927 (.A1(n_1_737_5638), .A2(n_1_737_4346), .ZN(n_1_737_4345));
   AND2_X1 i_1_737_4928 (.A1(n_1_737_5637), .A2(n_1_737_4347), .ZN(n_1_737_4346));
   OAI21_X1 i_1_737_4929 (.A(\out_bs[3] [4]), .B1(\out_bs[3] [3]), .B2(
      n_1_737_4896), .ZN(n_1_737_4347));
   NOR2_X1 i_1_737_4930 (.A1(n_1_737_248), .A2(n_1_737_5215), .ZN(n_1_737_4348));
   INV_X1 i_1_737_4931 (.A(n_1_737_4350), .ZN(n_1_737_4349));
   OAI21_X1 i_1_737_4932 (.A(n_1_737_4351), .B1(n_1_737_5298), .B2(n_1_737_4352), 
      .ZN(n_1_737_4350));
   OAI21_X1 i_1_737_4933 (.A(n_1_737_4354), .B1(n_1_737_5297), .B2(n_1_737_4353), 
      .ZN(n_1_737_4351));
   INV_X1 i_1_737_4934 (.A(n_1_737_4353), .ZN(n_1_737_4352));
   NOR2_X1 i_1_737_4935 (.A1(n_1_737_246), .A2(n_1_737_5320), .ZN(n_1_737_4353));
   OAI21_X1 i_1_737_4936 (.A(n_1_737_4445), .B1(n_1_737_5662), .B2(n_1_737_4889), 
      .ZN(n_1_737_4354));
   OAI21_X1 i_1_737_4937 (.A(n_1_737_4356), .B1(n_1_737_5236), .B2(n_1_737_4357), 
      .ZN(n_1_737_4355));
   OAI21_X1 i_1_737_4938 (.A(n_1_737_4359), .B1(n_1_737_5235), .B2(n_1_737_4358), 
      .ZN(n_1_737_4356));
   INV_X1 i_1_737_4939 (.A(n_1_737_4358), .ZN(n_1_737_4357));
   NOR2_X1 i_1_737_4940 (.A1(n_1_737_247), .A2(n_1_737_5274), .ZN(n_1_737_4358));
   NAND3_X1 i_1_737_4941 (.A1(n_1_737_5650), .A2(n_1_737_4360), .A3(n_1_737_5651), 
      .ZN(n_1_737_4359));
   OAI21_X1 i_1_737_4942 (.A(\out_bs[2] [4]), .B1(\out_bs[2] [3]), .B2(
      n_1_737_4901), .ZN(n_1_737_4360));
   INV_X1 i_1_737_4943 (.A(n_1_737_4362), .ZN(n_1_737_4361));
   OAI21_X1 i_1_737_4944 (.A(n_1_737_4363), .B1(n_1_737_5366), .B2(n_1_737_4364), 
      .ZN(n_1_737_4362));
   OAI21_X1 i_1_737_4945 (.A(n_1_737_4366), .B1(n_1_737_5365), .B2(n_1_737_4365), 
      .ZN(n_1_737_4363));
   INV_X1 i_1_737_4946 (.A(n_1_737_4365), .ZN(n_1_737_4364));
   NOR2_X1 i_1_737_4947 (.A1(n_1_737_249), .A2(n_1_737_5386), .ZN(n_1_737_4365));
   OAI21_X1 i_1_737_4948 (.A(n_1_737_4458), .B1(n_1_737_5623), .B2(n_1_737_4911), 
      .ZN(n_1_737_4366));
   NOR2_X1 i_1_737_4949 (.A1(n_1_737_244), .A2(n_1_737_5155), .ZN(n_582));
   NOR3_X1 i_1_737_4950 (.A1(n_1_737_243), .A2(n_1_737_5167), .A3(n_1_737_4367), 
      .ZN(n_583));
   OAI21_X1 i_1_737_4951 (.A(n_1_737_4367), .B1(n_1_737_243), .B2(n_1_737_5167), 
      .ZN(n_584));
   AOI21_X1 i_1_737_4952 (.A(n_1_737_4401), .B1(n_848), .B2(n_1_737_4924), 
      .ZN(n_1_737_4367));
   OR4_X1 i_1_737_4953 (.A1(n_1_737_4393), .A2(n_1_737_4370), .A3(n_1_737_4376), 
      .A4(n_1_737_4368), .ZN(n_585));
   OAI211_X1 i_1_737_4954 (.A(n_1_737_4389), .B(n_1_737_4383), .C1(n_1_737_5337), 
      .C2(n_1_737_4390), .ZN(n_1_737_4368));
   INV_X1 i_1_737_4955 (.A(n_1_737_4370), .ZN(n_1_737_4369));
   OAI21_X1 i_1_737_4956 (.A(n_1_737_4371), .B1(n_1_737_5298), .B2(n_1_737_4372), 
      .ZN(n_1_737_4370));
   OAI22_X1 i_1_737_4957 (.A1(\out_bs[1] [6]), .A2(n_1_737_4374), .B1(
      n_1_737_5297), .B2(n_1_737_4373), .ZN(n_1_737_4371));
   INV_X1 i_1_737_4958 (.A(n_1_737_4373), .ZN(n_1_737_4372));
   NOR2_X1 i_1_737_4959 (.A1(n_1_737_239), .A2(n_1_737_5320), .ZN(n_1_737_4373));
   INV_X1 i_1_737_4960 (.A(n_1_737_4375), .ZN(n_1_737_4374));
   AOI21_X1 i_1_737_4961 (.A(n_1_737_4448), .B1(\out_bs[1] [4]), .B2(
      n_1_737_4933), .ZN(n_1_737_4375));
   INV_X1 i_1_737_4962 (.A(n_1_737_4377), .ZN(n_1_737_4376));
   AOI22_X1 i_1_737_4963 (.A1(n_1_737_4382), .A2(n_1_737_4379), .B1(n_1_737_5189), 
      .B2(n_1_737_4378), .ZN(n_1_737_4377));
   OR2_X1 i_1_737_4964 (.A1(n_1_737_4382), .A2(n_1_737_4379), .ZN(n_1_737_4378));
   NAND2_X1 i_1_737_4965 (.A1(n_1_737_5638), .A2(n_1_737_4380), .ZN(n_1_737_4379));
   NOR2_X1 i_1_737_4966 (.A1(n_1_737_4424), .A2(n_1_737_4381), .ZN(n_1_737_4380));
   NOR2_X1 i_1_737_4967 (.A1(n_1_737_5636), .A2(n_1_737_4940), .ZN(n_1_737_4381));
   NOR2_X1 i_1_737_4968 (.A1(n_1_737_241), .A2(n_1_737_5215), .ZN(n_1_737_4382));
   OAI22_X1 i_1_737_4969 (.A1(n_1_737_4388), .A2(n_1_737_4384), .B1(n_1_737_5235), 
      .B2(n_1_737_4385), .ZN(n_1_737_4383));
   AND2_X1 i_1_737_4970 (.A1(n_1_737_5235), .A2(n_1_737_4385), .ZN(n_1_737_4384));
   NAND2_X1 i_1_737_4971 (.A1(n_1_737_5651), .A2(n_1_737_4386), .ZN(n_1_737_4385));
   NOR2_X1 i_1_737_4972 (.A1(n_1_737_4413), .A2(n_1_737_4387), .ZN(n_1_737_4386));
   NOR2_X1 i_1_737_4973 (.A1(n_1_737_5649), .A2(n_1_737_4954), .ZN(n_1_737_4387));
   NOR2_X1 i_1_737_4974 (.A1(n_1_737_240), .A2(n_1_737_5274), .ZN(n_1_737_4388));
   OAI22_X1 i_1_737_4975 (.A1(n_1_737_4434), .A2(n_1_737_4392), .B1(n_1_737_5336), 
      .B2(n_1_737_4391), .ZN(n_1_737_4389));
   INV_X1 i_1_737_4976 (.A(n_1_737_4391), .ZN(n_1_737_4390));
   NOR2_X1 i_1_737_4977 (.A1(n_1_737_238), .A2(n_1_737_5358), .ZN(n_1_737_4391));
   NOR2_X1 i_1_737_4978 (.A1(n_1_737_5669), .A2(n_1_737_4947), .ZN(n_1_737_4392));
   AOI21_X1 i_1_737_4979 (.A(n_1_737_4394), .B1(n_1_737_5366), .B2(n_1_737_4395), 
      .ZN(n_1_737_4393));
   AOI21_X1 i_1_737_4980 (.A(n_1_737_4399), .B1(n_1_737_5365), .B2(n_1_737_4396), 
      .ZN(n_1_737_4394));
   INV_X1 i_1_737_4981 (.A(n_1_737_4396), .ZN(n_1_737_4395));
   NAND2_X1 i_1_737_4982 (.A1(n_1_737_5625), .A2(n_1_737_4397), .ZN(n_1_737_4396));
   NOR2_X1 i_1_737_4983 (.A1(n_1_737_4460), .A2(n_1_737_4398), .ZN(n_1_737_4397));
   NOR2_X1 i_1_737_4984 (.A1(n_1_737_5623), .A2(n_1_737_4961), .ZN(n_1_737_4398));
   NOR2_X1 i_1_737_4985 (.A1(n_1_737_242), .A2(n_1_737_5386), .ZN(n_1_737_4399));
   NOR2_X1 i_1_737_4986 (.A1(n_1_737_237), .A2(n_1_737_5155), .ZN(n_586));
   INV_X1 i_1_737_4992 (.A(n_1_737_4404), .ZN(n_1_737_4403));
   OR4_X1 i_1_737_4994 (.A1(n_1_737_4417), .A2(n_1_737_4405), .A3(n_1_737_4430), 
      .A4(n_1_737_4453), .ZN(n_587));
   OAI21_X1 i_1_737_4995 (.A(n_1_737_4406), .B1(n_1_737_5236), .B2(n_1_737_4407), 
      .ZN(n_1_737_4405));
   OAI22_X1 i_1_737_4996 (.A1(\out_bs[2] [6]), .A2(n_1_737_4412), .B1(
      n_1_737_5235), .B2(n_1_737_4408), .ZN(n_1_737_4406));
   INV_X1 i_1_737_4997 (.A(n_1_737_4408), .ZN(n_1_737_4407));
   NOR2_X1 i_1_737_4998 (.A1(n_1_737_233), .A2(n_1_737_5274), .ZN(n_1_737_4408));
   INV_X1 i_1_737_4999 (.A(n_1_737_4410), .ZN(n_1_737_4409));
   NOR2_X1 i_1_737_5000 (.A1(\out_bs[2] [6]), .A2(n_1_737_4413), .ZN(
      n_1_737_4410));
   INV_X1 i_1_737_5001 (.A(n_1_737_4412), .ZN(n_1_737_4411));
   OAI21_X1 i_1_737_5002 (.A(n_1_737_5650), .B1(n_1_737_5649), .B2(n_1_737_4985), 
      .ZN(n_1_737_4412));
   INV_X1 i_1_737_5003 (.A(n_1_737_4414), .ZN(n_1_737_4413));
   NOR2_X1 i_1_737_5004 (.A1(\out_bs[2] [5]), .A2(n_1_737_4416), .ZN(
      n_1_737_4414));
   INV_X1 i_1_737_5005 (.A(n_1_737_4416), .ZN(n_1_737_4415));
   NOR2_X1 i_1_737_5006 (.A1(n_1_737_5649), .A2(n_1_737_5648), .ZN(n_1_737_4416));
   AOI21_X1 i_1_737_5007 (.A(n_1_737_4418), .B1(n_1_737_5190), .B2(n_1_737_4419), 
      .ZN(n_1_737_4417));
   AOI21_X1 i_1_737_5008 (.A(n_1_737_4429), .B1(n_1_737_5189), .B2(n_1_737_4420), 
      .ZN(n_1_737_4418));
   INV_X1 i_1_737_5009 (.A(n_1_737_4420), .ZN(n_1_737_4419));
   NAND2_X1 i_1_737_5010 (.A1(n_1_737_5638), .A2(n_1_737_4423), .ZN(n_1_737_4420));
   INV_X1 i_1_737_5011 (.A(n_1_737_4422), .ZN(n_1_737_4421));
   NOR2_X1 i_1_737_5012 (.A1(\out_bs[3] [6]), .A2(n_1_737_4424), .ZN(
      n_1_737_4422));
   NOR2_X1 i_1_737_5013 (.A1(n_1_737_4428), .A2(n_1_737_4424), .ZN(n_1_737_4423));
   INV_X1 i_1_737_5014 (.A(n_1_737_4425), .ZN(n_1_737_4424));
   NOR2_X1 i_1_737_5015 (.A1(\out_bs[3] [5]), .A2(n_1_737_4427), .ZN(
      n_1_737_4425));
   INV_X1 i_1_737_5016 (.A(n_1_737_4427), .ZN(n_1_737_4426));
   NOR2_X1 i_1_737_5017 (.A1(n_1_737_5636), .A2(n_1_737_5635), .ZN(n_1_737_4427));
   NOR2_X1 i_1_737_5018 (.A1(n_1_737_5636), .A2(n_1_737_4979), .ZN(n_1_737_4428));
   NOR2_X1 i_1_737_5019 (.A1(n_1_737_234), .A2(n_1_737_5215), .ZN(n_1_737_4429));
   OAI211_X1 i_1_737_5020 (.A(n_1_737_4431), .B(n_1_737_4440), .C1(n_1_737_5337), 
      .C2(n_1_737_4432), .ZN(n_1_737_4430));
   OAI22_X1 i_1_737_5021 (.A1(n_1_737_4439), .A2(n_1_737_4434), .B1(n_1_737_5336), 
      .B2(n_1_737_4433), .ZN(n_1_737_4431));
   INV_X1 i_1_737_5022 (.A(n_1_737_4433), .ZN(n_1_737_4432));
   NOR2_X1 i_1_737_5023 (.A1(n_1_737_231), .A2(n_1_737_5358), .ZN(n_1_737_4433));
   NAND2_X1 i_1_737_5024 (.A1(n_1_737_5671), .A2(n_1_737_4436), .ZN(n_1_737_4434));
   INV_X1 i_1_737_5025 (.A(n_1_737_4436), .ZN(n_1_737_4435));
   NOR2_X1 i_1_737_5026 (.A1(\out_bs[0] [5]), .A2(n_1_737_4438), .ZN(
      n_1_737_4436));
   INV_X1 i_1_737_5027 (.A(n_1_737_4438), .ZN(n_1_737_4437));
   NOR2_X1 i_1_737_5028 (.A1(n_1_737_5669), .A2(n_1_737_5668), .ZN(n_1_737_4438));
   NOR2_X1 i_1_737_5029 (.A1(n_1_737_5669), .A2(n_1_737_4992), .ZN(n_1_737_4439));
   INV_X1 i_1_737_5030 (.A(n_1_737_4441), .ZN(n_1_737_4440));
   OAI21_X1 i_1_737_5031 (.A(n_1_737_4442), .B1(n_1_737_5298), .B2(n_1_737_4443), 
      .ZN(n_1_737_4441));
   OAI22_X1 i_1_737_5032 (.A1(\out_bs[1] [6]), .A2(n_1_737_4446), .B1(
      n_1_737_5297), .B2(n_1_737_4444), .ZN(n_1_737_4442));
   INV_X1 i_1_737_5033 (.A(n_1_737_4444), .ZN(n_1_737_4443));
   NOR2_X1 i_1_737_5034 (.A1(n_1_737_232), .A2(n_1_737_5320), .ZN(n_1_737_4444));
   NOR2_X1 i_1_737_5035 (.A1(\out_bs[1] [6]), .A2(n_1_737_4448), .ZN(
      n_1_737_4445));
   INV_X1 i_1_737_5036 (.A(n_1_737_4447), .ZN(n_1_737_4446));
   NOR2_X1 i_1_737_5037 (.A1(n_1_737_4452), .A2(n_1_737_4448), .ZN(n_1_737_4447));
   INV_X1 i_1_737_5038 (.A(n_1_737_4449), .ZN(n_1_737_4448));
   NOR2_X1 i_1_737_5039 (.A1(\out_bs[1] [5]), .A2(n_1_737_4451), .ZN(
      n_1_737_4449));
   INV_X1 i_1_737_5040 (.A(n_1_737_4451), .ZN(n_1_737_4450));
   NOR2_X1 i_1_737_5041 (.A1(n_1_737_5662), .A2(n_1_737_5661), .ZN(n_1_737_4451));
   NOR2_X1 i_1_737_5042 (.A1(n_1_737_5662), .A2(n_1_737_4971), .ZN(n_1_737_4452));
   OAI22_X1 i_1_737_5044 (.A1(\out_bs[4] [6]), .A2(n_1_737_4459), .B1(
      n_1_737_5365), .B2(n_1_737_4456), .ZN(n_1_737_4454));
   INV_X1 i_1_737_5045 (.A(n_1_737_4456), .ZN(n_1_737_4455));
   NOR2_X1 i_1_737_5046 (.A1(n_1_737_235), .A2(n_1_737_5386), .ZN(n_1_737_4456));
   INV_X1 i_1_737_5047 (.A(n_1_737_4458), .ZN(n_1_737_4457));
   NOR2_X1 i_1_737_5048 (.A1(\out_bs[4] [6]), .A2(n_1_737_4460), .ZN(
      n_1_737_4458));
   OAI21_X1 i_1_737_5049 (.A(n_1_737_5624), .B1(n_1_737_5623), .B2(n_1_737_4999), 
      .ZN(n_1_737_4459));
   INV_X1 i_1_737_5050 (.A(n_1_737_4461), .ZN(n_1_737_4460));
   NOR2_X1 i_1_737_5051 (.A1(\out_bs[4] [5]), .A2(n_1_737_4462), .ZN(
      n_1_737_4461));
   NOR2_X1 i_1_737_5052 (.A1(n_1_737_5623), .A2(n_1_737_5622), .ZN(n_1_737_4462));
   NOR2_X1 i_1_737_5053 (.A1(n_1_737_230), .A2(n_1_737_5155), .ZN(n_588));
   NOR3_X1 i_1_737_5054 (.A1(n_1_737_229), .A2(n_1_737_5167), .A3(n_1_737_4518), 
      .ZN(n_589));
   OAI21_X1 i_1_737_5055 (.A(n_1_737_4518), .B1(n_1_737_229), .B2(n_1_737_5167), 
      .ZN(n_590));
   OAI211_X1 i_1_737_5056 (.A(n_1_737_4463), .B(n_1_737_4478), .C1(n_1_737_4476), 
      .C2(n_1_737_4475), .ZN(n_591));
   AND3_X1 i_1_737_5057 (.A1(n_1_737_4469), .A2(n_1_737_4465), .A3(n_1_737_4472), 
      .ZN(n_1_737_4463));
   INV_X1 i_1_737_5058 (.A(n_1_737_4465), .ZN(n_1_737_4464));
   OAI21_X1 i_1_737_5059 (.A(n_1_737_4466), .B1(n_1_737_5297), .B2(n_1_737_4468), 
      .ZN(n_1_737_4465));
   OAI211_X1 i_1_737_5060 (.A(n_1_737_5285), .B(n_1_737_4528), .C1(n_1_737_5298), 
      .C2(n_1_737_4467), .ZN(n_1_737_4466));
   INV_X1 i_1_737_5061 (.A(n_1_737_4468), .ZN(n_1_737_4467));
   NOR2_X1 i_1_737_5062 (.A1(n_1_737_225), .A2(n_1_737_5320), .ZN(n_1_737_4468));
   AOI22_X1 i_1_737_5063 (.A1(n_1_737_4533), .A2(n_1_737_4471), .B1(n_1_737_5189), 
      .B2(n_1_737_4470), .ZN(n_1_737_4469));
   OAI21_X1 i_1_737_5064 (.A(n_1_737_4534), .B1(n_1_737_227), .B2(n_1_737_5215), 
      .ZN(n_1_737_4470));
   NOR2_X1 i_1_737_5065 (.A1(n_1_737_227), .A2(n_1_737_5215), .ZN(n_1_737_4471));
   OAI22_X1 i_1_737_5066 (.A1(n_1_737_4552), .A2(n_1_737_4473), .B1(n_1_737_5235), 
      .B2(n_1_737_4474), .ZN(n_1_737_4472));
   AND2_X1 i_1_737_5067 (.A1(n_1_737_5235), .A2(n_1_737_4474), .ZN(n_1_737_4473));
   NOR2_X1 i_1_737_5068 (.A1(n_1_737_226), .A2(n_1_737_5274), .ZN(n_1_737_4474));
   NOR2_X1 i_1_737_5069 (.A1(n_1_737_4543), .A2(n_1_737_4477), .ZN(n_1_737_4475));
   AOI21_X1 i_1_737_5070 (.A(n_1_737_5336), .B1(n_1_737_4543), .B2(n_1_737_4477), 
      .ZN(n_1_737_4476));
   NOR2_X1 i_1_737_5071 (.A1(n_1_737_224), .A2(n_1_737_5358), .ZN(n_1_737_4477));
   OAI22_X1 i_1_737_5072 (.A1(n_1_737_4562), .A2(n_1_737_4479), .B1(n_1_737_5365), 
      .B2(n_1_737_4480), .ZN(n_1_737_4478));
   AND2_X1 i_1_737_5073 (.A1(n_1_737_5365), .A2(n_1_737_4480), .ZN(n_1_737_4479));
   NOR2_X1 i_1_737_5074 (.A1(n_1_737_228), .A2(n_1_737_5386), .ZN(n_1_737_4480));
   NOR2_X1 i_1_737_5075 (.A1(n_1_737_223), .A2(n_1_737_5155), .ZN(n_592));
   NOR3_X1 i_1_737_5076 (.A1(n_1_737_222), .A2(n_1_737_5167), .A3(n_1_737_4481), 
      .ZN(n_593));
   OAI21_X1 i_1_737_5077 (.A(n_1_737_4481), .B1(n_1_737_222), .B2(n_1_737_5167), 
      .ZN(n_594));
   AOI21_X1 i_1_737_5078 (.A(n_1_737_5181), .B1(n_848), .B2(n_1_737_5020), 
      .ZN(n_1_737_4481));
   OR4_X1 i_1_737_5079 (.A1(n_1_737_4500), .A2(n_1_737_4494), .A3(n_1_737_4482), 
      .A4(n_1_737_4506), .ZN(n_595));
   OAI211_X1 i_1_737_5080 (.A(n_1_737_4483), .B(n_1_737_4487), .C1(n_1_737_5337), 
      .C2(n_1_737_4484), .ZN(n_1_737_4482));
   OAI22_X1 i_1_737_5081 (.A1(n_1_737_5083), .A2(n_1_737_4486), .B1(n_1_737_5336), 
      .B2(n_1_737_4485), .ZN(n_1_737_4483));
   INV_X1 i_1_737_5082 (.A(n_1_737_4485), .ZN(n_1_737_4484));
   NOR2_X1 i_1_737_5083 (.A1(n_1_737_217), .A2(n_1_737_5358), .ZN(n_1_737_4485));
   NOR2_X1 i_1_737_5084 (.A1(n_1_737_5669), .A2(n_1_737_5028), .ZN(n_1_737_4486));
   OAI22_X1 i_1_737_5085 (.A1(n_1_737_4492), .A2(n_1_737_4488), .B1(n_1_737_5189), 
      .B2(n_1_737_4489), .ZN(n_1_737_4487));
   NOR2_X1 i_1_737_5086 (.A1(n_1_737_5190), .A2(n_1_737_4490), .ZN(n_1_737_4488));
   INV_X1 i_1_737_5087 (.A(n_1_737_4490), .ZN(n_1_737_4489));
   NOR2_X1 i_1_737_5088 (.A1(n_1_737_5221), .A2(n_1_737_4491), .ZN(n_1_737_4490));
   NOR2_X1 i_1_737_5089 (.A1(n_1_737_5636), .A2(n_1_737_5036), .ZN(n_1_737_4491));
   NOR2_X1 i_1_737_5090 (.A1(n_1_737_220), .A2(n_1_737_5215), .ZN(n_1_737_4492));
   INV_X1 i_1_737_5091 (.A(n_1_737_4494), .ZN(n_1_737_4493));
   OAI21_X1 i_1_737_5092 (.A(n_1_737_4495), .B1(n_1_737_5298), .B2(n_1_737_4496), 
      .ZN(n_1_737_4494));
   OAI22_X1 i_1_737_5093 (.A1(n_1_737_5284), .A2(n_1_737_4498), .B1(n_1_737_5297), 
      .B2(n_1_737_4497), .ZN(n_1_737_4495));
   INV_X1 i_1_737_5094 (.A(n_1_737_4497), .ZN(n_1_737_4496));
   NOR2_X1 i_1_737_5095 (.A1(n_1_737_218), .A2(n_1_737_5320), .ZN(n_1_737_4497));
   NOR2_X1 i_1_737_5096 (.A1(n_1_737_5662), .A2(n_1_737_5045), .ZN(n_1_737_4498));
   INV_X1 i_1_737_5097 (.A(n_1_737_4500), .ZN(n_1_737_4499));
   OAI21_X1 i_1_737_5098 (.A(n_1_737_4501), .B1(n_1_737_5236), .B2(n_1_737_4502), 
      .ZN(n_1_737_4500));
   OAI22_X1 i_1_737_5099 (.A1(n_1_737_5252), .A2(n_1_737_4504), .B1(n_1_737_5235), 
      .B2(n_1_737_4503), .ZN(n_1_737_4501));
   INV_X1 i_1_737_5100 (.A(n_1_737_4503), .ZN(n_1_737_4502));
   NOR2_X1 i_1_737_5101 (.A1(n_1_737_219), .A2(n_1_737_5274), .ZN(n_1_737_4503));
   NOR2_X1 i_1_737_5102 (.A1(n_1_737_5649), .A2(n_1_737_5054), .ZN(n_1_737_4504));
   INV_X1 i_1_737_5103 (.A(n_1_737_4506), .ZN(n_1_737_4505));
   OAI21_X1 i_1_737_5104 (.A(n_1_737_4507), .B1(n_1_737_5366), .B2(n_1_737_4508), 
      .ZN(n_1_737_4506));
   OAI22_X1 i_1_737_5105 (.A1(n_1_737_5392), .A2(n_1_737_4510), .B1(n_1_737_5365), 
      .B2(n_1_737_4509), .ZN(n_1_737_4507));
   INV_X1 i_1_737_5106 (.A(n_1_737_4509), .ZN(n_1_737_4508));
   NOR2_X1 i_1_737_5107 (.A1(n_1_737_221), .A2(n_1_737_5386), .ZN(n_1_737_4509));
   NOR2_X1 i_1_737_5108 (.A1(n_1_737_5623), .A2(n_1_737_5063), .ZN(n_1_737_4510));
   NOR3_X1 i_1_737_5109 (.A1(n_1_737_216), .A2(n_1_737_5155), .A3(n_1_737_4511), 
      .ZN(n_596));
   OAI21_X1 i_1_737_5110 (.A(n_1_737_4511), .B1(n_1_737_216), .B2(n_1_737_5155), 
      .ZN(n_597));
   NOR2_X1 i_1_737_5111 (.A1(n_1_737_4914), .A2(n_1_737_4512), .ZN(n_1_737_4511));
   AOI21_X1 i_1_737_5112 (.A(n_1_737_5605), .B1(n_1_737_5604), .B2(n_1_737_4515), 
      .ZN(n_1_737_4512));
   NOR2_X1 i_1_737_5113 (.A1(n_847), .A2(n_851), .ZN(n_1_737_4513));
   INV_X1 i_1_737_5114 (.A(n_1_737_4515), .ZN(n_1_737_4514));
   NOR2_X1 i_1_737_5115 (.A1(n_851), .A2(n_1311), .ZN(n_1_737_4515));
   AOI211_X1 i_1_737_5116 (.A(n_1_737_215), .B(n_1_737_5167), .C1(n_1_737_5182), 
      .C2(n_1_737_4517), .ZN(n_598));
   OAI211_X1 i_1_737_5117 (.A(n_1_737_5182), .B(n_1_737_4517), .C1(n_1_737_215), 
      .C2(n_1_737_5167), .ZN(n_599));
   INV_X1 i_1_737_5118 (.A(n_1_737_4517), .ZN(n_1_737_4516));
   OAI21_X1 i_1_737_5119 (.A(n_848), .B1(n_846), .B2(n_1_737_5073), .ZN(
      n_1_737_4517));
   NOR2_X1 i_1_737_5120 (.A1(n_1_737_5181), .A2(n_1_737_4519), .ZN(n_1_737_4518));
   NOR2_X1 i_1_737_5121 (.A1(n_1_737_5610), .A2(n_1_737_5175), .ZN(n_1_737_4519));
   NAND3_X1 i_1_737_5122 (.A1(n_1_737_4546), .A2(n_1_737_4529), .A3(n_1_737_4520), 
      .ZN(n_600));
   NOR3_X1 i_1_737_5123 (.A1(n_1_737_4556), .A2(n_1_737_4522), .A3(n_1_737_4537), 
      .ZN(n_1_737_4520));
   INV_X1 i_1_737_5124 (.A(n_1_737_4522), .ZN(n_1_737_4521));
   OAI21_X1 i_1_737_5125 (.A(n_1_737_4523), .B1(n_1_737_5298), .B2(n_1_737_4524), 
      .ZN(n_1_737_4522));
   OAI22_X1 i_1_737_5126 (.A1(\out_bs[1] [6]), .A2(n_1_737_4526), .B1(
      n_1_737_5297), .B2(n_1_737_4525), .ZN(n_1_737_4523));
   INV_X1 i_1_737_5127 (.A(n_1_737_4525), .ZN(n_1_737_4524));
   NOR2_X1 i_1_737_5128 (.A1(n_1_737_211), .A2(n_1_737_5320), .ZN(n_1_737_4525));
   NAND2_X1 i_1_737_5129 (.A1(n_1_737_5663), .A2(n_1_737_4527), .ZN(n_1_737_4526));
   OAI21_X1 i_1_737_5130 (.A(\out_bs[1] [4]), .B1(\out_bs[1] [3]), .B2(
      n_1_737_5112), .ZN(n_1_737_4527));
   OAI21_X1 i_1_737_5131 (.A(\out_bs[1] [4]), .B1(\out_bs[1] [3]), .B2(
      \out_bs[1] [2]), .ZN(n_1_737_4528));
   AOI22_X1 i_1_737_5132 (.A1(n_1_737_4536), .A2(n_1_737_4531), .B1(n_1_737_5189), 
      .B2(n_1_737_4530), .ZN(n_1_737_4529));
   OR2_X1 i_1_737_5133 (.A1(n_1_737_4536), .A2(n_1_737_4531), .ZN(n_1_737_4530));
   NAND2_X1 i_1_737_5134 (.A1(n_1_737_5222), .A2(n_1_737_4532), .ZN(n_1_737_4531));
   OAI21_X1 i_1_737_5135 (.A(\out_bs[3] [4]), .B1(\out_bs[3] [3]), .B2(
      n_1_737_5123), .ZN(n_1_737_4532));
   INV_X1 i_1_737_5136 (.A(n_1_737_4534), .ZN(n_1_737_4533));
   NOR2_X1 i_1_737_5137 (.A1(n_1_737_5221), .A2(n_1_737_4535), .ZN(n_1_737_4534));
   NOR2_X1 i_1_737_5138 (.A1(n_1_737_5636), .A2(n_1_737_5225), .ZN(n_1_737_4535));
   NOR2_X1 i_1_737_5139 (.A1(n_1_737_213), .A2(n_1_737_5215), .ZN(n_1_737_4536));
   OAI21_X1 i_1_737_5140 (.A(n_1_737_4538), .B1(n_1_737_5337), .B2(n_1_737_4539), 
      .ZN(n_1_737_4537));
   OAI22_X1 i_1_737_5141 (.A1(n_1_737_4545), .A2(n_1_737_4543), .B1(n_1_737_5336), 
      .B2(n_1_737_4540), .ZN(n_1_737_4538));
   INV_X1 i_1_737_5142 (.A(n_1_737_4540), .ZN(n_1_737_4539));
   NOR2_X1 i_1_737_5143 (.A1(n_1_737_210), .A2(n_1_737_5358), .ZN(n_1_737_4540));
   AND2_X1 i_1_737_5144 (.A1(n_1_737_5670), .A2(n_1_737_4542), .ZN(n_1_737_4541));
   NOR2_X1 i_1_737_5145 (.A1(n_1_737_4545), .A2(n_1_737_4544), .ZN(n_1_737_4542));
   OR2_X1 i_1_737_5146 (.A1(n_1_737_5083), .A2(n_1_737_4544), .ZN(n_1_737_4543));
   NOR2_X1 i_1_737_5147 (.A1(n_1_737_5669), .A2(n_1_737_5329), .ZN(n_1_737_4544));
   NOR2_X1 i_1_737_5148 (.A1(n_1_737_5669), .A2(n_1_737_5666), .ZN(n_1_737_4545));
   AOI21_X1 i_1_737_5149 (.A(n_1_737_4547), .B1(n_1_737_5235), .B2(n_1_737_4549), 
      .ZN(n_1_737_4546));
   INV_X1 i_1_737_5150 (.A(n_1_737_4548), .ZN(n_1_737_4547));
   OAI22_X1 i_1_737_5151 (.A1(\out_bs[2] [6]), .A2(n_1_737_4550), .B1(
      n_1_737_5235), .B2(n_1_737_4549), .ZN(n_1_737_4548));
   NOR2_X1 i_1_737_5152 (.A1(n_1_737_212), .A2(n_1_737_5274), .ZN(n_1_737_4549));
   NAND2_X1 i_1_737_5153 (.A1(n_1_737_5650), .A2(n_1_737_4551), .ZN(n_1_737_4550));
   OAI21_X1 i_1_737_5154 (.A(\out_bs[2] [4]), .B1(\out_bs[2] [3]), .B2(
      n_1_737_5096), .ZN(n_1_737_4551));
   NAND2_X1 i_1_737_5155 (.A1(n_1_737_5651), .A2(n_1_737_4553), .ZN(n_1_737_4552));
   NOR2_X1 i_1_737_5156 (.A1(\out_bs[2] [5]), .A2(n_1_737_4554), .ZN(
      n_1_737_4553));
   NOR2_X1 i_1_737_5157 (.A1(n_1_737_5649), .A2(n_1_737_5257), .ZN(n_1_737_4554));
   INV_X1 i_1_737_5158 (.A(n_1_737_4556), .ZN(n_1_737_4555));
   OAI21_X1 i_1_737_5159 (.A(n_1_737_4557), .B1(n_1_737_5366), .B2(n_1_737_4558), 
      .ZN(n_1_737_4556));
   OAI22_X1 i_1_737_5160 (.A1(n_1_737_5392), .A2(n_1_737_4560), .B1(n_1_737_5365), 
      .B2(n_1_737_4559), .ZN(n_1_737_4557));
   INV_X1 i_1_737_5161 (.A(n_1_737_4559), .ZN(n_1_737_4558));
   NOR2_X1 i_1_737_5162 (.A1(n_1_737_214), .A2(n_1_737_5386), .ZN(n_1_737_4559));
   INV_X1 i_1_737_5163 (.A(n_1_737_4561), .ZN(n_1_737_4560));
   OAI21_X1 i_1_737_5164 (.A(\out_bs[4] [4]), .B1(\out_bs[4] [3]), .B2(
      n_1_737_5131), .ZN(n_1_737_4561));
   NAND2_X1 i_1_737_5165 (.A1(n_1_737_5625), .A2(n_1_737_4563), .ZN(n_1_737_4562));
   NOR2_X1 i_1_737_5166 (.A1(\out_bs[4] [5]), .A2(n_1_737_4564), .ZN(
      n_1_737_4563));
   NOR2_X1 i_1_737_5167 (.A1(n_1_737_5623), .A2(n_1_737_5398), .ZN(n_1_737_4564));
   NOR2_X1 i_1_737_5168 (.A1(n_1_737_209), .A2(n_1_737_5155), .ZN(n_601));
   NOR3_X1 i_1_737_5169 (.A1(n_1_737_208), .A2(n_1_737_5167), .A3(n_1_737_4565), 
      .ZN(n_602));
   OAI21_X1 i_1_737_5170 (.A(n_1_737_4565), .B1(n_1_737_208), .B2(n_1_737_5167), 
      .ZN(n_603));
   AOI21_X1 i_1_737_5171 (.A(n_1_737_5181), .B1(n_848), .B2(n_1_737_5172), 
      .ZN(n_1_737_4565));
   NAND3_X1 i_1_737_5172 (.A1(n_1_737_4584), .A2(n_1_737_4572), .A3(n_1_737_4566), 
      .ZN(n_604));
   NOR3_X1 i_1_737_5173 (.A1(n_1_737_4579), .A2(n_1_737_4567), .A3(n_1_737_4590), 
      .ZN(n_1_737_4566));
   OAI21_X1 i_1_737_5174 (.A(n_1_737_4568), .B1(n_1_737_5337), .B2(n_1_737_4569), 
      .ZN(n_1_737_4567));
   OAI22_X1 i_1_737_5175 (.A1(n_1_737_5083), .A2(n_1_737_4571), .B1(n_1_737_5336), 
      .B2(n_1_737_4570), .ZN(n_1_737_4568));
   INV_X1 i_1_737_5176 (.A(n_1_737_4570), .ZN(n_1_737_4569));
   NOR2_X1 i_1_737_5177 (.A1(n_1_737_203), .A2(n_1_737_5358), .ZN(n_1_737_4570));
   NOR2_X1 i_1_737_5178 (.A1(n_1_737_5669), .A2(n_1_737_5325), .ZN(n_1_737_4571));
   OAI22_X1 i_1_737_5179 (.A1(n_1_737_4577), .A2(n_1_737_4573), .B1(n_1_737_5189), 
      .B2(n_1_737_4574), .ZN(n_1_737_4572));
   NOR2_X1 i_1_737_5180 (.A1(n_1_737_5190), .A2(n_1_737_4575), .ZN(n_1_737_4573));
   INV_X1 i_1_737_5181 (.A(n_1_737_4575), .ZN(n_1_737_4574));
   NOR2_X1 i_1_737_5182 (.A1(n_1_737_5221), .A2(n_1_737_4576), .ZN(n_1_737_4575));
   AND2_X1 i_1_737_5183 (.A1(\out_bs[3] [4]), .A2(n_1_737_5223), .ZN(
      n_1_737_4576));
   NOR2_X1 i_1_737_5184 (.A1(n_1_737_206), .A2(n_1_737_5215), .ZN(n_1_737_4577));
   INV_X1 i_1_737_5185 (.A(n_1_737_4579), .ZN(n_1_737_4578));
   OAI21_X1 i_1_737_5186 (.A(n_1_737_4580), .B1(n_1_737_5298), .B2(n_1_737_4581), 
      .ZN(n_1_737_4579));
   OAI22_X1 i_1_737_5187 (.A1(n_1_737_5284), .A2(n_1_737_4583), .B1(n_1_737_5297), 
      .B2(n_1_737_4582), .ZN(n_1_737_4580));
   INV_X1 i_1_737_5188 (.A(n_1_737_4582), .ZN(n_1_737_4581));
   NOR2_X1 i_1_737_5189 (.A1(n_1_737_204), .A2(n_1_737_5320), .ZN(n_1_737_4582));
   NOR2_X1 i_1_737_5190 (.A1(n_1_737_5662), .A2(n_1_737_5286), .ZN(n_1_737_4583));
   AOI21_X1 i_1_737_5191 (.A(n_1_737_4585), .B1(n_1_737_5235), .B2(n_1_737_4587), 
      .ZN(n_1_737_4584));
   INV_X1 i_1_737_5192 (.A(n_1_737_4586), .ZN(n_1_737_4585));
   OAI22_X1 i_1_737_5193 (.A1(n_1_737_5252), .A2(n_1_737_4588), .B1(n_1_737_5235), 
      .B2(n_1_737_4587), .ZN(n_1_737_4586));
   NOR2_X1 i_1_737_5194 (.A1(n_1_737_205), .A2(n_1_737_5274), .ZN(n_1_737_4587));
   AND2_X1 i_1_737_5195 (.A1(\out_bs[2] [4]), .A2(n_1_737_5254), .ZN(
      n_1_737_4588));
   INV_X1 i_1_737_5196 (.A(n_1_737_4590), .ZN(n_1_737_4589));
   OAI21_X1 i_1_737_5197 (.A(n_1_737_4591), .B1(n_1_737_5366), .B2(n_1_737_4592), 
      .ZN(n_1_737_4590));
   OAI22_X1 i_1_737_5198 (.A1(n_1_737_5392), .A2(n_1_737_4594), .B1(n_1_737_5365), 
      .B2(n_1_737_4593), .ZN(n_1_737_4591));
   INV_X1 i_1_737_5199 (.A(n_1_737_4593), .ZN(n_1_737_4592));
   NOR2_X1 i_1_737_5200 (.A1(n_1_737_207), .A2(n_1_737_5386), .ZN(n_1_737_4593));
   NOR2_X1 i_1_737_5201 (.A1(n_1_737_5623), .A2(n_1_737_5395), .ZN(n_1_737_4594));
   NOR2_X1 i_1_737_5202 (.A1(n_1_737_202), .A2(n_1_737_5155), .ZN(n_605));
   NOR3_X1 i_1_737_5203 (.A1(n_1_737_201), .A2(n_1_737_5167), .A3(n_1_737_5180), 
      .ZN(n_606));
   OAI21_X1 i_1_737_5204 (.A(n_1_737_5180), .B1(n_1_737_201), .B2(n_1_737_5167), 
      .ZN(n_607));
   NAND4_X1 i_1_737_5205 (.A1(n_1_737_4606), .A2(n_1_737_4601), .A3(n_1_737_4598), 
      .A4(n_1_737_4595), .ZN(n_608));
   AOI211_X1 i_1_737_5206 (.A(n_1_737_4596), .B(n_1_737_4609), .C1(n_1_737_5336), 
      .C2(n_1_737_4604), .ZN(n_1_737_4595));
   INV_X1 i_1_737_5207 (.A(n_1_737_4597), .ZN(n_1_737_4596));
   OAI21_X1 i_1_737_5208 (.A(n_1_737_5082), .B1(n_1_737_5336), .B2(n_1_737_4604), 
      .ZN(n_1_737_4597));
   AOI22_X1 i_1_737_5209 (.A1(n_1_737_5219), .A2(n_1_737_4600), .B1(n_1_737_5189), 
      .B2(n_1_737_4599), .ZN(n_1_737_4598));
   OAI21_X1 i_1_737_5210 (.A(n_1_737_5220), .B1(n_1_737_199), .B2(n_1_737_5215), 
      .ZN(n_1_737_4599));
   NOR2_X1 i_1_737_5211 (.A1(n_1_737_199), .A2(n_1_737_5215), .ZN(n_1_737_4600));
   AOI22_X1 i_1_737_5212 (.A1(n_1_737_5390), .A2(n_1_737_4603), .B1(n_1_737_5365), 
      .B2(n_1_737_4602), .ZN(n_1_737_4601));
   OAI21_X1 i_1_737_5213 (.A(n_1_737_5391), .B1(n_1_737_200), .B2(n_1_737_5386), 
      .ZN(n_1_737_4602));
   NOR2_X1 i_1_737_5214 (.A1(n_1_737_200), .A2(n_1_737_5386), .ZN(n_1_737_4603));
   NOR2_X1 i_1_737_5215 (.A1(n_1_737_196), .A2(n_1_737_5358), .ZN(n_1_737_4604));
   INV_X1 i_1_737_5216 (.A(n_1_737_4606), .ZN(n_1_737_4605));
   AOI22_X1 i_1_737_5217 (.A1(n_1_737_5250), .A2(n_1_737_4608), .B1(n_1_737_5235), 
      .B2(n_1_737_4607), .ZN(n_1_737_4606));
   OAI21_X1 i_1_737_5218 (.A(n_1_737_5251), .B1(n_1_737_198), .B2(n_1_737_5274), 
      .ZN(n_1_737_4607));
   NOR2_X1 i_1_737_5219 (.A1(n_1_737_198), .A2(n_1_737_5274), .ZN(n_1_737_4608));
   INV_X1 i_1_737_5220 (.A(n_1_737_4610), .ZN(n_1_737_4609));
   OAI21_X1 i_1_737_5221 (.A(n_1_737_4611), .B1(n_1_737_5297), .B2(n_1_737_4613), 
      .ZN(n_1_737_4610));
   OAI21_X1 i_1_737_5222 (.A(n_1_737_5283), .B1(n_1_737_5298), .B2(n_1_737_4612), 
      .ZN(n_1_737_4611));
   INV_X1 i_1_737_5223 (.A(n_1_737_4613), .ZN(n_1_737_4612));
   NOR2_X1 i_1_737_5224 (.A1(n_1_737_197), .A2(n_1_737_5320), .ZN(n_1_737_4613));
   AOI21_X1 i_1_737_5225 (.A(n_1_737_5166), .B1(n_1_737_5180), .B2(n_1_737_4614), 
      .ZN(n_609));
   NAND3_X1 i_1_737_5226 (.A1(n_1_737_5180), .A2(n_1_737_4614), .A3(n_1_737_5166), 
      .ZN(n_610));
   INV_X1 i_1_737_5227 (.A(n_1_737_4615), .ZN(n_1_737_4614));
   NOR2_X1 i_1_737_5228 (.A1(n_1_737_5609), .A2(n_1_737_4882), .ZN(n_1_737_4615));
   NAND4_X1 i_1_737_5229 (.A1(n_1_737_4618), .A2(n_1_737_4616), .A3(n_1_737_4633), 
      .A4(n_1_737_4639), .ZN(n_611));
   AOI211_X1 i_1_737_5230 (.A(n_1_737_4617), .B(n_1_737_4628), .C1(n_1_737_5356), 
      .C2(n_1_737_5336), .ZN(n_1_737_4616));
   AOI21_X1 i_1_737_5231 (.A(n_1_737_4624), .B1(n_1_737_5357), .B2(n_1_737_5337), 
      .ZN(n_1_737_4617));
   INV_X1 i_1_737_5232 (.A(n_1_737_4619), .ZN(n_1_737_4618));
   OAI21_X1 i_1_737_5233 (.A(n_1_737_4621), .B1(n_1_737_5190), .B2(n_1_737_4620), 
      .ZN(n_1_737_4619));
   NOR3_X1 i_1_737_5234 (.A1(n_1_737_5219), .A2(n_1_737_4623), .A3(n_1_737_5214), 
      .ZN(n_1_737_4620));
   OAI21_X1 i_1_737_5235 (.A(n_1_737_5214), .B1(n_1_737_5219), .B2(n_1_737_4623), 
      .ZN(n_1_737_4621));
   INV_X1 i_1_737_5236 (.A(n_1_737_4623), .ZN(n_1_737_4622));
   NOR2_X1 i_1_737_5237 (.A1(n_1_737_5635), .A2(n_1_737_4895), .ZN(n_1_737_4623));
   NOR2_X1 i_1_737_5238 (.A1(n_1_737_5082), .A2(n_1_737_4625), .ZN(n_1_737_4624));
   INV_X1 i_1_737_5239 (.A(n_1_737_4626), .ZN(n_1_737_4625));
   NAND2_X1 i_1_737_5240 (.A1(\out_bs[0] [3]), .A2(n_1_737_4905), .ZN(
      n_1_737_4626));
   INV_X1 i_1_737_5241 (.A(n_1_737_4628), .ZN(n_1_737_4627));
   OAI22_X1 i_1_737_5242 (.A1(n_1_737_4630), .A2(n_1_737_4629), .B1(n_1_737_5318), 
      .B2(n_1_737_5298), .ZN(n_1_737_4628));
   NOR2_X1 i_1_737_5243 (.A1(n_1_737_5319), .A2(n_1_737_5297), .ZN(n_1_737_4629));
   NOR2_X1 i_1_737_5244 (.A1(n_1_737_5282), .A2(n_1_737_4632), .ZN(n_1_737_4630));
   INV_X1 i_1_737_5245 (.A(n_1_737_4632), .ZN(n_1_737_4631));
   NOR2_X1 i_1_737_5246 (.A1(n_1_737_5661), .A2(n_1_737_4889), .ZN(n_1_737_4632));
   OAI21_X1 i_1_737_5247 (.A(n_1_737_4634), .B1(n_1_737_5235), .B2(n_1_737_4635), 
      .ZN(n_1_737_4633));
   OAI21_X1 i_1_737_5248 (.A(n_1_737_5273), .B1(n_1_737_5236), .B2(n_1_737_4636), 
      .ZN(n_1_737_4634));
   INV_X1 i_1_737_5249 (.A(n_1_737_4636), .ZN(n_1_737_4635));
   NOR2_X1 i_1_737_5250 (.A1(n_1_737_5250), .A2(n_1_737_4637), .ZN(n_1_737_4636));
   INV_X1 i_1_737_5251 (.A(n_1_737_4638), .ZN(n_1_737_4637));
   NAND2_X1 i_1_737_5252 (.A1(\out_bs[2] [3]), .A2(n_1_737_4901), .ZN(
      n_1_737_4638));
   OAI21_X1 i_1_737_5253 (.A(n_1_737_4640), .B1(n_1_737_5365), .B2(n_1_737_4641), 
      .ZN(n_1_737_4639));
   OAI21_X1 i_1_737_5254 (.A(n_1_737_5385), .B1(n_1_737_5366), .B2(n_1_737_4642), 
      .ZN(n_1_737_4640));
   INV_X1 i_1_737_5255 (.A(n_1_737_4642), .ZN(n_1_737_4641));
   NOR2_X1 i_1_737_5256 (.A1(n_1_737_5390), .A2(n_1_737_4644), .ZN(n_1_737_4642));
   INV_X1 i_1_737_5257 (.A(n_1_737_4644), .ZN(n_1_737_4643));
   NOR2_X1 i_1_737_5258 (.A1(n_1_737_5622), .A2(n_1_737_4911), .ZN(n_1_737_4644));
   NOR2_X1 i_1_737_5259 (.A1(n_1_737_195), .A2(n_1_737_5154), .ZN(n_612));
   AOI211_X1 i_1_737_5260 (.A(n_1_737_194), .B(n_1_737_5166), .C1(n_1_737_5180), 
      .C2(n_1_737_4645), .ZN(n_613));
   OAI211_X1 i_1_737_5261 (.A(n_1_737_5180), .B(n_1_737_4645), .C1(n_1_737_194), 
      .C2(n_1_737_5166), .ZN(n_614));
   INV_X1 i_1_737_5262 (.A(n_1_737_4646), .ZN(n_1_737_4645));
   NOR2_X1 i_1_737_5263 (.A1(n_1_737_5609), .A2(n_1_737_4925), .ZN(n_1_737_4646));
   NAND3_X1 i_1_737_5264 (.A1(n_1_737_4660), .A2(n_1_737_4654), .A3(n_1_737_4647), 
      .ZN(n_615));
   AOI211_X1 i_1_737_5265 (.A(n_1_737_4671), .B(n_1_737_4649), .C1(n_1_737_4667), 
      .C2(n_1_737_4666), .ZN(n_1_737_4647));
   INV_X1 i_1_737_5266 (.A(n_1_737_4649), .ZN(n_1_737_4648));
   OAI21_X1 i_1_737_5267 (.A(n_1_737_4651), .B1(n_1_737_5298), .B2(n_1_737_4650), 
      .ZN(n_1_737_4649));
   AOI211_X1 i_1_737_5268 (.A(n_1_737_5282), .B(n_1_737_4652), .C1(n_1_737_5588), 
      .C2(n_1_737_5319), .ZN(n_1_737_4650));
   OAI211_X1 i_1_737_5269 (.A(n_1_737_5588), .B(n_1_737_5319), .C1(n_1_737_5282), 
      .C2(n_1_737_4652), .ZN(n_1_737_4651));
   INV_X1 i_1_737_5270 (.A(n_1_737_4653), .ZN(n_1_737_4652));
   NAND2_X1 i_1_737_5271 (.A1(\out_bs[1] [3]), .A2(n_1_737_4933), .ZN(
      n_1_737_4653));
   INV_X1 i_1_737_5272 (.A(n_1_737_4655), .ZN(n_1_737_4654));
   OAI21_X1 i_1_737_5273 (.A(n_1_737_4657), .B1(n_1_737_5190), .B2(n_1_737_4656), 
      .ZN(n_1_737_4655));
   AOI211_X1 i_1_737_5274 (.A(n_1_737_5219), .B(n_1_737_4659), .C1(n_1_737_5587), 
      .C2(n_1_737_5214), .ZN(n_1_737_4656));
   OAI211_X1 i_1_737_5275 (.A(n_1_737_5587), .B(n_1_737_5214), .C1(n_1_737_5219), 
      .C2(n_1_737_4659), .ZN(n_1_737_4657));
   INV_X1 i_1_737_5276 (.A(n_1_737_4659), .ZN(n_1_737_4658));
   NOR2_X1 i_1_737_5277 (.A1(n_1_737_5635), .A2(n_1_737_4940), .ZN(n_1_737_4659));
   OAI21_X1 i_1_737_5278 (.A(n_1_737_4661), .B1(n_1_737_5235), .B2(n_1_737_4663), 
      .ZN(n_1_737_4660));
   OAI211_X1 i_1_737_5279 (.A(n_1_737_5251), .B(n_1_737_4664), .C1(n_1_737_5236), 
      .C2(n_1_737_4662), .ZN(n_1_737_4661));
   INV_X1 i_1_737_5280 (.A(n_1_737_4663), .ZN(n_1_737_4662));
   NOR2_X1 i_1_737_5281 (.A1(n_1_737_191), .A2(n_1_737_5273), .ZN(n_1_737_4663));
   INV_X1 i_1_737_5282 (.A(n_1_737_4665), .ZN(n_1_737_4664));
   NOR2_X1 i_1_737_5283 (.A1(n_1_737_5648), .A2(n_1_737_4954), .ZN(n_1_737_4665));
   NAND2_X1 i_1_737_5284 (.A1(n_1_737_5337), .A2(n_1_737_4668), .ZN(n_1_737_4666));
   OAI22_X1 i_1_737_5285 (.A1(n_1_737_189), .A2(n_1_737_5357), .B1(n_1_737_5337), 
      .B2(n_1_737_4668), .ZN(n_1_737_4667));
   NOR2_X1 i_1_737_5286 (.A1(n_1_737_5082), .A2(n_1_737_4670), .ZN(n_1_737_4668));
   INV_X1 i_1_737_5287 (.A(n_1_737_4670), .ZN(n_1_737_4669));
   NOR2_X1 i_1_737_5288 (.A1(n_1_737_5668), .A2(n_1_737_4947), .ZN(n_1_737_4670));
   INV_X1 i_1_737_5289 (.A(n_1_737_4672), .ZN(n_1_737_4671));
   OAI21_X1 i_1_737_5290 (.A(n_1_737_4673), .B1(n_1_737_5365), .B2(n_1_737_4675), 
      .ZN(n_1_737_4672));
   OAI211_X1 i_1_737_5291 (.A(n_1_737_5391), .B(n_1_737_4676), .C1(n_1_737_5366), 
      .C2(n_1_737_4674), .ZN(n_1_737_4673));
   INV_X1 i_1_737_5292 (.A(n_1_737_4675), .ZN(n_1_737_4674));
   NOR2_X1 i_1_737_5293 (.A1(n_1_737_193), .A2(n_1_737_5385), .ZN(n_1_737_4675));
   INV_X1 i_1_737_5294 (.A(n_1_737_4677), .ZN(n_1_737_4676));
   NOR2_X1 i_1_737_5295 (.A1(n_1_737_5622), .A2(n_1_737_4961), .ZN(n_1_737_4677));
   NOR2_X1 i_1_737_5296 (.A1(n_1_737_188), .A2(n_1_737_5154), .ZN(n_616));
   AOI211_X1 i_1_737_5297 (.A(n_1_737_187), .B(n_1_737_5166), .C1(n_1_737_5180), 
      .C2(n_1_737_4678), .ZN(n_617));
   OAI211_X1 i_1_737_5298 (.A(n_1_737_5180), .B(n_1_737_4678), .C1(n_1_737_187), 
      .C2(n_1_737_5166), .ZN(n_618));
   INV_X1 i_1_737_5299 (.A(n_1_737_4679), .ZN(n_1_737_4678));
   NOR2_X1 i_1_737_5300 (.A1(n_1_737_5609), .A2(n_1_737_4964), .ZN(n_1_737_4679));
   NAND4_X1 i_1_737_5301 (.A1(n_1_737_4708), .A2(n_1_737_4693), .A3(n_1_737_4687), 
      .A4(n_1_737_4680), .ZN(n_619));
   AOI21_X1 i_1_737_5302 (.A(n_1_737_4701), .B1(n_1_737_4682), .B2(n_1_737_4681), 
      .ZN(n_1_737_4680));
   NAND2_X1 i_1_737_5303 (.A1(n_1_737_5337), .A2(n_1_737_4683), .ZN(n_1_737_4681));
   OAI22_X1 i_1_737_5304 (.A1(n_1_737_182), .A2(n_1_737_5357), .B1(n_1_737_5337), 
      .B2(n_1_737_4683), .ZN(n_1_737_4682));
   NOR2_X1 i_1_737_5305 (.A1(n_1_737_5082), .A2(n_1_737_4686), .ZN(n_1_737_4683));
   NOR2_X1 i_1_737_5306 (.A1(\out_bs[0] [4]), .A2(n_1_737_4686), .ZN(
      n_1_737_4684));
   INV_X1 i_1_737_5307 (.A(n_1_737_4686), .ZN(n_1_737_4685));
   NOR2_X1 i_1_737_5308 (.A1(n_1_737_5668), .A2(n_1_737_4992), .ZN(n_1_737_4686));
   OAI21_X1 i_1_737_5309 (.A(n_1_737_4688), .B1(n_1_737_5189), .B2(n_1_737_4690), 
      .ZN(n_1_737_4687));
   OAI211_X1 i_1_737_5310 (.A(n_1_737_5220), .B(n_1_737_4691), .C1(n_1_737_5190), 
      .C2(n_1_737_4689), .ZN(n_1_737_4688));
   INV_X1 i_1_737_5311 (.A(n_1_737_4690), .ZN(n_1_737_4689));
   NOR2_X1 i_1_737_5312 (.A1(n_1_737_185), .A2(n_1_737_5213), .ZN(n_1_737_4690));
   INV_X1 i_1_737_5313 (.A(n_1_737_4692), .ZN(n_1_737_4691));
   NOR2_X1 i_1_737_5314 (.A1(n_1_737_5635), .A2(n_1_737_4979), .ZN(n_1_737_4692));
   INV_X1 i_1_737_5315 (.A(n_1_737_4694), .ZN(n_1_737_4693));
   OAI21_X1 i_1_737_5316 (.A(n_1_737_4696), .B1(n_1_737_5298), .B2(n_1_737_4695), 
      .ZN(n_1_737_4694));
   AOI211_X1 i_1_737_5317 (.A(n_1_737_5282), .B(n_1_737_4699), .C1(n_1_737_5589), 
      .C2(n_1_737_5319), .ZN(n_1_737_4695));
   OAI211_X1 i_1_737_5318 (.A(n_1_737_5589), .B(n_1_737_5319), .C1(n_1_737_5282), 
      .C2(n_1_737_4699), .ZN(n_1_737_4696));
   NOR2_X1 i_1_737_5319 (.A1(\out_bs[1] [4]), .A2(n_1_737_4699), .ZN(
      n_1_737_4697));
   INV_X1 i_1_737_5320 (.A(n_1_737_4699), .ZN(n_1_737_4698));
   NOR2_X1 i_1_737_5321 (.A1(n_1_737_5661), .A2(n_1_737_4971), .ZN(n_1_737_4699));
   INV_X1 i_1_737_5322 (.A(n_1_737_4701), .ZN(n_1_737_4700));
   OAI21_X1 i_1_737_5323 (.A(n_1_737_4702), .B1(n_1_737_5236), .B2(n_1_737_4703), 
      .ZN(n_1_737_4701));
   OAI22_X1 i_1_737_5324 (.A1(n_1_737_5250), .A2(n_1_737_4707), .B1(n_1_737_5235), 
      .B2(n_1_737_4704), .ZN(n_1_737_4702));
   INV_X1 i_1_737_5325 (.A(n_1_737_4704), .ZN(n_1_737_4703));
   NOR2_X1 i_1_737_5326 (.A1(n_1_737_184), .A2(n_1_737_5273), .ZN(n_1_737_4704));
   NOR2_X1 i_1_737_5327 (.A1(\out_bs[2] [4]), .A2(n_1_737_4707), .ZN(
      n_1_737_4705));
   INV_X1 i_1_737_5328 (.A(n_1_737_4707), .ZN(n_1_737_4706));
   NOR2_X1 i_1_737_5329 (.A1(n_1_737_5648), .A2(n_1_737_4986), .ZN(n_1_737_4707));
   INV_X1 i_1_737_5330 (.A(n_1_737_4709), .ZN(n_1_737_4708));
   OAI21_X1 i_1_737_5331 (.A(n_1_737_4710), .B1(n_1_737_5366), .B2(n_1_737_4711), 
      .ZN(n_1_737_4709));
   OAI22_X1 i_1_737_5332 (.A1(n_1_737_5390), .A2(n_1_737_4715), .B1(n_1_737_5365), 
      .B2(n_1_737_4712), .ZN(n_1_737_4710));
   INV_X1 i_1_737_5333 (.A(n_1_737_4712), .ZN(n_1_737_4711));
   NOR2_X1 i_1_737_5334 (.A1(n_1_737_186), .A2(n_1_737_5385), .ZN(n_1_737_4712));
   NOR2_X1 i_1_737_5335 (.A1(\out_bs[4] [4]), .A2(n_1_737_4715), .ZN(
      n_1_737_4713));
   INV_X1 i_1_737_5336 (.A(n_1_737_4715), .ZN(n_1_737_4714));
   NOR2_X1 i_1_737_5337 (.A1(n_1_737_5622), .A2(n_1_737_5000), .ZN(n_1_737_4715));
   NOR2_X1 i_1_737_5338 (.A1(n_1_737_181), .A2(n_1_737_5154), .ZN(n_620));
   NOR3_X1 i_1_737_5339 (.A1(n_1_737_180), .A2(n_1_737_5166), .A3(n_1_737_4739), 
      .ZN(n_621));
   OAI21_X1 i_1_737_5340 (.A(n_1_737_4739), .B1(n_1_737_180), .B2(n_1_737_5166), 
      .ZN(n_622));
   NAND3_X1 i_1_737_5341 (.A1(n_1_737_4720), .A2(n_1_737_4716), .A3(n_1_737_4723), 
      .ZN(n_623));
   OAI21_X1 i_1_737_5342 (.A(n_1_737_4717), .B1(n_1_737_5336), .B2(n_1_737_4719), 
      .ZN(n_1_737_4716));
   OAI22_X1 i_1_737_5343 (.A1(n_1_737_175), .A2(n_1_737_5357), .B1(n_1_737_5337), 
      .B2(n_1_737_4718), .ZN(n_1_737_4717));
   INV_X1 i_1_737_5344 (.A(n_1_737_4719), .ZN(n_1_737_4718));
   NAND2_X1 i_1_737_5345 (.A1(n_1_737_5671), .A2(n_1_737_4776), .ZN(n_1_737_4719));
   AOI21_X1 i_1_737_5346 (.A(n_1_737_4722), .B1(n_1_737_5365), .B2(n_1_737_4721), 
      .ZN(n_1_737_4720));
   OAI211_X1 i_1_737_5347 (.A(n_1_737_5625), .B(n_1_737_4786), .C1(n_1_737_179), 
      .C2(n_1_737_5385), .ZN(n_1_737_4721));
   AOI211_X1 i_1_737_5348 (.A(n_1_737_179), .B(n_1_737_5385), .C1(n_1_737_5625), 
      .C2(n_1_737_4786), .ZN(n_1_737_4722));
   NOR3_X1 i_1_737_5349 (.A1(n_1_737_4728), .A2(n_1_737_4724), .A3(n_1_737_4732), 
      .ZN(n_1_737_4723));
   INV_X1 i_1_737_5350 (.A(n_1_737_4725), .ZN(n_1_737_4724));
   AOI21_X1 i_1_737_5351 (.A(n_1_737_4727), .B1(n_1_737_5297), .B2(n_1_737_4726), 
      .ZN(n_1_737_4725));
   OAI211_X1 i_1_737_5352 (.A(n_1_737_5664), .B(n_1_737_4749), .C1(n_1_737_176), 
      .C2(n_1_737_5318), .ZN(n_1_737_4726));
   AOI211_X1 i_1_737_5353 (.A(n_1_737_176), .B(n_1_737_5318), .C1(n_1_737_5664), 
      .C2(n_1_737_4749), .ZN(n_1_737_4727));
   INV_X1 i_1_737_5354 (.A(n_1_737_4729), .ZN(n_1_737_4728));
   AOI21_X1 i_1_737_5355 (.A(n_1_737_4731), .B1(n_1_737_5189), .B2(n_1_737_4730), 
      .ZN(n_1_737_4729));
   OAI211_X1 i_1_737_5356 (.A(n_1_737_5638), .B(n_1_737_4759), .C1(n_1_737_178), 
      .C2(n_1_737_5213), .ZN(n_1_737_4730));
   AOI211_X1 i_1_737_5357 (.A(n_1_737_178), .B(n_1_737_5213), .C1(n_1_737_5638), 
      .C2(n_1_737_4759), .ZN(n_1_737_4731));
   AOI21_X1 i_1_737_5358 (.A(n_1_737_4733), .B1(n_1_737_5236), .B2(n_1_737_4734), 
      .ZN(n_1_737_4732));
   AOI211_X1 i_1_737_5359 (.A(n_1_737_5250), .B(n_1_737_4772), .C1(n_1_737_5235), 
      .C2(n_1_737_4735), .ZN(n_1_737_4733));
   INV_X1 i_1_737_5360 (.A(n_1_737_4735), .ZN(n_1_737_4734));
   NOR2_X1 i_1_737_5361 (.A1(n_1_737_177), .A2(n_1_737_5273), .ZN(n_1_737_4735));
   NOR2_X1 i_1_737_5362 (.A1(n_1_737_174), .A2(n_1_737_5154), .ZN(n_624));
   NOR3_X1 i_1_737_5363 (.A1(n_1_737_173), .A2(n_1_737_5166), .A3(n_1_737_4736), 
      .ZN(n_625));
   OAI21_X1 i_1_737_5364 (.A(n_1_737_4736), .B1(n_1_737_173), .B2(n_1_737_5166), 
      .ZN(n_626));
   NOR2_X1 i_1_737_5365 (.A1(n_1_737_5181), .A2(n_1_737_4738), .ZN(n_1_737_4736));
   INV_X1 i_1_737_5366 (.A(n_1_737_4738), .ZN(n_1_737_4737));
   OAI21_X1 i_1_737_5367 (.A(n_1_737_4740), .B1(n_1_737_5609), .B2(n_1_737_5023), 
      .ZN(n_1_737_4738));
   NOR2_X1 i_1_737_5368 (.A1(n_1_737_5181), .A2(n_1_737_4741), .ZN(n_1_737_4739));
   INV_X1 i_1_737_5369 (.A(n_1_737_4741), .ZN(n_1_737_4740));
   OAI21_X1 i_1_737_5370 (.A(n_1_737_5610), .B1(n_1_737_5609), .B2(n_1_737_5608), 
      .ZN(n_1_737_4741));
   NAND3_X1 i_1_737_5371 (.A1(n_1_737_4764), .A2(n_1_737_4754), .A3(n_1_737_4742), 
      .ZN(n_627));
   AOI211_X1 i_1_737_5372 (.A(n_1_737_4781), .B(n_1_737_4743), .C1(n_1_737_4774), 
      .C2(n_1_737_4773), .ZN(n_1_737_4742));
   INV_X1 i_1_737_5373 (.A(n_1_737_4744), .ZN(n_1_737_4743));
   AOI22_X1 i_1_737_5374 (.A1(n_1_737_4747), .A2(n_1_737_4746), .B1(n_1_737_5297), 
      .B2(n_1_737_4745), .ZN(n_1_737_4744));
   OAI21_X1 i_1_737_5375 (.A(n_1_737_4748), .B1(n_1_737_169), .B2(n_1_737_5318), 
      .ZN(n_1_737_4745));
   NOR2_X1 i_1_737_5376 (.A1(n_1_737_169), .A2(n_1_737_5318), .ZN(n_1_737_4746));
   INV_X1 i_1_737_5377 (.A(n_1_737_4748), .ZN(n_1_737_4747));
   NOR2_X1 i_1_737_5378 (.A1(n_1_737_5284), .A2(n_1_737_4751), .ZN(n_1_737_4748));
   NOR2_X1 i_1_737_5379 (.A1(n_1_737_5292), .A2(n_1_737_4753), .ZN(n_1_737_4749));
   INV_X1 i_1_737_5380 (.A(n_1_737_4751), .ZN(n_1_737_4750));
   OAI21_X1 i_1_737_5381 (.A(n_1_737_4752), .B1(n_1_737_5661), .B2(n_1_737_5048), 
      .ZN(n_1_737_4751));
   NOR2_X1 i_1_737_5382 (.A1(\out_bs[1] [4]), .A2(n_1_737_4753), .ZN(
      n_1_737_4752));
   NOR2_X1 i_1_737_5383 (.A1(n_1_737_5661), .A2(n_1_737_5660), .ZN(n_1_737_4753));
   AOI22_X1 i_1_737_5384 (.A1(n_1_737_4757), .A2(n_1_737_4756), .B1(n_1_737_5189), 
      .B2(n_1_737_4755), .ZN(n_1_737_4754));
   OAI21_X1 i_1_737_5385 (.A(n_1_737_4758), .B1(n_1_737_171), .B2(n_1_737_5213), 
      .ZN(n_1_737_4755));
   NOR2_X1 i_1_737_5386 (.A1(n_1_737_171), .A2(n_1_737_5213), .ZN(n_1_737_4756));
   INV_X1 i_1_737_5387 (.A(n_1_737_4758), .ZN(n_1_737_4757));
   NOR2_X1 i_1_737_5388 (.A1(n_1_737_5221), .A2(n_1_737_4761), .ZN(n_1_737_4758));
   NOR2_X1 i_1_737_5389 (.A1(n_1_737_5228), .A2(n_1_737_4763), .ZN(n_1_737_4759));
   INV_X1 i_1_737_5390 (.A(n_1_737_4761), .ZN(n_1_737_4760));
   OAI21_X1 i_1_737_5391 (.A(n_1_737_4762), .B1(n_1_737_5635), .B2(n_1_737_5039), 
      .ZN(n_1_737_4761));
   NOR2_X1 i_1_737_5392 (.A1(\out_bs[3] [4]), .A2(n_1_737_4763), .ZN(
      n_1_737_4762));
   NOR2_X1 i_1_737_5393 (.A1(n_1_737_5635), .A2(n_1_737_5634), .ZN(n_1_737_4763));
   OAI21_X1 i_1_737_5394 (.A(n_1_737_4765), .B1(n_1_737_5235), .B2(n_1_737_4767), 
      .ZN(n_1_737_4764));
   OAI211_X1 i_1_737_5395 (.A(n_1_737_5253), .B(n_1_737_4769), .C1(n_1_737_5236), 
      .C2(n_1_737_4766), .ZN(n_1_737_4765));
   INV_X1 i_1_737_5396 (.A(n_1_737_4767), .ZN(n_1_737_4766));
   NOR2_X1 i_1_737_5397 (.A1(n_1_737_170), .A2(n_1_737_5273), .ZN(n_1_737_4767));
   NOR2_X1 i_1_737_5398 (.A1(n_1_737_5259), .A2(n_1_737_4772), .ZN(n_1_737_4768));
   INV_X1 i_1_737_5399 (.A(n_1_737_4770), .ZN(n_1_737_4769));
   OAI21_X1 i_1_737_5400 (.A(n_1_737_4771), .B1(n_1_737_5648), .B2(n_1_737_5056), 
      .ZN(n_1_737_4770));
   NOR2_X1 i_1_737_5401 (.A1(\out_bs[2] [4]), .A2(n_1_737_4772), .ZN(
      n_1_737_4771));
   NOR2_X1 i_1_737_5402 (.A1(n_1_737_5648), .A2(n_1_737_5647), .ZN(n_1_737_4772));
   NAND2_X1 i_1_737_5403 (.A1(n_1_737_5337), .A2(n_1_737_4775), .ZN(n_1_737_4773));
   OAI22_X1 i_1_737_5404 (.A1(n_1_737_168), .A2(n_1_737_5357), .B1(n_1_737_5337), 
      .B2(n_1_737_4775), .ZN(n_1_737_4774));
   NOR2_X1 i_1_737_5405 (.A1(n_1_737_5083), .A2(n_1_737_4778), .ZN(n_1_737_4775));
   NOR2_X1 i_1_737_5406 (.A1(n_1_737_5331), .A2(n_1_737_4780), .ZN(n_1_737_4776));
   INV_X1 i_1_737_5407 (.A(n_1_737_4778), .ZN(n_1_737_4777));
   OAI21_X1 i_1_737_5408 (.A(n_1_737_4779), .B1(n_1_737_5668), .B2(n_1_737_5029), 
      .ZN(n_1_737_4778));
   NOR2_X1 i_1_737_5409 (.A1(\out_bs[0] [4]), .A2(n_1_737_4780), .ZN(
      n_1_737_4779));
   NOR2_X1 i_1_737_5410 (.A1(n_1_737_5668), .A2(n_1_737_5667), .ZN(n_1_737_4780));
   INV_X1 i_1_737_5411 (.A(n_1_737_4782), .ZN(n_1_737_4781));
   OAI22_X1 i_1_737_5412 (.A1(n_1_737_4785), .A2(n_1_737_4783), .B1(n_1_737_5365), 
      .B2(n_1_737_4784), .ZN(n_1_737_4782));
   AND2_X1 i_1_737_5413 (.A1(n_1_737_5365), .A2(n_1_737_4784), .ZN(n_1_737_4783));
   NOR2_X1 i_1_737_5414 (.A1(n_1_737_172), .A2(n_1_737_5385), .ZN(n_1_737_4784));
   NAND2_X1 i_1_737_5415 (.A1(n_1_737_5393), .A2(n_1_737_4787), .ZN(n_1_737_4785));
   NOR2_X1 i_1_737_5416 (.A1(n_1_737_5400), .A2(n_1_737_4790), .ZN(n_1_737_4786));
   INV_X1 i_1_737_5417 (.A(n_1_737_4788), .ZN(n_1_737_4787));
   OAI21_X1 i_1_737_5418 (.A(n_1_737_4789), .B1(n_1_737_5622), .B2(n_1_737_5066), 
      .ZN(n_1_737_4788));
   NOR2_X1 i_1_737_5419 (.A1(\out_bs[4] [4]), .A2(n_1_737_4790), .ZN(
      n_1_737_4789));
   NOR2_X1 i_1_737_5420 (.A1(n_1_737_5622), .A2(n_1_737_5621), .ZN(n_1_737_4790));
   NOR2_X1 i_1_737_5421 (.A1(n_1_737_167), .A2(n_1_737_5154), .ZN(n_628));
   NOR3_X1 i_1_737_5422 (.A1(n_1_737_166), .A2(n_1_737_5166), .A3(n_1_737_4811), 
      .ZN(n_629));
   OAI21_X1 i_1_737_5423 (.A(n_1_737_4811), .B1(n_1_737_166), .B2(n_1_737_5166), 
      .ZN(n_630));
   NAND4_X1 i_1_737_5424 (.A1(n_1_737_4795), .A2(n_1_737_4791), .A3(n_1_737_4801), 
      .A4(n_1_737_4805), .ZN(n_631));
   AOI211_X1 i_1_737_5425 (.A(n_1_737_4798), .B(n_1_737_4792), .C1(n_1_737_4821), 
      .C2(n_1_737_4800), .ZN(n_1_737_4791));
   INV_X1 i_1_737_5426 (.A(n_1_737_4793), .ZN(n_1_737_4792));
   OAI21_X1 i_1_737_5427 (.A(n_1_737_4794), .B1(n_1_737_5297), .B2(n_1_737_4842), 
      .ZN(n_1_737_4793));
   OAI22_X1 i_1_737_5428 (.A1(n_1_737_162), .A2(n_1_737_5318), .B1(n_1_737_5298), 
      .B2(n_1_737_4843), .ZN(n_1_737_4794));
   AOI22_X1 i_1_737_5429 (.A1(n_1_737_4832), .A2(n_1_737_4797), .B1(n_1_737_5189), 
      .B2(n_1_737_4796), .ZN(n_1_737_4795));
   OAI21_X1 i_1_737_5430 (.A(n_1_737_4833), .B1(n_1_737_164), .B2(n_1_737_5213), 
      .ZN(n_1_737_4796));
   NOR2_X1 i_1_737_5431 (.A1(n_1_737_164), .A2(n_1_737_5213), .ZN(n_1_737_4797));
   INV_X1 i_1_737_5432 (.A(n_1_737_4799), .ZN(n_1_737_4798));
   OAI21_X1 i_1_737_5433 (.A(n_1_737_5336), .B1(n_1_737_4821), .B2(n_1_737_4800), 
      .ZN(n_1_737_4799));
   NOR2_X1 i_1_737_5434 (.A1(n_1_737_161), .A2(n_1_737_5357), .ZN(n_1_737_4800));
   OAI21_X1 i_1_737_5435 (.A(n_1_737_4802), .B1(n_1_737_5235), .B2(n_1_737_4804), 
      .ZN(n_1_737_4801));
   OAI211_X1 i_1_737_5436 (.A(n_1_737_5251), .B(n_1_737_4853), .C1(n_1_737_5236), 
      .C2(n_1_737_4803), .ZN(n_1_737_4802));
   INV_X1 i_1_737_5437 (.A(n_1_737_4804), .ZN(n_1_737_4803));
   NOR2_X1 i_1_737_5438 (.A1(n_1_737_163), .A2(n_1_737_5273), .ZN(n_1_737_4804));
   OAI21_X1 i_1_737_5439 (.A(n_1_737_4806), .B1(n_1_737_5365), .B2(n_1_737_4808), 
      .ZN(n_1_737_4805));
   OAI211_X1 i_1_737_5440 (.A(n_1_737_5391), .B(n_1_737_4862), .C1(n_1_737_5366), 
      .C2(n_1_737_4807), .ZN(n_1_737_4806));
   INV_X1 i_1_737_5441 (.A(n_1_737_4808), .ZN(n_1_737_4807));
   NOR2_X1 i_1_737_5442 (.A1(n_1_737_165), .A2(n_1_737_5385), .ZN(n_1_737_4808));
   NOR2_X1 i_1_737_5443 (.A1(n_1_737_160), .A2(n_1_737_5154), .ZN(n_632));
   AOI211_X1 i_1_737_5444 (.A(n_1_737_159), .B(n_1_737_5166), .C1(n_1_737_5180), 
      .C2(n_1_737_4809), .ZN(n_633));
   OAI211_X1 i_1_737_5445 (.A(n_1_737_5180), .B(n_1_737_4809), .C1(n_1_737_159), 
      .C2(n_1_737_5166), .ZN(n_634));
   INV_X1 i_1_737_5446 (.A(n_1_737_4810), .ZN(n_1_737_4809));
   AOI21_X1 i_1_737_5447 (.A(n_1_737_5609), .B1(n_1_737_5608), .B2(n_1_737_5183), 
      .ZN(n_1_737_4810));
   NOR2_X1 i_1_737_5448 (.A1(n_1_737_5179), .A2(n_1_737_4814), .ZN(n_1_737_4811));
   NAND2_X1 i_1_737_5449 (.A1(n_1_737_5610), .A2(n_1_737_4813), .ZN(n_1_737_4812));
   INV_X1 i_1_737_5450 (.A(n_1_737_4814), .ZN(n_1_737_4813));
   NOR2_X1 i_1_737_5451 (.A1(n_1_737_5609), .A2(n_1_737_5074), .ZN(n_1_737_4814));
   NAND4_X1 i_1_737_5452 (.A1(n_1_737_4855), .A2(n_1_737_4836), .A3(n_1_737_4825), 
      .A4(n_1_737_4815), .ZN(n_635));
   AOI21_X1 i_1_737_5453 (.A(n_1_737_4846), .B1(n_1_737_4817), .B2(n_1_737_4816), 
      .ZN(n_1_737_4815));
   NAND2_X1 i_1_737_5454 (.A1(n_1_737_5337), .A2(n_1_737_4818), .ZN(n_1_737_4816));
   OAI22_X1 i_1_737_5455 (.A1(n_1_737_154), .A2(n_1_737_5357), .B1(n_1_737_5337), 
      .B2(n_1_737_4818), .ZN(n_1_737_4817));
   NOR2_X1 i_1_737_5456 (.A1(n_1_737_5082), .A2(n_1_737_4819), .ZN(n_1_737_4818));
   INV_X1 i_1_737_5457 (.A(n_1_737_4820), .ZN(n_1_737_4819));
   NOR2_X1 i_1_737_5458 (.A1(n_1_737_4824), .A2(n_1_737_4823), .ZN(n_1_737_4820));
   NAND3_X1 i_1_737_5459 (.A1(n_1_737_5671), .A2(n_1_737_5332), .A3(n_1_737_4822), 
      .ZN(n_1_737_4821));
   INV_X1 i_1_737_5460 (.A(n_1_737_4823), .ZN(n_1_737_4822));
   NOR2_X1 i_1_737_5461 (.A1(n_1_737_5668), .A2(n_1_737_5085), .ZN(n_1_737_4823));
   NOR2_X1 i_1_737_5462 (.A1(n_1_737_5668), .A2(n_1_737_5665), .ZN(n_1_737_4824));
   OAI21_X1 i_1_737_5463 (.A(n_1_737_4826), .B1(n_1_737_5189), .B2(n_1_737_4828), 
      .ZN(n_1_737_4825));
   OAI211_X1 i_1_737_5464 (.A(n_1_737_5220), .B(n_1_737_4830), .C1(n_1_737_5190), 
      .C2(n_1_737_4827), .ZN(n_1_737_4826));
   INV_X1 i_1_737_5465 (.A(n_1_737_4828), .ZN(n_1_737_4827));
   NOR2_X1 i_1_737_5466 (.A1(n_1_737_157), .A2(n_1_737_5213), .ZN(n_1_737_4828));
   NOR2_X1 i_1_737_5467 (.A1(\out_bs[3] [4]), .A2(n_1_737_4831), .ZN(
      n_1_737_4829));
   INV_X1 i_1_737_5468 (.A(n_1_737_4831), .ZN(n_1_737_4830));
   AOI21_X1 i_1_737_5469 (.A(n_1_737_5635), .B1(n_1_737_5634), .B2(n_1_737_5232), 
      .ZN(n_1_737_4831));
   INV_X1 i_1_737_5470 (.A(n_1_737_4833), .ZN(n_1_737_4832));
   NOR2_X1 i_1_737_5471 (.A1(n_1_737_5219), .A2(n_1_737_4835), .ZN(n_1_737_4833));
   INV_X1 i_1_737_5472 (.A(n_1_737_4835), .ZN(n_1_737_4834));
   NOR2_X1 i_1_737_5473 (.A1(n_1_737_5635), .A2(n_1_737_5124), .ZN(n_1_737_4835));
   INV_X1 i_1_737_5474 (.A(n_1_737_4837), .ZN(n_1_737_4836));
   OAI21_X1 i_1_737_5475 (.A(n_1_737_4839), .B1(n_1_737_5298), .B2(n_1_737_4838), 
      .ZN(n_1_737_4837));
   AOI211_X1 i_1_737_5476 (.A(n_1_737_5282), .B(n_1_737_4841), .C1(n_1_737_5590), 
      .C2(n_1_737_5319), .ZN(n_1_737_4838));
   OAI211_X1 i_1_737_5477 (.A(n_1_737_5590), .B(n_1_737_5319), .C1(n_1_737_5282), 
      .C2(n_1_737_4841), .ZN(n_1_737_4839));
   INV_X1 i_1_737_5478 (.A(n_1_737_4841), .ZN(n_1_737_4840));
   AOI21_X1 i_1_737_5479 (.A(n_1_737_5661), .B1(n_1_737_5660), .B2(n_1_737_5296), 
      .ZN(n_1_737_4841));
   INV_X1 i_1_737_5480 (.A(n_1_737_4843), .ZN(n_1_737_4842));
   NOR2_X1 i_1_737_5481 (.A1(n_1_737_5282), .A2(n_1_737_4845), .ZN(n_1_737_4843));
   INV_X1 i_1_737_5482 (.A(n_1_737_4845), .ZN(n_1_737_4844));
   NOR2_X1 i_1_737_5483 (.A1(n_1_737_5661), .A2(n_1_737_5113), .ZN(n_1_737_4845));
   OAI21_X1 i_1_737_5484 (.A(n_1_737_4847), .B1(n_1_737_5236), .B2(n_1_737_4848), 
      .ZN(n_1_737_4846));
   OAI22_X1 i_1_737_5485 (.A1(n_1_737_5250), .A2(n_1_737_4852), .B1(n_1_737_5235), 
      .B2(n_1_737_4849), .ZN(n_1_737_4847));
   INV_X1 i_1_737_5486 (.A(n_1_737_4849), .ZN(n_1_737_4848));
   NOR2_X1 i_1_737_5487 (.A1(n_1_737_156), .A2(n_1_737_5273), .ZN(n_1_737_4849));
   NOR2_X1 i_1_737_5488 (.A1(\out_bs[2] [4]), .A2(n_1_737_4852), .ZN(
      n_1_737_4850));
   INV_X1 i_1_737_5489 (.A(n_1_737_4852), .ZN(n_1_737_4851));
   AOI21_X1 i_1_737_5490 (.A(n_1_737_5648), .B1(n_1_737_5647), .B2(n_1_737_5263), 
      .ZN(n_1_737_4852));
   INV_X1 i_1_737_5491 (.A(n_1_737_4854), .ZN(n_1_737_4853));
   NOR2_X1 i_1_737_5492 (.A1(n_1_737_5648), .A2(n_1_737_5097), .ZN(n_1_737_4854));
   INV_X1 i_1_737_5493 (.A(n_1_737_4856), .ZN(n_1_737_4855));
   OAI21_X1 i_1_737_5494 (.A(n_1_737_4857), .B1(n_1_737_5366), .B2(n_1_737_4858), 
      .ZN(n_1_737_4856));
   OAI22_X1 i_1_737_5495 (.A1(n_1_737_5390), .A2(n_1_737_4860), .B1(n_1_737_5365), 
      .B2(n_1_737_4859), .ZN(n_1_737_4857));
   INV_X1 i_1_737_5496 (.A(n_1_737_4859), .ZN(n_1_737_4858));
   NOR2_X1 i_1_737_5497 (.A1(n_1_737_158), .A2(n_1_737_5385), .ZN(n_1_737_4859));
   INV_X1 i_1_737_5498 (.A(n_1_737_4861), .ZN(n_1_737_4860));
   OAI21_X1 i_1_737_5499 (.A(\out_bs[4] [3]), .B1(\out_bs[4] [2]), .B2(
      n_1_737_5404), .ZN(n_1_737_4861));
   INV_X1 i_1_737_5500 (.A(n_1_737_4863), .ZN(n_1_737_4862));
   NOR2_X1 i_1_737_5501 (.A1(n_1_737_5622), .A2(n_1_737_5132), .ZN(n_1_737_4863));
   NOR2_X1 i_1_737_5502 (.A1(n_1_737_153), .A2(n_1_737_5154), .ZN(n_636));
   NOR3_X1 i_1_737_5503 (.A1(n_1_737_152), .A2(n_1_737_5166), .A3(n_1_737_5176), 
      .ZN(n_637));
   OAI21_X1 i_1_737_5504 (.A(n_1_737_5176), .B1(n_1_737_152), .B2(n_1_737_5166), 
      .ZN(n_638));
   NAND3_X1 i_1_737_5505 (.A1(n_1_737_4877), .A2(n_1_737_4867), .A3(n_1_737_4864), 
      .ZN(n_639));
   AND3_X1 i_1_737_5506 (.A1(n_1_737_4874), .A2(n_1_737_4870), .A3(n_1_737_4865), 
      .ZN(n_1_737_4864));
   OAI22_X1 i_1_737_5507 (.A1(n_1_737_4880), .A2(n_1_737_4866), .B1(n_1_737_5336), 
      .B2(n_1_737_5080), .ZN(n_1_737_4865));
   NOR2_X1 i_1_737_5508 (.A1(n_1_737_5337), .A2(n_1_737_5081), .ZN(n_1_737_4866));
   AOI22_X1 i_1_737_5509 (.A1(n_1_737_5121), .A2(n_1_737_4869), .B1(n_1_737_5189), 
      .B2(n_1_737_4868), .ZN(n_1_737_4867));
   OAI21_X1 i_1_737_5510 (.A(n_1_737_5122), .B1(n_1_737_150), .B2(n_1_737_5213), 
      .ZN(n_1_737_4868));
   NOR2_X1 i_1_737_5511 (.A1(n_1_737_150), .A2(n_1_737_5213), .ZN(n_1_737_4869));
   AOI22_X1 i_1_737_5512 (.A1(n_1_737_5129), .A2(n_1_737_4872), .B1(n_1_737_5365), 
      .B2(n_1_737_4871), .ZN(n_1_737_4870));
   OAI21_X1 i_1_737_5513 (.A(n_1_737_5130), .B1(n_1_737_151), .B2(n_1_737_5385), 
      .ZN(n_1_737_4871));
   NOR2_X1 i_1_737_5514 (.A1(n_1_737_151), .A2(n_1_737_5385), .ZN(n_1_737_4872));
   INV_X1 i_1_737_5515 (.A(n_1_737_4874), .ZN(n_1_737_4873));
   OAI22_X1 i_1_737_5516 (.A1(n_1_737_4876), .A2(n_1_737_4875), .B1(n_1_737_5297), 
      .B2(n_1_737_5110), .ZN(n_1_737_4874));
   NOR2_X1 i_1_737_5517 (.A1(n_1_737_5298), .A2(n_1_737_5111), .ZN(n_1_737_4875));
   NOR2_X1 i_1_737_5518 (.A1(n_1_737_148), .A2(n_1_737_5318), .ZN(n_1_737_4876));
   AOI22_X1 i_1_737_5519 (.A1(n_1_737_5094), .A2(n_1_737_4879), .B1(n_1_737_5235), 
      .B2(n_1_737_4878), .ZN(n_1_737_4877));
   OAI21_X1 i_1_737_5520 (.A(n_1_737_5095), .B1(n_1_737_149), .B2(n_1_737_5273), 
      .ZN(n_1_737_4878));
   NOR2_X1 i_1_737_5521 (.A1(n_1_737_149), .A2(n_1_737_5273), .ZN(n_1_737_4879));
   NOR2_X1 i_1_737_5522 (.A1(n_1_737_147), .A2(n_1_737_5357), .ZN(n_1_737_4880));
   AOI21_X1 i_1_737_5523 (.A(n_1_737_5163), .B1(n_1_737_5176), .B2(n_1_737_4882), 
      .ZN(n_640));
   NAND3_X1 i_1_737_5524 (.A1(n_1_737_5176), .A2(n_1_737_4882), .A3(n_1_737_5163), 
      .ZN(n_641));
   NAND2_X1 i_1_737_5525 (.A1(n_1_737_5178), .A2(n_1_737_4882), .ZN(n_1_737_4881));
   INV_X1 i_1_737_5526 (.A(n_1_737_4883), .ZN(n_1_737_4882));
   NOR2_X1 i_1_737_5527 (.A1(n_1_737_5608), .A2(n_1_737_5023), .ZN(n_1_737_4883));
   NAND3_X1 i_1_737_5528 (.A1(n_1_737_4897), .A2(n_1_737_4891), .A3(n_1_737_4884), 
      .ZN(n_642));
   NOR3_X1 i_1_737_5529 (.A1(n_1_737_4906), .A2(n_1_737_4886), .A3(n_1_737_4902), 
      .ZN(n_1_737_4884));
   INV_X1 i_1_737_5530 (.A(n_1_737_4886), .ZN(n_1_737_4885));
   OAI22_X1 i_1_737_5531 (.A1(n_1_737_4888), .A2(n_1_737_4887), .B1(n_1_737_5314), 
      .B2(n_1_737_5298), .ZN(n_1_737_4886));
   NOR2_X1 i_1_737_5532 (.A1(n_1_737_5315), .A2(n_1_737_5297), .ZN(n_1_737_4887));
   NOR2_X1 i_1_737_5533 (.A1(n_1_737_5110), .A2(n_1_737_4890), .ZN(n_1_737_4888));
   INV_X1 i_1_737_5534 (.A(n_1_737_4890), .ZN(n_1_737_4889));
   NOR2_X1 i_1_737_5535 (.A1(n_1_737_5660), .A2(n_1_737_5048), .ZN(n_1_737_4890));
   OAI21_X1 i_1_737_5536 (.A(n_1_737_4892), .B1(n_1_737_5210), .B2(n_1_737_4893), 
      .ZN(n_1_737_4891));
   OAI21_X1 i_1_737_5537 (.A(n_1_737_5190), .B1(n_1_737_5209), .B2(n_1_737_4894), 
      .ZN(n_1_737_4892));
   INV_X1 i_1_737_5538 (.A(n_1_737_4894), .ZN(n_1_737_4893));
   NOR2_X1 i_1_737_5539 (.A1(n_1_737_5121), .A2(n_1_737_4896), .ZN(n_1_737_4894));
   INV_X1 i_1_737_5540 (.A(n_1_737_4896), .ZN(n_1_737_4895));
   NOR2_X1 i_1_737_5541 (.A1(n_1_737_5634), .A2(n_1_737_5039), .ZN(n_1_737_4896));
   OAI21_X1 i_1_737_5542 (.A(n_1_737_4898), .B1(n_1_737_5235), .B2(n_1_737_4899), 
      .ZN(n_1_737_4897));
   OAI21_X1 i_1_737_5543 (.A(n_1_737_5270), .B1(n_1_737_5236), .B2(n_1_737_4900), 
      .ZN(n_1_737_4898));
   INV_X1 i_1_737_5544 (.A(n_1_737_4900), .ZN(n_1_737_4899));
   NOR2_X1 i_1_737_5545 (.A1(n_1_737_5094), .A2(n_1_737_4901), .ZN(n_1_737_4900));
   NOR2_X1 i_1_737_5546 (.A1(n_1_737_5647), .A2(n_1_737_5056), .ZN(n_1_737_4901));
   OAI21_X1 i_1_737_5547 (.A(n_1_737_4903), .B1(n_1_737_5352), .B2(n_1_737_5337), 
      .ZN(n_1_737_4902));
   OAI22_X1 i_1_737_5548 (.A1(n_1_737_5080), .A2(n_1_737_4905), .B1(n_1_737_5353), 
      .B2(n_1_737_5336), .ZN(n_1_737_4903));
   NOR2_X1 i_1_737_5549 (.A1(n_1_737_5333), .A2(n_1_737_4905), .ZN(n_1_737_4904));
   NOR2_X1 i_1_737_5550 (.A1(n_1_737_5667), .A2(n_1_737_5029), .ZN(n_1_737_4905));
   INV_X1 i_1_737_5551 (.A(n_1_737_4907), .ZN(n_1_737_4906));
   OAI21_X1 i_1_737_5552 (.A(n_1_737_4908), .B1(n_1_737_5365), .B2(n_1_737_4909), 
      .ZN(n_1_737_4907));
   OAI21_X1 i_1_737_5553 (.A(n_1_737_5382), .B1(n_1_737_5366), .B2(n_1_737_4910), 
      .ZN(n_1_737_4908));
   INV_X1 i_1_737_5554 (.A(n_1_737_4910), .ZN(n_1_737_4909));
   NOR2_X1 i_1_737_5555 (.A1(n_1_737_5129), .A2(n_1_737_4912), .ZN(n_1_737_4910));
   INV_X1 i_1_737_5556 (.A(n_1_737_4912), .ZN(n_1_737_4911));
   NOR2_X1 i_1_737_5557 (.A1(n_1_737_5621), .A2(n_1_737_5066), .ZN(n_1_737_4912));
   NOR3_X1 i_1_737_5558 (.A1(n_1_737_146), .A2(n_1_737_5151), .A3(n_1_737_4913), 
      .ZN(n_643));
   OAI21_X1 i_1_737_5559 (.A(n_1_737_4913), .B1(n_1_737_146), .B2(n_1_737_5151), 
      .ZN(n_644));
   NOR2_X1 i_1_737_5560 (.A1(n_1_737_4917), .A2(n_1_737_4914), .ZN(n_1_737_4913));
   INV_X1 i_1_737_5561 (.A(n_1_737_4915), .ZN(n_1_737_4914));
   NOR2_X1 i_1_737_5562 (.A1(\out_bs[6] [6]), .A2(\out_bs[6] [5]), .ZN(
      n_1_737_4915));
   INV_X1 i_1_737_5563 (.A(n_1_737_4917), .ZN(n_1_737_4916));
   NAND2_X1 i_1_737_5564 (.A1(n_1_737_5605), .A2(n_1_737_4920), .ZN(n_1_737_4917));
   INV_X1 i_1_737_5565 (.A(n_1_737_4919), .ZN(n_1_737_4918));
   NOR2_X1 i_1_737_5566 (.A1(\out_bs[6] [4]), .A2(n_847), .ZN(n_1_737_4919));
   NOR2_X1 i_1_737_5567 (.A1(n_847), .A2(n_1_737_4921), .ZN(n_1_737_4920));
   AND2_X1 i_1_737_5568 (.A1(n_851), .A2(n_1311), .ZN(n_1_737_4921));
   AOI211_X1 i_1_737_5569 (.A(n_1_737_145), .B(n_1_737_5163), .C1(n_1_737_5182), 
      .C2(n_1_737_4923), .ZN(n_645));
   OAI211_X1 i_1_737_5570 (.A(n_1_737_5182), .B(n_1_737_4923), .C1(n_1_737_145), 
      .C2(n_1_737_5163), .ZN(n_646));
   INV_X1 i_1_737_5571 (.A(n_1_737_4923), .ZN(n_1_737_4922));
   NOR2_X1 i_1_737_5572 (.A1(n_1_737_5177), .A2(n_1_737_4924), .ZN(n_1_737_4923));
   INV_X1 i_1_737_5573 (.A(n_1_737_4925), .ZN(n_1_737_4924));
   NAND2_X1 i_1_737_5574 (.A1(n_849), .A2(n_1313), .ZN(n_1_737_4925));
   NAND3_X1 i_1_737_5575 (.A1(n_1_737_4949), .A2(n_1_737_4926), .A3(n_1_737_4956), 
      .ZN(n_647));
   AOI211_X1 i_1_737_5576 (.A(n_1_737_4935), .B(n_1_737_4928), .C1(n_1_737_4943), 
      .C2(n_1_737_4942), .ZN(n_1_737_4926));
   INV_X1 i_1_737_5577 (.A(n_1_737_4928), .ZN(n_1_737_4927));
   OAI21_X1 i_1_737_5578 (.A(n_1_737_4930), .B1(n_1_737_5298), .B2(n_1_737_4929), 
      .ZN(n_1_737_4928));
   AOI211_X1 i_1_737_5579 (.A(n_1_737_5284), .B(n_1_737_4931), .C1(n_1_737_5592), 
      .C2(n_1_737_5315), .ZN(n_1_737_4929));
   OAI211_X1 i_1_737_5580 (.A(n_1_737_5592), .B(n_1_737_5315), .C1(n_1_737_5284), 
      .C2(n_1_737_4931), .ZN(n_1_737_4930));
   INV_X1 i_1_737_5581 (.A(n_1_737_4932), .ZN(n_1_737_4931));
   NOR2_X1 i_1_737_5582 (.A1(n_1_737_5294), .A2(n_1_737_4933), .ZN(n_1_737_4932));
   NOR2_X1 i_1_737_5583 (.A1(n_1_737_5660), .A2(n_1_737_5659), .ZN(n_1_737_4933));
   INV_X1 i_1_737_5584 (.A(n_1_737_4935), .ZN(n_1_737_4934));
   OAI21_X1 i_1_737_5585 (.A(n_1_737_4937), .B1(n_1_737_5190), .B2(n_1_737_4936), 
      .ZN(n_1_737_4935));
   AOI211_X1 i_1_737_5586 (.A(n_1_737_5221), .B(n_1_737_4938), .C1(n_1_737_5591), 
      .C2(n_1_737_5210), .ZN(n_1_737_4936));
   OAI211_X1 i_1_737_5587 (.A(n_1_737_5591), .B(n_1_737_5210), .C1(n_1_737_5221), 
      .C2(n_1_737_4938), .ZN(n_1_737_4937));
   INV_X1 i_1_737_5588 (.A(n_1_737_4939), .ZN(n_1_737_4938));
   NOR2_X1 i_1_737_5589 (.A1(n_1_737_5230), .A2(n_1_737_4941), .ZN(n_1_737_4939));
   INV_X1 i_1_737_5590 (.A(n_1_737_4941), .ZN(n_1_737_4940));
   NOR2_X1 i_1_737_5591 (.A1(n_1_737_5634), .A2(n_1_737_5633), .ZN(n_1_737_4941));
   NAND2_X1 i_1_737_5592 (.A1(n_1_737_5337), .A2(n_1_737_4944), .ZN(n_1_737_4942));
   OAI22_X1 i_1_737_5593 (.A1(n_1_737_140), .A2(n_1_737_5352), .B1(n_1_737_5337), 
      .B2(n_1_737_4944), .ZN(n_1_737_4943));
   NOR2_X1 i_1_737_5594 (.A1(n_1_737_5083), .A2(n_1_737_4945), .ZN(n_1_737_4944));
   INV_X1 i_1_737_5595 (.A(n_1_737_4946), .ZN(n_1_737_4945));
   NOR2_X1 i_1_737_5596 (.A1(n_1_737_5333), .A2(n_1_737_4948), .ZN(n_1_737_4946));
   INV_X1 i_1_737_5597 (.A(n_1_737_4948), .ZN(n_1_737_4947));
   NOR2_X1 i_1_737_5598 (.A1(n_1_737_5667), .A2(n_1_737_5666), .ZN(n_1_737_4948));
   OAI21_X1 i_1_737_5599 (.A(n_1_737_4950), .B1(n_1_737_5235), .B2(n_1_737_4952), 
      .ZN(n_1_737_4949));
   OAI211_X1 i_1_737_5600 (.A(n_1_737_5253), .B(n_1_737_4953), .C1(n_1_737_5236), 
      .C2(n_1_737_4951), .ZN(n_1_737_4950));
   INV_X1 i_1_737_5601 (.A(n_1_737_4952), .ZN(n_1_737_4951));
   NOR2_X1 i_1_737_5602 (.A1(n_1_737_142), .A2(n_1_737_5270), .ZN(n_1_737_4952));
   NOR2_X1 i_1_737_5603 (.A1(n_1_737_5261), .A2(n_1_737_4955), .ZN(n_1_737_4953));
   INV_X1 i_1_737_5604 (.A(n_1_737_4955), .ZN(n_1_737_4954));
   NOR2_X1 i_1_737_5605 (.A1(n_1_737_5647), .A2(n_1_737_5646), .ZN(n_1_737_4955));
   OAI21_X1 i_1_737_5606 (.A(n_1_737_4957), .B1(n_1_737_5365), .B2(n_1_737_4959), 
      .ZN(n_1_737_4956));
   OAI211_X1 i_1_737_5607 (.A(n_1_737_5393), .B(n_1_737_4960), .C1(n_1_737_5366), 
      .C2(n_1_737_4958), .ZN(n_1_737_4957));
   INV_X1 i_1_737_5608 (.A(n_1_737_4959), .ZN(n_1_737_4958));
   NOR2_X1 i_1_737_5609 (.A1(n_1_737_144), .A2(n_1_737_5382), .ZN(n_1_737_4959));
   NOR2_X1 i_1_737_5610 (.A1(n_1_737_5402), .A2(n_1_737_4962), .ZN(n_1_737_4960));
   INV_X1 i_1_737_5611 (.A(n_1_737_4962), .ZN(n_1_737_4961));
   NOR2_X1 i_1_737_5612 (.A1(n_1_737_5621), .A2(n_1_737_5620), .ZN(n_1_737_4962));
   NOR2_X1 i_1_737_5613 (.A1(n_1_737_139), .A2(n_1_737_5151), .ZN(n_648));
   AOI211_X1 i_1_737_5614 (.A(n_1_737_138), .B(n_1_737_5163), .C1(n_1_737_5176), 
      .C2(n_1_737_4964), .ZN(n_649));
   OAI211_X1 i_1_737_5615 (.A(n_1_737_5176), .B(n_1_737_4964), .C1(n_1_737_138), 
      .C2(n_1_737_5163), .ZN(n_650));
   NAND2_X1 i_1_737_5616 (.A1(n_1_737_5178), .A2(n_1_737_4964), .ZN(n_1_737_4963));
   INV_X1 i_1_737_5617 (.A(n_1_737_4965), .ZN(n_1_737_4964));
   NAND4_X1 i_1_737_5619 (.A1(n_1_737_4988), .A2(n_1_737_4981), .A3(n_1_737_4974), 
      .A4(n_1_737_4966), .ZN(n_651));
   NOR2_X1 i_1_737_5620 (.A1(n_1_737_4994), .A2(n_1_737_4968), .ZN(n_1_737_4966));
   INV_X1 i_1_737_5621 (.A(n_1_737_4968), .ZN(n_1_737_4967));
   OAI21_X1 i_1_737_5622 (.A(n_1_737_4970), .B1(n_1_737_5298), .B2(n_1_737_4969), 
      .ZN(n_1_737_4968));
   AOI211_X1 i_1_737_5623 (.A(n_1_737_5110), .B(n_1_737_4972), .C1(n_1_737_5593), 
      .C2(n_1_737_5315), .ZN(n_1_737_4969));
   OAI211_X1 i_1_737_5624 (.A(n_1_737_5593), .B(n_1_737_5315), .C1(n_1_737_5110), 
      .C2(n_1_737_4972), .ZN(n_1_737_4970));
   INV_X1 i_1_737_5625 (.A(n_1_737_4972), .ZN(n_1_737_4971));
   NOR2_X1 i_1_737_5626 (.A1(n_1_737_5660), .A2(n_1_737_5296), .ZN(n_1_737_4972));
   INV_X1 i_1_737_5627 (.A(n_1_737_4974), .ZN(n_1_737_4973));
   AOI22_X1 i_1_737_5628 (.A1(n_1_737_4977), .A2(n_1_737_4976), .B1(n_1_737_5189), 
      .B2(n_1_737_4975), .ZN(n_1_737_4974));
   OAI21_X1 i_1_737_5629 (.A(n_1_737_4978), .B1(n_1_737_136), .B2(n_1_737_5209), 
      .ZN(n_1_737_4975));
   NOR2_X1 i_1_737_5630 (.A1(n_1_737_136), .A2(n_1_737_5209), .ZN(n_1_737_4976));
   INV_X1 i_1_737_5631 (.A(n_1_737_4978), .ZN(n_1_737_4977));
   NOR2_X1 i_1_737_5632 (.A1(n_1_737_5121), .A2(n_1_737_4980), .ZN(n_1_737_4978));
   INV_X1 i_1_737_5633 (.A(n_1_737_4980), .ZN(n_1_737_4979));
   NOR2_X1 i_1_737_5634 (.A1(n_1_737_5634), .A2(n_1_737_5232), .ZN(n_1_737_4980));
   OAI21_X1 i_1_737_5635 (.A(n_1_737_4982), .B1(n_1_737_5235), .B2(n_1_737_4984), 
      .ZN(n_1_737_4981));
   OAI211_X1 i_1_737_5636 (.A(n_1_737_5095), .B(n_1_737_4986), .C1(n_1_737_5236), 
      .C2(n_1_737_4983), .ZN(n_1_737_4982));
   INV_X1 i_1_737_5637 (.A(n_1_737_4984), .ZN(n_1_737_4983));
   NOR2_X1 i_1_737_5638 (.A1(n_1_737_135), .A2(n_1_737_5270), .ZN(n_1_737_4984));
   NOR2_X1 i_1_737_5639 (.A1(\out_bs[2] [3]), .A2(n_1_737_4987), .ZN(
      n_1_737_4985));
   INV_X1 i_1_737_5640 (.A(n_1_737_4987), .ZN(n_1_737_4986));
   NOR2_X1 i_1_737_5641 (.A1(n_1_737_5647), .A2(n_1_737_5263), .ZN(n_1_737_4987));
   OAI21_X1 i_1_737_5642 (.A(n_1_737_4989), .B1(n_1_737_5336), .B2(n_1_737_4990), 
      .ZN(n_1_737_4988));
   OAI22_X1 i_1_737_5643 (.A1(n_1_737_133), .A2(n_1_737_5352), .B1(n_1_737_5337), 
      .B2(n_1_737_4991), .ZN(n_1_737_4989));
   INV_X1 i_1_737_5644 (.A(n_1_737_4991), .ZN(n_1_737_4990));
   NOR2_X1 i_1_737_5645 (.A1(n_1_737_5080), .A2(n_1_737_4993), .ZN(n_1_737_4991));
   INV_X1 i_1_737_5646 (.A(n_1_737_4993), .ZN(n_1_737_4992));
   NOR2_X1 i_1_737_5647 (.A1(n_1_737_5667), .A2(n_1_737_5335), .ZN(n_1_737_4993));
   INV_X1 i_1_737_5648 (.A(n_1_737_4995), .ZN(n_1_737_4994));
   OAI21_X1 i_1_737_5649 (.A(n_1_737_4996), .B1(n_1_737_5365), .B2(n_1_737_4998), 
      .ZN(n_1_737_4995));
   OAI211_X1 i_1_737_5650 (.A(n_1_737_5130), .B(n_1_737_5000), .C1(n_1_737_5366), 
      .C2(n_1_737_4997), .ZN(n_1_737_4996));
   INV_X1 i_1_737_5651 (.A(n_1_737_4998), .ZN(n_1_737_4997));
   NOR2_X1 i_1_737_5652 (.A1(n_1_737_137), .A2(n_1_737_5382), .ZN(n_1_737_4998));
   NOR2_X1 i_1_737_5653 (.A1(\out_bs[4] [3]), .A2(n_1_737_5001), .ZN(
      n_1_737_4999));
   INV_X1 i_1_737_5654 (.A(n_1_737_5001), .ZN(n_1_737_5000));
   NOR2_X1 i_1_737_5655 (.A1(n_1_737_5621), .A2(n_1_737_5405), .ZN(n_1_737_5001));
   NOR2_X1 i_1_737_5656 (.A1(n_1_737_132), .A2(n_1_737_5151), .ZN(n_652));
   NOR3_X1 i_1_737_5657 (.A1(n_1_737_131), .A2(n_1_737_5163), .A3(n_1_737_5173), 
      .ZN(n_653));
   OAI21_X1 i_1_737_5658 (.A(n_1_737_5173), .B1(n_1_737_131), .B2(n_1_737_5163), 
      .ZN(n_654));
   NAND3_X1 i_1_737_5659 (.A1(n_1_737_5013), .A2(n_1_737_5002), .A3(n_1_737_5017), 
      .ZN(n_655));
   AND3_X1 i_1_737_5660 (.A1(n_1_737_5007), .A2(n_1_737_5004), .A3(n_1_737_5010), 
      .ZN(n_1_737_5002));
   INV_X1 i_1_737_5661 (.A(n_1_737_5004), .ZN(n_1_737_5003));
   OAI22_X1 i_1_737_5662 (.A1(n_1_737_5006), .A2(n_1_737_5005), .B1(n_1_737_5297), 
      .B2(n_1_737_5047), .ZN(n_1_737_5004));
   AND2_X1 i_1_737_5663 (.A1(n_1_737_5297), .A2(n_1_737_5047), .ZN(n_1_737_5005));
   NOR2_X1 i_1_737_5664 (.A1(n_1_737_127), .A2(n_1_737_5314), .ZN(n_1_737_5006));
   AOI22_X1 i_1_737_5665 (.A1(n_1_737_5037), .A2(n_1_737_5009), .B1(n_1_737_5189), 
      .B2(n_1_737_5008), .ZN(n_1_737_5007));
   OAI21_X1 i_1_737_5666 (.A(n_1_737_5038), .B1(n_1_737_129), .B2(n_1_737_5209), 
      .ZN(n_1_737_5008));
   NOR2_X1 i_1_737_5667 (.A1(n_1_737_129), .A2(n_1_737_5209), .ZN(n_1_737_5009));
   OAI22_X1 i_1_737_5668 (.A1(n_1_737_5055), .A2(n_1_737_5011), .B1(n_1_737_5235), 
      .B2(n_1_737_5012), .ZN(n_1_737_5010));
   AND2_X1 i_1_737_5669 (.A1(n_1_737_5235), .A2(n_1_737_5012), .ZN(n_1_737_5011));
   NOR2_X1 i_1_737_5670 (.A1(n_1_737_128), .A2(n_1_737_5270), .ZN(n_1_737_5012));
   OAI21_X1 i_1_737_5671 (.A(n_1_737_5014), .B1(n_1_737_5336), .B2(n_1_737_5016), 
      .ZN(n_1_737_5013));
   OAI22_X1 i_1_737_5672 (.A1(n_1_737_126), .A2(n_1_737_5352), .B1(n_1_737_5337), 
      .B2(n_1_737_5015), .ZN(n_1_737_5014));
   INV_X1 i_1_737_5673 (.A(n_1_737_5016), .ZN(n_1_737_5015));
   NAND2_X1 i_1_737_5674 (.A1(n_1_737_5671), .A2(n_1_737_5327), .ZN(n_1_737_5016));
   OAI22_X1 i_1_737_5675 (.A1(n_1_737_5064), .A2(n_1_737_5018), .B1(n_1_737_5365), 
      .B2(n_1_737_5019), .ZN(n_1_737_5017));
   AND2_X1 i_1_737_5676 (.A1(n_1_737_5365), .A2(n_1_737_5019), .ZN(n_1_737_5018));
   NOR2_X1 i_1_737_5677 (.A1(n_1_737_130), .A2(n_1_737_5382), .ZN(n_1_737_5019));
   AOI211_X1 i_1_737_5678 (.A(\out_as[5] [6]), .B(n_1_737_5070), .C1(
      n_1_737_5180), .C2(n_1_737_5021), .ZN(n_656));
   OAI211_X1 i_1_737_5679 (.A(n_1_737_5180), .B(n_1_737_5021), .C1(
      \out_as[5] [6]), .C2(n_1_737_5070), .ZN(n_657));
   INV_X1 i_1_737_5680 (.A(n_1_737_5021), .ZN(n_1_737_5020));
   NOR2_X1 i_1_737_5681 (.A1(n_1_737_5174), .A2(n_1_737_5022), .ZN(n_1_737_5021));
   INV_X1 i_1_737_5682 (.A(n_1_737_5023), .ZN(n_1_737_5022));
   NAND2_X1 i_1_737_5683 (.A1(n_1313), .A2(\out_bs[5] [0]), .ZN(n_1_737_5023));
   NAND3_X1 i_1_737_5684 (.A1(n_1_737_5049), .A2(n_1_737_5031), .A3(n_1_737_5024), 
      .ZN(n_658));
   NOR3_X1 i_1_737_5685 (.A1(n_1_737_5042), .A2(n_1_737_5025), .A3(n_1_737_5059), 
      .ZN(n_1_737_5024));
   OAI21_X1 i_1_737_5686 (.A(n_1_737_5026), .B1(n_1_737_5337), .B2(n_1_737_5086), 
      .ZN(n_1_737_5025));
   OAI22_X1 i_1_737_5687 (.A1(n_1_737_5082), .A2(n_1_737_5027), .B1(n_1_737_5336), 
      .B2(n_1_737_5087), .ZN(n_1_737_5026));
   INV_X1 i_1_737_5688 (.A(n_1_737_5028), .ZN(n_1_737_5027));
   NOR2_X1 i_1_737_5689 (.A1(n_1_737_5328), .A2(n_1_737_5030), .ZN(n_1_737_5028));
   INV_X1 i_1_737_5690 (.A(n_1_737_5030), .ZN(n_1_737_5029));
   NOR2_X1 i_1_737_5691 (.A1(n_1_737_5666), .A2(n_1_737_5665), .ZN(n_1_737_5030));
   OAI21_X1 i_1_737_5692 (.A(n_1_737_5032), .B1(n_1_737_5189), .B2(n_1_737_5033), 
      .ZN(n_1_737_5031));
   OAI21_X1 i_1_737_5693 (.A(n_1_737_5117), .B1(n_1_737_5190), .B2(n_1_737_5034), 
      .ZN(n_1_737_5032));
   INV_X1 i_1_737_5694 (.A(n_1_737_5034), .ZN(n_1_737_5033));
   NOR2_X1 i_1_737_5695 (.A1(n_1_737_5219), .A2(n_1_737_5035), .ZN(n_1_737_5034));
   INV_X1 i_1_737_5696 (.A(n_1_737_5036), .ZN(n_1_737_5035));
   NOR2_X1 i_1_737_5697 (.A1(n_1_737_5224), .A2(n_1_737_5040), .ZN(n_1_737_5036));
   INV_X1 i_1_737_5698 (.A(n_1_737_5038), .ZN(n_1_737_5037));
   NOR2_X1 i_1_737_5699 (.A1(n_1_737_5224), .A2(n_1_737_5219), .ZN(n_1_737_5038));
   INV_X1 i_1_737_5700 (.A(n_1_737_5040), .ZN(n_1_737_5039));
   NOR2_X1 i_1_737_5701 (.A1(n_1_737_5633), .A2(n_1_737_5632), .ZN(n_1_737_5040));
   INV_X1 i_1_737_5702 (.A(n_1_737_5042), .ZN(n_1_737_5041));
   OAI22_X1 i_1_737_5703 (.A1(n_1_737_5044), .A2(n_1_737_5043), .B1(n_1_737_5298), 
      .B2(n_1_737_5106), .ZN(n_1_737_5042));
   NOR2_X1 i_1_737_5704 (.A1(n_1_737_5297), .A2(n_1_737_5107), .ZN(n_1_737_5043));
   NOR2_X1 i_1_737_5705 (.A1(n_1_737_5282), .A2(n_1_737_5046), .ZN(n_1_737_5044));
   INV_X1 i_1_737_5706 (.A(n_1_737_5046), .ZN(n_1_737_5045));
   NAND2_X1 i_1_737_5707 (.A1(n_1_737_5289), .A2(n_1_737_5048), .ZN(n_1_737_5046));
   NAND2_X1 i_1_737_5708 (.A1(n_1_737_5664), .A2(n_1_737_5288), .ZN(n_1_737_5047));
   NAND2_X1 i_1_737_5709 (.A1(\out_bs[1] [1]), .A2(\out_bs[1] [0]), .ZN(
      n_1_737_5048));
   AOI21_X1 i_1_737_5710 (.A(n_1_737_5050), .B1(n_1_737_5100), .B2(n_1_737_5051), 
      .ZN(n_1_737_5049));
   AOI21_X1 i_1_737_5711 (.A(n_1_737_5236), .B1(n_1_737_5099), .B2(n_1_737_5052), 
      .ZN(n_1_737_5050));
   INV_X1 i_1_737_5712 (.A(n_1_737_5052), .ZN(n_1_737_5051));
   NOR2_X1 i_1_737_5713 (.A1(n_1_737_5250), .A2(n_1_737_5053), .ZN(n_1_737_5052));
   INV_X1 i_1_737_5714 (.A(n_1_737_5054), .ZN(n_1_737_5053));
   NOR2_X1 i_1_737_5715 (.A1(n_1_737_5256), .A2(n_1_737_5057), .ZN(n_1_737_5054));
   NAND2_X1 i_1_737_5716 (.A1(n_1_737_5651), .A2(n_1_737_5255), .ZN(n_1_737_5055));
   INV_X1 i_1_737_5717 (.A(n_1_737_5057), .ZN(n_1_737_5056));
   NOR2_X1 i_1_737_5718 (.A1(n_1_737_5646), .A2(n_1_737_5645), .ZN(n_1_737_5057));
   INV_X1 i_1_737_5719 (.A(n_1_737_5059), .ZN(n_1_737_5058));
   OAI22_X1 i_1_737_5720 (.A1(n_1_737_5061), .A2(n_1_737_5060), .B1(n_1_737_5366), 
      .B2(n_1_737_5134), .ZN(n_1_737_5059));
   NOR2_X1 i_1_737_5721 (.A1(n_1_737_5365), .A2(n_1_737_5135), .ZN(n_1_737_5060));
   NOR2_X1 i_1_737_5722 (.A1(n_1_737_5390), .A2(n_1_737_5062), .ZN(n_1_737_5061));
   INV_X1 i_1_737_5723 (.A(n_1_737_5063), .ZN(n_1_737_5062));
   NOR2_X1 i_1_737_5724 (.A1(n_1_737_5397), .A2(n_1_737_5065), .ZN(n_1_737_5063));
   NAND2_X1 i_1_737_5725 (.A1(n_1_737_5625), .A2(n_1_737_5396), .ZN(n_1_737_5064));
   INV_X1 i_1_737_5726 (.A(n_1_737_5066), .ZN(n_1_737_5065));
   NAND2_X1 i_1_737_5727 (.A1(\out_bs[4] [1]), .A2(\out_bs[4] [0]), .ZN(
      n_1_737_5066));
   NOR3_X1 i_1_737_5728 (.A1(\out_as[6] [6]), .A2(n_1_737_5067), .A3(n_1_737_125), 
      .ZN(n_659));
   NOR2_X1 i_1_737_5729 (.A1(\out_as[6] [6]), .A2(n_1_737_5067), .ZN(n_660));
   OR2_X1 i_1_737_5730 (.A1(\out_as[6] [5]), .A2(n_1_737_5148), .ZN(n_1_737_5067));
   INV_X1 i_1_737_5731 (.A(n_1_737_5068), .ZN(n_661));
   OAI21_X1 i_1_737_5732 (.A(n_1_737_5069), .B1(n_1_737_5181), .B2(n_1_737_5071), 
      .ZN(n_1_737_5068));
   OR3_X1 i_1_737_5733 (.A1(n_1_737_5181), .A2(n_1_737_5071), .A3(n_1_737_5069), 
      .ZN(n_662));
   NOR3_X1 i_1_737_5734 (.A1(\out_as[5] [6]), .A2(n_1_737_5070), .A3(n_1_737_124), 
      .ZN(n_1_737_5069));
   OR2_X1 i_1_737_5735 (.A1(\out_as[5] [5]), .A2(n_1_737_5160), .ZN(n_1_737_5070));
   INV_X1 i_1_737_5736 (.A(n_1_737_5072), .ZN(n_1_737_5071));
   NOR2_X1 i_1_737_5737 (.A1(n_1_737_5177), .A2(n_1_737_5073), .ZN(n_1_737_5072));
   INV_X1 i_1_737_5738 (.A(n_1_737_5074), .ZN(n_1_737_5073));
   NOR2_X1 i_1_737_5739 (.A1(n_849), .A2(n_1313), .ZN(n_1_737_5074));
   NAND4_X1 i_1_737_5740 (.A1(n_1_737_5114), .A2(n_1_737_5103), .A3(n_1_737_5075), 
      .A4(n_1_737_5125), .ZN(n_663));
   AOI21_X1 i_1_737_5741 (.A(n_1_737_5089), .B1(n_1_737_5077), .B2(n_1_737_5076), 
      .ZN(n_1_737_5075));
   NAND2_X1 i_1_737_5742 (.A1(n_1_737_5337), .A2(n_1_737_5078), .ZN(n_1_737_5076));
   OAI22_X1 i_1_737_5743 (.A1(n_1_737_119), .A2(n_1_737_5086), .B1(n_1_737_5337), 
      .B2(n_1_737_5078), .ZN(n_1_737_5077));
   NOR2_X1 i_1_737_5744 (.A1(n_1_737_5084), .A2(n_1_737_5080), .ZN(n_1_737_5078));
   NOR2_X1 i_1_737_5745 (.A1(n_1_737_5333), .A2(n_1_737_5084), .ZN(n_1_737_5079));
   INV_X1 i_1_737_5746 (.A(n_1_737_5081), .ZN(n_1_737_5080));
   NOR2_X1 i_1_737_5747 (.A1(\out_bs[0] [6]), .A2(n_1_737_5330), .ZN(
      n_1_737_5081));
   NAND2_X1 i_1_737_5748 (.A1(n_1_737_5671), .A2(n_1_737_5332), .ZN(n_1_737_5082));
   NAND2_X1 i_1_737_5749 (.A1(n_1_737_5671), .A2(n_1_737_5670), .ZN(n_1_737_5083));
   INV_X1 i_1_737_5750 (.A(n_1_737_5085), .ZN(n_1_737_5084));
   NOR2_X1 i_1_737_5751 (.A1(\out_bs[0] [2]), .A2(\out_bs[0] [1]), .ZN(
      n_1_737_5085));
   INV_X1 i_1_737_5752 (.A(n_1_737_5087), .ZN(n_1_737_5086));
   NOR2_X1 i_1_737_5753 (.A1(\out_as[0] [6]), .A2(n_1_737_5088), .ZN(
      n_1_737_5087));
   OR2_X1 i_1_737_5754 (.A1(\out_as[0] [5]), .A2(n_1_737_5349), .ZN(n_1_737_5088));
   INV_X1 i_1_737_5755 (.A(n_1_737_5090), .ZN(n_1_737_5089));
   OAI22_X1 i_1_737_5756 (.A1(n_1_737_5098), .A2(n_1_737_5091), .B1(n_1_737_5235), 
      .B2(n_1_737_5092), .ZN(n_1_737_5090));
   AND2_X1 i_1_737_5757 (.A1(n_1_737_5235), .A2(n_1_737_5092), .ZN(n_1_737_5091));
   NAND2_X1 i_1_737_5758 (.A1(n_1_737_5253), .A2(n_1_737_5093), .ZN(n_1_737_5092));
   NOR2_X1 i_1_737_5759 (.A1(n_1_737_5261), .A2(n_1_737_5096), .ZN(n_1_737_5093));
   INV_X1 i_1_737_5760 (.A(n_1_737_5095), .ZN(n_1_737_5094));
   NOR2_X1 i_1_737_5761 (.A1(\out_bs[2] [6]), .A2(n_1_737_5258), .ZN(
      n_1_737_5095));
   INV_X1 i_1_737_5762 (.A(n_1_737_5097), .ZN(n_1_737_5096));
   NOR2_X1 i_1_737_5763 (.A1(\out_bs[2] [2]), .A2(\out_bs[2] [1]), .ZN(
      n_1_737_5097));
   NOR2_X1 i_1_737_5764 (.A1(n_1_737_121), .A2(n_1_737_5099), .ZN(n_1_737_5098));
   INV_X1 i_1_737_5765 (.A(n_1_737_5100), .ZN(n_1_737_5099));
   NOR2_X1 i_1_737_5766 (.A1(\out_as[2] [6]), .A2(n_1_737_5101), .ZN(
      n_1_737_5100));
   OR2_X1 i_1_737_5767 (.A1(\out_as[2] [5]), .A2(n_1_737_5267), .ZN(n_1_737_5101));
   INV_X1 i_1_737_5768 (.A(n_1_737_5103), .ZN(n_1_737_5102));
   AOI21_X1 i_1_737_5769 (.A(n_1_737_5105), .B1(n_1_737_5297), .B2(n_1_737_5104), 
      .ZN(n_1_737_5103));
   OAI211_X1 i_1_737_5770 (.A(n_1_737_5285), .B(n_1_737_5109), .C1(n_1_737_120), 
      .C2(n_1_737_5106), .ZN(n_1_737_5104));
   AOI211_X1 i_1_737_5771 (.A(n_1_737_120), .B(n_1_737_5106), .C1(n_1_737_5285), 
      .C2(n_1_737_5109), .ZN(n_1_737_5105));
   INV_X1 i_1_737_5772 (.A(n_1_737_5107), .ZN(n_1_737_5106));
   NOR2_X1 i_1_737_5773 (.A1(\out_as[1] [6]), .A2(n_1_737_5108), .ZN(
      n_1_737_5107));
   OR2_X1 i_1_737_5774 (.A1(\out_as[1] [5]), .A2(n_1_737_5311), .ZN(n_1_737_5108));
   NOR2_X1 i_1_737_5775 (.A1(n_1_737_5294), .A2(n_1_737_5112), .ZN(n_1_737_5109));
   INV_X1 i_1_737_5776 (.A(n_1_737_5111), .ZN(n_1_737_5110));
   NOR2_X1 i_1_737_5777 (.A1(\out_bs[1] [6]), .A2(n_1_737_5290), .ZN(
      n_1_737_5111));
   INV_X1 i_1_737_5778 (.A(n_1_737_5113), .ZN(n_1_737_5112));
   NOR2_X1 i_1_737_5779 (.A1(\out_bs[1] [2]), .A2(\out_bs[1] [1]), .ZN(
      n_1_737_5113));
   OAI22_X1 i_1_737_5780 (.A1(n_1_737_5119), .A2(n_1_737_5115), .B1(n_1_737_5189), 
      .B2(n_1_737_5116), .ZN(n_1_737_5114));
   AND2_X1 i_1_737_5781 (.A1(n_1_737_5189), .A2(n_1_737_5116), .ZN(n_1_737_5115));
   NOR2_X1 i_1_737_5782 (.A1(n_1_737_122), .A2(n_1_737_5117), .ZN(n_1_737_5116));
   OR2_X1 i_1_737_5783 (.A1(\out_as[3] [6]), .A2(n_1_737_5118), .ZN(n_1_737_5117));
   OR2_X1 i_1_737_5784 (.A1(\out_as[3] [5]), .A2(n_1_737_5206), .ZN(n_1_737_5118));
   NAND2_X1 i_1_737_5785 (.A1(n_1_737_5222), .A2(n_1_737_5120), .ZN(n_1_737_5119));
   NOR2_X1 i_1_737_5786 (.A1(n_1_737_5230), .A2(n_1_737_5123), .ZN(n_1_737_5120));
   INV_X1 i_1_737_5787 (.A(n_1_737_5122), .ZN(n_1_737_5121));
   NOR2_X1 i_1_737_5788 (.A1(\out_bs[3] [6]), .A2(n_1_737_5226), .ZN(
      n_1_737_5122));
   INV_X1 i_1_737_5789 (.A(n_1_737_5124), .ZN(n_1_737_5123));
   NOR2_X1 i_1_737_5790 (.A1(\out_bs[3] [2]), .A2(\out_bs[3] [1]), .ZN(
      n_1_737_5124));
   OAI22_X1 i_1_737_5791 (.A1(n_1_737_5133), .A2(n_1_737_5126), .B1(n_1_737_5365), 
      .B2(n_1_737_5127), .ZN(n_1_737_5125));
   AND2_X1 i_1_737_5792 (.A1(n_1_737_5365), .A2(n_1_737_5127), .ZN(n_1_737_5126));
   NAND2_X1 i_1_737_5793 (.A1(n_1_737_5393), .A2(n_1_737_5128), .ZN(n_1_737_5127));
   NOR2_X1 i_1_737_5794 (.A1(n_1_737_5402), .A2(n_1_737_5131), .ZN(n_1_737_5128));
   INV_X1 i_1_737_5795 (.A(n_1_737_5130), .ZN(n_1_737_5129));
   NOR2_X1 i_1_737_5796 (.A1(\out_bs[4] [6]), .A2(n_1_737_5399), .ZN(
      n_1_737_5130));
   INV_X1 i_1_737_5797 (.A(n_1_737_5132), .ZN(n_1_737_5131));
   NOR2_X1 i_1_737_5798 (.A1(\out_bs[4] [2]), .A2(\out_bs[4] [1]), .ZN(
      n_1_737_5132));
   NOR2_X1 i_1_737_5799 (.A1(n_1_737_123), .A2(n_1_737_5134), .ZN(n_1_737_5133));
   INV_X1 i_1_737_5800 (.A(n_1_737_5135), .ZN(n_1_737_5134));
   NOR2_X1 i_1_737_5801 (.A1(\out_as[4] [6]), .A2(n_1_737_5136), .ZN(
      n_1_737_5135));
   OR2_X1 i_1_737_5802 (.A1(\out_as[4] [5]), .A2(n_1_737_5379), .ZN(n_1_737_5136));
   OR2_X1 i_1_737_5803 (.A1(n_958), .A2(n_771), .ZN(n_664));
   OR2_X1 i_1_737_5804 (.A1(n_953), .A2(n_772), .ZN(n_665));
   OR2_X1 i_1_737_5805 (.A1(n_963), .A2(n_773), .ZN(n_666));
   OR2_X1 i_1_737_5806 (.A1(n_954), .A2(n_776), .ZN(n_667));
   OR2_X1 i_1_737_5807 (.A1(n_966), .A2(n_777), .ZN(n_668));
   OR2_X1 i_1_737_5808 (.A1(n_959), .A2(n_779), .ZN(n_669));
   OR2_X1 i_1_737_5810 (.A1(n_964), .A2(n_780), .ZN(n_670));
   OR2_X1 i_1_737_5811 (.A1(n_956), .A2(n_781), .ZN(n_671));
   OR2_X1 i_1_737_5812 (.A1(n_960), .A2(n_782), .ZN(n_672));
   OR2_X1 i_1_737_5813 (.A1(n_967), .A2(n_784), .ZN(n_673));
   OR2_X1 i_1_737_5814 (.A1(n_965), .A2(n_788), .ZN(n_674));
   OR2_X1 i_1_737_5815 (.A1(n_961), .A2(n_790), .ZN(n_675));
   OR2_X1 i_1_737_5816 (.A1(n_957), .A2(n_793), .ZN(n_676));
   OR2_X1 i_1_737_5818 (.A1(n_968), .A2(n_815), .ZN(n_677));
   NOR2_X1 i_1_737_5820 (.A1(\out_as[7] [6]), .A2(n_1_737_117), .ZN(n_678));
   NOR2_X1 i_1_737_5821 (.A1(\out_as[7] [6]), .A2(n_1_737_111), .ZN(n_679));
   NOR2_X1 i_1_737_5822 (.A1(\out_as[7] [6]), .A2(n_1_737_106), .ZN(n_680));
   NOR2_X1 i_1_737_5823 (.A1(\out_as[7] [6]), .A2(n_1_737_101), .ZN(n_681));
   NOR2_X1 i_1_737_5824 (.A1(\out_as[7] [6]), .A2(n_1_737_97), .ZN(n_682));
   NOR2_X1 i_1_737_5825 (.A1(\out_as[7] [6]), .A2(n_1_737_93), .ZN(n_683));
   NOR2_X1 i_1_737_5826 (.A1(\out_as[7] [6]), .A2(n_1_737_89), .ZN(n_684));
   NOR2_X1 i_1_737_5827 (.A1(\out_as[7] [6]), .A2(n_1_737_85), .ZN(n_685));
   NOR2_X1 i_1_737_5828 (.A1(\out_as[7] [6]), .A2(n_1_737_82), .ZN(n_686));
   NOR2_X1 i_1_737_5829 (.A1(\out_as[7] [6]), .A2(n_1_737_79), .ZN(n_687));
   NOR2_X1 i_1_737_5830 (.A1(\out_as[7] [6]), .A2(n_1_737_76), .ZN(n_688));
   NOR2_X1 i_1_737_5831 (.A1(\out_as[7] [6]), .A2(n_1_737_73), .ZN(n_689));
   NOR2_X1 i_1_737_5832 (.A1(\out_as[7] [6]), .A2(n_1_737_70), .ZN(n_690));
   NOR2_X1 i_1_737_5833 (.A1(\out_as[7] [6]), .A2(n_1_737_67), .ZN(n_691));
   NOR2_X1 i_1_737_5834 (.A1(\out_as[7] [6]), .A2(n_1_737_64), .ZN(n_692));
   NOR2_X1 i_1_737_5835 (.A1(\out_as[7] [6]), .A2(n_1_737_61), .ZN(n_693));
   NOR2_X1 i_1_737_5836 (.A1(\out_as[7] [6]), .A2(n_1_737_59), .ZN(n_694));
   NOR2_X1 i_1_737_5837 (.A1(\out_as[7] [6]), .A2(n_1_737_57), .ZN(n_695));
   NOR2_X1 i_1_737_5838 (.A1(\out_as[7] [6]), .A2(n_1_737_55), .ZN(n_696));
   NOR2_X1 i_1_737_5839 (.A1(\out_as[7] [6]), .A2(n_1_737_53), .ZN(n_697));
   NOR2_X1 i_1_737_5840 (.A1(\out_as[7] [6]), .A2(n_1_737_51), .ZN(n_698));
   NOR2_X1 i_1_737_5841 (.A1(\out_as[7] [6]), .A2(n_1_737_49), .ZN(n_699));
   NOR2_X1 i_1_737_5842 (.A1(\out_as[7] [6]), .A2(n_1_737_47), .ZN(n_700));
   NOR2_X1 i_1_737_5843 (.A1(\out_as[7] [6]), .A2(n_1_737_45), .ZN(n_701));
   NOR2_X1 i_1_737_5844 (.A1(\out_as[7] [6]), .A2(n_1_737_43), .ZN(n_702));
   NOR2_X1 i_1_737_5845 (.A1(\out_as[7] [6]), .A2(n_1_737_41), .ZN(n_703));
   NOR2_X1 i_1_737_5846 (.A1(\out_as[7] [6]), .A2(n_1_737_39), .ZN(n_704));
   NOR2_X1 i_1_737_5847 (.A1(\out_as[7] [6]), .A2(n_1_737_37), .ZN(n_705));
   NOR2_X1 i_1_737_5848 (.A1(\out_as[7] [6]), .A2(n_1_737_35), .ZN(n_706));
   NOR2_X1 i_1_737_5849 (.A1(\out_as[7] [6]), .A2(n_1_737_33), .ZN(n_707));
   OR2_X1 i_1_737_5850 (.A1(n_969), .A2(n_709), .ZN(n_708));
   NOR2_X1 i_1_737_5851 (.A1(\out_as[7] [6]), .A2(n_1_737_31), .ZN(n_709));
   NOR2_X1 i_1_737_5852 (.A1(n_1_737_116), .A2(n_1_737_5140), .ZN(n_710));
   NOR2_X1 i_1_737_5853 (.A1(n_1_737_110), .A2(n_1_737_5140), .ZN(n_711));
   NOR2_X1 i_1_737_5854 (.A1(n_1_737_105), .A2(n_1_737_5140), .ZN(n_712));
   NOR2_X1 i_1_737_5855 (.A1(n_1_737_100), .A2(n_1_737_5140), .ZN(n_713));
   NOR2_X1 i_1_737_5856 (.A1(n_1_737_96), .A2(n_1_737_5140), .ZN(n_714));
   NOR2_X1 i_1_737_5857 (.A1(n_1_737_92), .A2(n_1_737_5140), .ZN(n_715));
   NOR2_X1 i_1_737_5858 (.A1(n_1_737_88), .A2(n_1_737_5140), .ZN(n_716));
   NOR2_X1 i_1_737_5859 (.A1(n_1_737_84), .A2(n_1_737_5140), .ZN(n_717));
   NOR2_X1 i_1_737_5860 (.A1(n_1_737_81), .A2(n_1_737_5140), .ZN(n_718));
   NOR2_X1 i_1_737_5861 (.A1(n_1_737_78), .A2(n_1_737_5140), .ZN(n_719));
   NOR2_X1 i_1_737_5862 (.A1(n_1_737_75), .A2(n_1_737_5140), .ZN(n_720));
   NOR2_X1 i_1_737_5863 (.A1(n_1_737_72), .A2(n_1_737_5140), .ZN(n_721));
   NOR2_X1 i_1_737_5864 (.A1(n_1_737_69), .A2(n_1_737_5140), .ZN(n_722));
   NOR2_X1 i_1_737_5865 (.A1(n_1_737_66), .A2(n_1_737_5140), .ZN(n_723));
   NOR2_X1 i_1_737_5866 (.A1(n_1_737_63), .A2(n_1_737_5140), .ZN(n_724));
   NOR2_X1 i_1_737_5867 (.A1(n_1_737_115), .A2(n_1_737_5139), .ZN(n_725));
   NOR2_X1 i_1_737_5868 (.A1(n_1_737_109), .A2(n_1_737_5139), .ZN(n_726));
   NOR2_X1 i_1_737_5869 (.A1(n_1_737_104), .A2(n_1_737_5139), .ZN(n_727));
   NOR2_X1 i_1_737_5870 (.A1(n_1_737_99), .A2(n_1_737_5139), .ZN(n_728));
   NOR2_X1 i_1_737_5871 (.A1(n_1_737_95), .A2(n_1_737_5139), .ZN(n_729));
   NOR2_X1 i_1_737_5872 (.A1(n_1_737_91), .A2(n_1_737_5139), .ZN(n_730));
   NOR2_X1 i_1_737_5873 (.A1(n_1_737_87), .A2(n_1_737_5139), .ZN(n_731));
   NOR2_X1 i_1_737_5874 (.A1(n_1_737_114), .A2(n_1_737_5137), .ZN(n_732));
   NOR2_X1 i_1_737_5875 (.A1(n_1_737_108), .A2(n_1_737_5137), .ZN(n_733));
   NOR2_X1 i_1_737_5876 (.A1(n_1_737_103), .A2(n_1_737_5137), .ZN(n_734));
   INV_X1 i_1_737_5877 (.A(n_735), .ZN(n_1_737_5137));
   NOR2_X1 i_1_737_5878 (.A1(\out_as[7] [6]), .A2(n_1_737_5138), .ZN(n_735));
   OR2_X1 i_1_737_5879 (.A1(\out_as[7] [5]), .A2(n_1_737_5144), .ZN(n_1_737_5138));
   NOR3_X1 i_1_737_5880 (.A1(n_1_737_113), .A2(n_1_737_5141), .A3(\out_as[7] [6]), 
      .ZN(n_736));
   INV_X1 i_1_737_5881 (.A(n_737), .ZN(n_1_737_5139));
   NOR2_X1 i_1_737_5882 (.A1(\out_as[7] [6]), .A2(n_1_737_5142), .ZN(n_737));
   INV_X1 i_1_737_5883 (.A(n_738), .ZN(n_1_737_5140));
   NOR2_X1 i_1_737_5884 (.A1(\out_as[7] [6]), .A2(\out_as[7] [5]), .ZN(n_738));
   OR2_X1 i_1_737_5885 (.A1(\out_as[7] [5]), .A2(n_1_737_5143), .ZN(n_1_737_5141));
   OR2_X1 i_1_737_5886 (.A1(\out_as[7] [5]), .A2(\out_as[7] [4]), .ZN(
      n_1_737_5142));
   OR2_X1 i_1_737_5887 (.A1(\out_as[7] [4]), .A2(n_1_737_5145), .ZN(n_1_737_5143));
   OR2_X1 i_1_737_5888 (.A1(\out_as[7] [4]), .A2(\out_as[7] [3]), .ZN(
      n_1_737_5144));
   OR2_X1 i_1_737_5889 (.A1(\out_as[7] [3]), .A2(\out_as[7] [2]), .ZN(
      n_1_737_5145));
   NOR2_X1 i_1_737_5890 (.A1(\out_as[6] [6]), .A2(n_1_737_5146), .ZN(n_739));
   OR2_X1 i_1_737_5891 (.A1(\out_as[6] [5]), .A2(n_1_737_5147), .ZN(n_1_737_5146));
   OR2_X1 i_1_737_5892 (.A1(\out_as[6] [4]), .A2(n_1_737_5149), .ZN(n_1_737_5147));
   OR2_X1 i_1_737_5893 (.A1(\out_as[6] [4]), .A2(n_1_737_5150), .ZN(n_1_737_5148));
   OR2_X1 i_1_737_5894 (.A1(\out_as[6] [3]), .A2(n_1_737_5157), .ZN(n_1_737_5149));
   OR2_X1 i_1_737_5895 (.A1(\out_as[6] [3]), .A2(\out_as[6] [2]), .ZN(
      n_1_737_5150));
   INV_X1 i_1_737_5896 (.A(n_740), .ZN(n_1_737_5151));
   NOR2_X1 i_1_737_5897 (.A1(\out_as[6] [6]), .A2(n_1_737_5152), .ZN(n_740));
   OR2_X1 i_1_737_5898 (.A1(\out_as[6] [5]), .A2(n_1_737_5153), .ZN(n_1_737_5152));
   OR2_X1 i_1_737_5899 (.A1(\out_as[6] [4]), .A2(\out_as[6] [3]), .ZN(
      n_1_737_5153));
   INV_X1 i_1_737_5900 (.A(n_741), .ZN(n_1_737_5154));
   NOR2_X1 i_1_737_5901 (.A1(\out_as[6] [6]), .A2(n_1_737_5156), .ZN(n_741));
   INV_X1 i_1_737_5902 (.A(n_742), .ZN(n_1_737_5155));
   NOR2_X1 i_1_737_5903 (.A1(\out_as[6] [6]), .A2(\out_as[6] [5]), .ZN(n_742));
   OR2_X1 i_1_737_5904 (.A1(\out_as[6] [5]), .A2(\out_as[6] [4]), .ZN(
      n_1_737_5156));
   OR2_X1 i_1_737_5905 (.A1(\out_as[6] [2]), .A2(\out_as[6] [1]), .ZN(
      n_1_737_5157));
   AOI211_X1 i_1_737_5906 (.A(\out_as[5] [6]), .B(n_1_737_5158), .C1(
      n_1_737_5180), .C2(n_1_737_5171), .ZN(n_743));
   OAI211_X1 i_1_737_5907 (.A(n_1_737_5180), .B(n_1_737_5171), .C1(
      \out_as[5] [6]), .C2(n_1_737_5158), .ZN(n_744));
   OR2_X1 i_1_737_5908 (.A1(\out_as[5] [5]), .A2(n_1_737_5159), .ZN(n_1_737_5158));
   OR2_X1 i_1_737_5909 (.A1(\out_as[5] [4]), .A2(n_1_737_5161), .ZN(n_1_737_5159));
   OR2_X1 i_1_737_5910 (.A1(\out_as[5] [4]), .A2(n_1_737_5162), .ZN(n_1_737_5160));
   OR2_X1 i_1_737_5911 (.A1(\out_as[5] [3]), .A2(n_1_737_5170), .ZN(n_1_737_5161));
   OR2_X1 i_1_737_5912 (.A1(\out_as[5] [3]), .A2(\out_as[5] [2]), .ZN(
      n_1_737_5162));
   OR2_X1 i_1_737_5913 (.A1(\out_as[5] [6]), .A2(n_1_737_5164), .ZN(n_1_737_5163));
   OR2_X1 i_1_737_5914 (.A1(\out_as[5] [5]), .A2(n_1_737_5165), .ZN(n_1_737_5164));
   OR2_X1 i_1_737_5915 (.A1(\out_as[5] [4]), .A2(\out_as[5] [3]), .ZN(
      n_1_737_5165));
   OR2_X1 i_1_737_5916 (.A1(\out_as[5] [6]), .A2(n_1_737_5169), .ZN(n_1_737_5166));
   NOR2_X1 i_1_737_5918 (.A1(\out_as[5] [6]), .A2(\out_as[5] [5]), .ZN(
      n_1_737_5168));
   OR2_X1 i_1_737_5919 (.A1(\out_as[5] [5]), .A2(\out_as[5] [4]), .ZN(
      n_1_737_5169));
   OR2_X1 i_1_737_5920 (.A1(\out_as[5] [2]), .A2(\out_as[5] [1]), .ZN(
      n_1_737_5170));
   INV_X1 i_1_737_5921 (.A(n_1_737_5172), .ZN(n_1_737_5171));
   NAND2_X1 i_1_737_5922 (.A1(n_1_737_5183), .A2(n_1_737_5175), .ZN(n_1_737_5172));
   NOR2_X1 i_1_737_5923 (.A1(n_1_737_5179), .A2(n_1_737_5174), .ZN(n_1_737_5173));
   INV_X1 i_1_737_5924 (.A(n_1_737_5175), .ZN(n_1_737_5174));
   NOR2_X1 i_1_737_5925 (.A1(n_846), .A2(n_849), .ZN(n_1_737_5175));
   NOR2_X1 i_1_737_5926 (.A1(n_1_737_5181), .A2(n_1_737_5177), .ZN(n_1_737_5176));
   INV_X1 i_1_737_5927 (.A(n_1_737_5178), .ZN(n_1_737_5177));
   NOR2_X1 i_1_737_5928 (.A1(n_848), .A2(n_846), .ZN(n_1_737_5178));
   INV_X1 i_1_737_5929 (.A(n_1_737_5180), .ZN(n_1_737_5179));
   NOR2_X1 i_1_737_5930 (.A1(n_848), .A2(n_1_737_5181), .ZN(n_1_737_5180));
   NOR2_X1 i_1_737_5933 (.A1(n_1313), .A2(\out_bs[5] [0]), .ZN(n_1_737_5183));
   NAND3_X1 i_1_737_5934 (.A1(n_1_737_5279), .A2(n_1_737_5233), .A3(n_1_737_5184), 
      .ZN(n_745));
   AOI211_X1 i_1_737_5935 (.A(n_1_737_5363), .B(n_1_737_5185), .C1(n_1_737_5346), 
      .C2(n_1_737_5336), .ZN(n_1_737_5184));
   NAND2_X1 i_1_737_5936 (.A1(n_1_737_5278), .A2(n_1_737_5186), .ZN(n_1_737_5185));
   INV_X1 i_1_737_5937 (.A(n_1_737_5187), .ZN(n_1_737_5186));
   OAI21_X1 i_1_737_5938 (.A(n_1_737_5188), .B1(n_1_737_5202), .B2(n_1_737_5190), 
      .ZN(n_1_737_5187));
   OAI22_X1 i_1_737_5939 (.A1(n_1_737_5223), .A2(n_1_737_5219), .B1(n_1_737_5203), 
      .B2(n_1_737_5189), .ZN(n_1_737_5188));
   INV_X1 i_1_737_5940 (.A(n_1_737_5190), .ZN(n_1_737_5189));
   OAI21_X1 i_1_737_5941 (.A(n_1_737_5191), .B1(\out_as[3] [6]), .B2(
      n_1_737_5192), .ZN(n_1_737_5190));
   OAI21_X1 i_1_737_5942 (.A(\out_bs[3] [6]), .B1(n_1_737_5631), .B2(
      n_1_737_5193), .ZN(n_1_737_5191));
   INV_X1 i_1_737_5943 (.A(n_1_737_5193), .ZN(n_1_737_5192));
   OAI21_X1 i_1_737_5944 (.A(n_1_737_5194), .B1(n_1_737_5637), .B2(
      \out_as[3] [5]), .ZN(n_1_737_5193));
   OAI221_X1 i_1_737_5945 (.A(n_1_737_5195), .B1(\out_bs[3] [4]), .B2(
      n_1_737_5629), .C1(\out_bs[3] [5]), .C2(n_1_737_5630), .ZN(n_1_737_5194));
   OAI221_X1 i_1_737_5946 (.A(n_1_737_5196), .B1(n_1_737_5635), .B2(
      \out_as[3] [3]), .C1(n_1_737_5636), .C2(\out_as[3] [4]), .ZN(n_1_737_5195));
   OAI222_X1 i_1_737_5947 (.A1(\out_bs[3] [3]), .A2(n_1_737_5628), .B1(
      \out_bs[3] [2]), .B2(n_1_737_5627), .C1(n_1_737_5198), .C2(n_1_737_5197), 
      .ZN(n_1_737_5196));
   NOR2_X1 i_1_737_5948 (.A1(n_1_737_5634), .A2(\out_as[3] [2]), .ZN(
      n_1_737_5197));
   OAI21_X1 i_1_737_5949 (.A(n_1_737_5199), .B1(\out_as[3] [1]), .B2(
      n_1_737_5200), .ZN(n_1_737_5198));
   OAI21_X1 i_1_737_5950 (.A(\out_bs[3] [1]), .B1(n_1_737_5626), .B2(
      n_1_737_5201), .ZN(n_1_737_5199));
   INV_X1 i_1_737_5951 (.A(n_1_737_5201), .ZN(n_1_737_5200));
   NAND2_X1 i_1_737_5952 (.A1(n_1_737_5632), .A2(\out_as[3] [0]), .ZN(
      n_1_737_5201));
   INV_X1 i_1_737_5953 (.A(n_1_737_5203), .ZN(n_1_737_5202));
   NOR2_X1 i_1_737_5954 (.A1(\out_as[3] [6]), .A2(n_1_737_5204), .ZN(
      n_1_737_5203));
   OR2_X1 i_1_737_5955 (.A1(\out_as[3] [5]), .A2(n_1_737_5205), .ZN(n_1_737_5204));
   OR2_X1 i_1_737_5956 (.A1(\out_as[3] [4]), .A2(n_1_737_5207), .ZN(n_1_737_5205));
   NAND3_X1 i_1_737_5957 (.A1(n_1_737_5629), .A2(n_1_737_5628), .A3(n_1_737_5627), 
      .ZN(n_1_737_5206));
   OR2_X1 i_1_737_5958 (.A1(\out_as[3] [3]), .A2(n_1_737_5218), .ZN(n_1_737_5207));
   NAND2_X1 i_1_737_5959 (.A1(n_1_737_5628), .A2(n_1_737_5627), .ZN(n_1_737_5208));
   INV_X1 i_1_737_5960 (.A(n_1_737_5210), .ZN(n_1_737_5209));
   NOR2_X1 i_1_737_5961 (.A1(\out_as[3] [6]), .A2(n_1_737_5211), .ZN(
      n_1_737_5210));
   NAND3_X1 i_1_737_5962 (.A1(n_1_737_5630), .A2(n_1_737_5629), .A3(n_1_737_5628), 
      .ZN(n_1_737_5211));
   NAND2_X1 i_1_737_5963 (.A1(n_1_737_5629), .A2(n_1_737_5628), .ZN(n_1_737_5212));
   INV_X1 i_1_737_5964 (.A(n_1_737_5214), .ZN(n_1_737_5213));
   NOR2_X1 i_1_737_5965 (.A1(\out_as[3] [6]), .A2(n_1_737_5217), .ZN(
      n_1_737_5214));
   INV_X1 i_1_737_5966 (.A(n_1_737_5216), .ZN(n_1_737_5215));
   NOR2_X1 i_1_737_5967 (.A1(\out_as[3] [6]), .A2(\out_as[3] [5]), .ZN(
      n_1_737_5216));
   NAND2_X1 i_1_737_5968 (.A1(n_1_737_5630), .A2(n_1_737_5629), .ZN(n_1_737_5217));
   NAND2_X1 i_1_737_5969 (.A1(n_1_737_5627), .A2(n_1_737_5626), .ZN(n_1_737_5218));
   INV_X1 i_1_737_5970 (.A(n_1_737_5220), .ZN(n_1_737_5219));
   NOR2_X1 i_1_737_5971 (.A1(\out_bs[3] [6]), .A2(n_1_737_5228), .ZN(
      n_1_737_5220));
   INV_X1 i_1_737_5972 (.A(n_1_737_5222), .ZN(n_1_737_5221));
   NOR2_X1 i_1_737_5973 (.A1(\out_bs[3] [6]), .A2(\out_bs[3] [5]), .ZN(
      n_1_737_5222));
   NAND2_X1 i_1_737_5974 (.A1(n_1_737_5232), .A2(n_1_737_5225), .ZN(n_1_737_5223));
   INV_X1 i_1_737_5975 (.A(n_1_737_5225), .ZN(n_1_737_5224));
   NOR2_X1 i_1_737_5976 (.A1(\out_bs[3] [3]), .A2(\out_bs[3] [2]), .ZN(
      n_1_737_5225));
   INV_X1 i_1_737_5977 (.A(n_1_737_5227), .ZN(n_1_737_5226));
   NOR2_X1 i_1_737_5978 (.A1(\out_bs[3] [5]), .A2(n_1_737_5230), .ZN(
      n_1_737_5227));
   INV_X1 i_1_737_5979 (.A(n_1_737_5229), .ZN(n_1_737_5228));
   NOR2_X1 i_1_737_5980 (.A1(\out_bs[3] [5]), .A2(\out_bs[3] [4]), .ZN(
      n_1_737_5229));
   INV_X1 i_1_737_5981 (.A(n_1_737_5231), .ZN(n_1_737_5230));
   NOR2_X1 i_1_737_5982 (.A1(\out_bs[3] [4]), .A2(\out_bs[3] [3]), .ZN(
      n_1_737_5231));
   NOR2_X1 i_1_737_5983 (.A1(\out_bs[3] [1]), .A2(\out_bs[3] [0]), .ZN(
      n_1_737_5232));
   OAI22_X1 i_1_737_5984 (.A1(n_1_737_5264), .A2(n_1_737_5234), .B1(n_1_737_5248), 
      .B2(n_1_737_5235), .ZN(n_1_737_5233));
   NOR2_X1 i_1_737_5985 (.A1(n_1_737_5249), .A2(n_1_737_5236), .ZN(n_1_737_5234));
   INV_X1 i_1_737_5986 (.A(n_1_737_5236), .ZN(n_1_737_5235));
   OAI21_X1 i_1_737_5987 (.A(n_1_737_5237), .B1(\out_as[2] [6]), .B2(
      n_1_737_5238), .ZN(n_1_737_5236));
   OAI21_X1 i_1_737_5988 (.A(\out_bs[2] [6]), .B1(n_1_737_5644), .B2(
      n_1_737_5239), .ZN(n_1_737_5237));
   INV_X1 i_1_737_5989 (.A(n_1_737_5239), .ZN(n_1_737_5238));
   OAI21_X1 i_1_737_5990 (.A(n_1_737_5240), .B1(n_1_737_5650), .B2(
      \out_as[2] [5]), .ZN(n_1_737_5239));
   OAI221_X1 i_1_737_5991 (.A(n_1_737_5241), .B1(\out_bs[2] [4]), .B2(
      n_1_737_5642), .C1(\out_bs[2] [5]), .C2(n_1_737_5643), .ZN(n_1_737_5240));
   OAI221_X1 i_1_737_5992 (.A(n_1_737_5242), .B1(n_1_737_5648), .B2(
      \out_as[2] [3]), .C1(n_1_737_5649), .C2(\out_as[2] [4]), .ZN(n_1_737_5241));
   OAI222_X1 i_1_737_5993 (.A1(\out_bs[2] [2]), .A2(n_1_737_5640), .B1(
      \out_bs[2] [3]), .B2(n_1_737_5641), .C1(n_1_737_5244), .C2(n_1_737_5243), 
      .ZN(n_1_737_5242));
   NOR2_X1 i_1_737_5994 (.A1(n_1_737_5647), .A2(\out_as[2] [2]), .ZN(
      n_1_737_5243));
   OAI21_X1 i_1_737_5995 (.A(n_1_737_5245), .B1(\out_as[2] [1]), .B2(
      n_1_737_5246), .ZN(n_1_737_5244));
   OAI21_X1 i_1_737_5996 (.A(\out_bs[2] [1]), .B1(n_1_737_5639), .B2(
      n_1_737_5247), .ZN(n_1_737_5245));
   INV_X1 i_1_737_5997 (.A(n_1_737_5247), .ZN(n_1_737_5246));
   NAND2_X1 i_1_737_5998 (.A1(n_1_737_5645), .A2(\out_as[2] [0]), .ZN(
      n_1_737_5247));
   INV_X1 i_1_737_5999 (.A(n_1_737_5249), .ZN(n_1_737_5248));
   NOR2_X1 i_1_737_6000 (.A1(n_1_737_5254), .A2(n_1_737_5250), .ZN(n_1_737_5249));
   INV_X1 i_1_737_6001 (.A(n_1_737_5251), .ZN(n_1_737_5250));
   NOR2_X1 i_1_737_6002 (.A1(\out_bs[2] [6]), .A2(n_1_737_5259), .ZN(
      n_1_737_5251));
   INV_X1 i_1_737_6003 (.A(n_1_737_5253), .ZN(n_1_737_5252));
   NOR2_X1 i_1_737_6004 (.A1(\out_bs[2] [6]), .A2(\out_bs[2] [5]), .ZN(
      n_1_737_5253));
   NAND2_X1 i_1_737_6005 (.A1(n_1_737_5263), .A2(n_1_737_5257), .ZN(n_1_737_5254));
   NOR2_X1 i_1_737_6006 (.A1(n_1_737_5259), .A2(n_1_737_5256), .ZN(n_1_737_5255));
   INV_X1 i_1_737_6007 (.A(n_1_737_5257), .ZN(n_1_737_5256));
   NOR2_X1 i_1_737_6008 (.A1(\out_bs[2] [3]), .A2(\out_bs[2] [2]), .ZN(
      n_1_737_5257));
   NAND2_X1 i_1_737_6009 (.A1(n_1_737_5650), .A2(n_1_737_5262), .ZN(n_1_737_5258));
   INV_X1 i_1_737_6010 (.A(n_1_737_5260), .ZN(n_1_737_5259));
   NOR2_X1 i_1_737_6011 (.A1(\out_bs[2] [5]), .A2(\out_bs[2] [4]), .ZN(
      n_1_737_5260));
   INV_X1 i_1_737_6012 (.A(n_1_737_5262), .ZN(n_1_737_5261));
   NOR2_X1 i_1_737_6013 (.A1(\out_bs[2] [4]), .A2(\out_bs[2] [3]), .ZN(
      n_1_737_5262));
   NOR2_X1 i_1_737_6014 (.A1(\out_bs[2] [1]), .A2(\out_bs[2] [0]), .ZN(
      n_1_737_5263));
   NOR2_X1 i_1_737_6015 (.A1(\out_as[2] [6]), .A2(n_1_737_5265), .ZN(
      n_1_737_5264));
   OR2_X1 i_1_737_6016 (.A1(\out_as[2] [5]), .A2(n_1_737_5266), .ZN(n_1_737_5265));
   OR2_X1 i_1_737_6017 (.A1(\out_as[2] [4]), .A2(n_1_737_5268), .ZN(n_1_737_5266));
   NAND3_X1 i_1_737_6018 (.A1(n_1_737_5642), .A2(n_1_737_5641), .A3(n_1_737_5640), 
      .ZN(n_1_737_5267));
   OR2_X1 i_1_737_6019 (.A1(\out_as[2] [3]), .A2(n_1_737_5277), .ZN(n_1_737_5268));
   NAND2_X1 i_1_737_6020 (.A1(n_1_737_5641), .A2(n_1_737_5640), .ZN(n_1_737_5269));
   OR2_X1 i_1_737_6021 (.A1(\out_as[2] [6]), .A2(n_1_737_5271), .ZN(n_1_737_5270));
   NAND3_X1 i_1_737_6022 (.A1(n_1_737_5643), .A2(n_1_737_5642), .A3(n_1_737_5641), 
      .ZN(n_1_737_5271));
   NAND2_X1 i_1_737_6023 (.A1(n_1_737_5642), .A2(n_1_737_5641), .ZN(n_1_737_5272));
   NAND2_X1 i_1_737_6024 (.A1(n_1_737_5642), .A2(n_1_737_5275), .ZN(n_1_737_5273));
   INV_X1 i_1_737_6025 (.A(n_1_737_5275), .ZN(n_1_737_5274));
   NOR2_X1 i_1_737_6026 (.A1(\out_as[2] [6]), .A2(\out_as[2] [5]), .ZN(
      n_1_737_5275));
   NAND2_X1 i_1_737_6027 (.A1(n_1_737_5643), .A2(n_1_737_5642), .ZN(n_1_737_5276));
   NAND2_X1 i_1_737_6028 (.A1(n_1_737_5640), .A2(n_1_737_5639), .ZN(n_1_737_5277));
   OAI21_X1 i_1_737_6029 (.A(n_1_737_5324), .B1(n_1_737_5346), .B2(n_1_737_5336), 
      .ZN(n_1_737_5278));
   INV_X1 i_1_737_6030 (.A(n_1_737_5280), .ZN(n_1_737_5279));
   OAI21_X1 i_1_737_6031 (.A(n_1_737_5281), .B1(n_1_737_5307), .B2(n_1_737_5298), 
      .ZN(n_1_737_5280));
   OAI22_X1 i_1_737_6032 (.A1(n_1_737_5287), .A2(n_1_737_5282), .B1(n_1_737_5308), 
      .B2(n_1_737_5297), .ZN(n_1_737_5281));
   INV_X1 i_1_737_6033 (.A(n_1_737_5283), .ZN(n_1_737_5282));
   NOR2_X1 i_1_737_6034 (.A1(\out_bs[1] [6]), .A2(n_1_737_5292), .ZN(
      n_1_737_5283));
   INV_X1 i_1_737_6035 (.A(n_1_737_5285), .ZN(n_1_737_5284));
   NOR2_X1 i_1_737_6036 (.A1(\out_bs[1] [6]), .A2(\out_bs[1] [5]), .ZN(
      n_1_737_5285));
   INV_X1 i_1_737_6037 (.A(n_1_737_5287), .ZN(n_1_737_5286));
   NAND2_X1 i_1_737_6038 (.A1(n_1_737_5296), .A2(n_1_737_5289), .ZN(n_1_737_5287));
   NOR2_X1 i_1_737_6039 (.A1(\out_bs[1] [2]), .A2(n_1_737_5290), .ZN(
      n_1_737_5288));
   NOR2_X1 i_1_737_6040 (.A1(\out_bs[1] [3]), .A2(\out_bs[1] [2]), .ZN(
      n_1_737_5289));
   INV_X1 i_1_737_6041 (.A(n_1_737_5291), .ZN(n_1_737_5290));
   NOR2_X1 i_1_737_6042 (.A1(\out_bs[1] [5]), .A2(n_1_737_5294), .ZN(
      n_1_737_5291));
   INV_X1 i_1_737_6043 (.A(n_1_737_5293), .ZN(n_1_737_5292));
   NOR2_X1 i_1_737_6044 (.A1(\out_bs[1] [5]), .A2(\out_bs[1] [4]), .ZN(
      n_1_737_5293));
   INV_X1 i_1_737_6045 (.A(n_1_737_5295), .ZN(n_1_737_5294));
   NOR2_X1 i_1_737_6046 (.A1(\out_bs[1] [4]), .A2(\out_bs[1] [3]), .ZN(
      n_1_737_5295));
   NOR2_X1 i_1_737_6047 (.A1(\out_bs[1] [1]), .A2(\out_bs[1] [0]), .ZN(
      n_1_737_5296));
   INV_X1 i_1_737_6048 (.A(n_1_737_5298), .ZN(n_1_737_5297));
   OAI21_X1 i_1_737_6049 (.A(n_1_737_5299), .B1(\out_as[1] [6]), .B2(
      n_1_737_5300), .ZN(n_1_737_5298));
   OAI21_X1 i_1_737_6050 (.A(\out_bs[1] [6]), .B1(n_1_737_5658), .B2(
      n_1_737_5301), .ZN(n_1_737_5299));
   INV_X1 i_1_737_6051 (.A(n_1_737_5301), .ZN(n_1_737_5300));
   OAI21_X1 i_1_737_6052 (.A(n_1_737_5302), .B1(n_1_737_5663), .B2(
      \out_as[1] [5]), .ZN(n_1_737_5301));
   OAI221_X1 i_1_737_6053 (.A(n_1_737_5303), .B1(\out_bs[1] [4]), .B2(
      n_1_737_5656), .C1(\out_bs[1] [5]), .C2(n_1_737_5657), .ZN(n_1_737_5302));
   OAI221_X1 i_1_737_6054 (.A(n_1_737_5304), .B1(n_1_737_5661), .B2(
      \out_as[1] [3]), .C1(n_1_737_5662), .C2(\out_as[1] [4]), .ZN(n_1_737_5303));
   OAI221_X1 i_1_737_6055 (.A(n_1_737_5305), .B1(\out_bs[1] [2]), .B2(
      n_1_737_5654), .C1(\out_bs[1] [3]), .C2(n_1_737_5655), .ZN(n_1_737_5304));
   OAI221_X1 i_1_737_6056 (.A(n_1_737_5306), .B1(n_1_737_5659), .B2(
      \out_as[1] [1]), .C1(n_1_737_5660), .C2(\out_as[1] [2]), .ZN(n_1_737_5305));
   OAI22_X1 i_1_737_6057 (.A1(\out_bs[1] [0]), .A2(n_1_737_5652), .B1(
      \out_bs[1] [1]), .B2(n_1_737_5653), .ZN(n_1_737_5306));
   INV_X1 i_1_737_6058 (.A(n_1_737_5308), .ZN(n_1_737_5307));
   NOR2_X1 i_1_737_6059 (.A1(\out_as[1] [6]), .A2(n_1_737_5309), .ZN(
      n_1_737_5308));
   OR2_X1 i_1_737_6060 (.A1(\out_as[1] [5]), .A2(n_1_737_5310), .ZN(n_1_737_5309));
   OR2_X1 i_1_737_6061 (.A1(\out_as[1] [4]), .A2(n_1_737_5312), .ZN(n_1_737_5310));
   NAND3_X1 i_1_737_6062 (.A1(n_1_737_5656), .A2(n_1_737_5655), .A3(n_1_737_5654), 
      .ZN(n_1_737_5311));
   OR2_X1 i_1_737_6063 (.A1(\out_as[1] [3]), .A2(n_1_737_5323), .ZN(n_1_737_5312));
   NAND2_X1 i_1_737_6064 (.A1(n_1_737_5655), .A2(n_1_737_5654), .ZN(n_1_737_5313));
   INV_X1 i_1_737_6065 (.A(n_1_737_5315), .ZN(n_1_737_5314));
   NOR2_X1 i_1_737_6066 (.A1(\out_as[1] [6]), .A2(n_1_737_5316), .ZN(
      n_1_737_5315));
   NAND3_X1 i_1_737_6067 (.A1(n_1_737_5657), .A2(n_1_737_5656), .A3(n_1_737_5655), 
      .ZN(n_1_737_5316));
   NAND2_X1 i_1_737_6068 (.A1(n_1_737_5656), .A2(n_1_737_5655), .ZN(n_1_737_5317));
   INV_X1 i_1_737_6069 (.A(n_1_737_5319), .ZN(n_1_737_5318));
   NOR2_X1 i_1_737_6070 (.A1(\out_as[1] [6]), .A2(n_1_737_5322), .ZN(
      n_1_737_5319));
   INV_X1 i_1_737_6071 (.A(n_1_737_5321), .ZN(n_1_737_5320));
   NOR2_X1 i_1_737_6072 (.A1(\out_as[1] [6]), .A2(\out_as[1] [5]), .ZN(
      n_1_737_5321));
   NAND2_X1 i_1_737_6073 (.A1(n_1_737_5657), .A2(n_1_737_5656), .ZN(n_1_737_5322));
   NAND2_X1 i_1_737_6074 (.A1(n_1_737_5654), .A2(n_1_737_5653), .ZN(n_1_737_5323));
   NAND3_X1 i_1_737_6075 (.A1(n_1_737_5332), .A2(n_1_737_5325), .A3(n_1_737_5671), 
      .ZN(n_1_737_5324));
   INV_X1 i_1_737_6076 (.A(n_1_737_5326), .ZN(n_1_737_5325));
   NAND2_X1 i_1_737_6077 (.A1(n_1_737_5335), .A2(n_1_737_5329), .ZN(n_1_737_5326));
   NOR2_X1 i_1_737_6078 (.A1(n_1_737_5331), .A2(n_1_737_5328), .ZN(n_1_737_5327));
   INV_X1 i_1_737_6079 (.A(n_1_737_5329), .ZN(n_1_737_5328));
   NOR2_X1 i_1_737_6080 (.A1(\out_bs[0] [3]), .A2(\out_bs[0] [2]), .ZN(
      n_1_737_5329));
   NAND2_X1 i_1_737_6081 (.A1(n_1_737_5670), .A2(n_1_737_5334), .ZN(n_1_737_5330));
   INV_X1 i_1_737_6082 (.A(n_1_737_5332), .ZN(n_1_737_5331));
   NOR2_X1 i_1_737_6083 (.A1(\out_bs[0] [5]), .A2(\out_bs[0] [4]), .ZN(
      n_1_737_5332));
   INV_X1 i_1_737_6084 (.A(n_1_737_5334), .ZN(n_1_737_5333));
   NOR2_X1 i_1_737_6085 (.A1(\out_bs[0] [4]), .A2(\out_bs[0] [3]), .ZN(
      n_1_737_5334));
   NOR2_X1 i_1_737_6086 (.A1(\out_bs[0] [1]), .A2(\out_bs[0] [0]), .ZN(
      n_1_737_5335));
   INV_X1 i_1_737_6087 (.A(n_1_737_5337), .ZN(n_1_737_5336));
   OAI21_X1 i_1_737_6089 (.A(\out_bs[0] [6]), .B1(n_1_737_5678), .B2(
      n_1_737_5340), .ZN(n_1_737_5338));
   INV_X1 i_1_737_6090 (.A(n_1_737_5340), .ZN(n_1_737_5339));
   OAI22_X1 i_1_737_6091 (.A1(\out_as[0] [5]), .A2(n_1_737_5670), .B1(
      n_1_737_5342), .B2(n_1_737_5341), .ZN(n_1_737_5340));
   OAI22_X1 i_1_737_6092 (.A1(n_1_737_5676), .A2(\out_bs[0] [4]), .B1(
      n_1_737_5677), .B2(\out_bs[0] [5]), .ZN(n_1_737_5341));
   AOI222_X1 i_1_737_6093 (.A1(n_1_737_5675), .A2(\out_bs[0] [3]), .B1(
      n_1_737_5676), .B2(\out_bs[0] [4]), .C1(n_1_737_5344), .C2(n_1_737_5343), 
      .ZN(n_1_737_5342));
   AOI22_X1 i_1_737_6094 (.A1(\out_as[0] [2]), .A2(n_1_737_5667), .B1(
      \out_as[0] [3]), .B2(n_1_737_5668), .ZN(n_1_737_5343));
   OAI221_X1 i_1_737_6095 (.A(n_1_737_5345), .B1(\out_as[0] [2]), .B2(
      n_1_737_5667), .C1(\out_as[0] [1]), .C2(n_1_737_5666), .ZN(n_1_737_5344));
   OAI22_X1 i_1_737_6096 (.A1(n_1_737_5672), .A2(\out_bs[0] [0]), .B1(
      n_1_737_5673), .B2(\out_bs[0] [1]), .ZN(n_1_737_5345));
   NOR2_X1 i_1_737_6097 (.A1(\out_as[0] [6]), .A2(n_1_737_5347), .ZN(
      n_1_737_5346));
   OR2_X1 i_1_737_6098 (.A1(\out_as[0] [5]), .A2(n_1_737_5348), .ZN(n_1_737_5347));
   OR2_X1 i_1_737_6099 (.A1(\out_as[0] [4]), .A2(n_1_737_5350), .ZN(n_1_737_5348));
   NAND3_X1 i_1_737_6100 (.A1(n_1_737_5676), .A2(n_1_737_5675), .A3(n_1_737_5674), 
      .ZN(n_1_737_5349));
   OR2_X1 i_1_737_6101 (.A1(\out_as[0] [3]), .A2(n_1_737_5361), .ZN(n_1_737_5350));
   NAND2_X1 i_1_737_6102 (.A1(n_1_737_5675), .A2(n_1_737_5674), .ZN(n_1_737_5351));
   INV_X1 i_1_737_6103 (.A(n_1_737_5353), .ZN(n_1_737_5352));
   NOR2_X1 i_1_737_6104 (.A1(\out_as[0] [6]), .A2(n_1_737_5354), .ZN(
      n_1_737_5353));
   NAND3_X1 i_1_737_6105 (.A1(n_1_737_5677), .A2(n_1_737_5676), .A3(n_1_737_5675), 
      .ZN(n_1_737_5354));
   NAND2_X1 i_1_737_6106 (.A1(n_1_737_5676), .A2(n_1_737_5675), .ZN(n_1_737_5355));
   INV_X1 i_1_737_6107 (.A(n_1_737_5357), .ZN(n_1_737_5356));
   NAND2_X1 i_1_737_6108 (.A1(n_1_737_5676), .A2(n_1_737_5359), .ZN(n_1_737_5357));
   INV_X1 i_1_737_6109 (.A(n_1_737_5359), .ZN(n_1_737_5358));
   NOR2_X1 i_1_737_6110 (.A1(\out_as[0] [6]), .A2(\out_as[0] [5]), .ZN(
      n_1_737_5359));
   NAND2_X1 i_1_737_6111 (.A1(n_1_737_5677), .A2(n_1_737_5676), .ZN(n_1_737_5360));
   NAND2_X1 i_1_737_6112 (.A1(n_1_737_5674), .A2(n_1_737_5673), .ZN(n_1_737_5361));
   INV_X1 i_1_737_6113 (.A(n_1_737_5363), .ZN(n_1_737_5362));
   OAI21_X1 i_1_737_6114 (.A(n_1_737_5364), .B1(n_1_737_5375), .B2(n_1_737_5366), 
      .ZN(n_1_737_5363));
   OAI22_X1 i_1_737_6115 (.A1(n_1_737_5394), .A2(n_1_737_5390), .B1(n_1_737_5376), 
      .B2(n_1_737_5365), .ZN(n_1_737_5364));
   INV_X1 i_1_737_6116 (.A(n_1_737_5366), .ZN(n_1_737_5365));
   OAI21_X1 i_1_737_6117 (.A(n_1_737_5367), .B1(\out_as[4] [6]), .B2(
      n_1_737_5368), .ZN(n_1_737_5366));
   OAI21_X1 i_1_737_6118 (.A(\out_bs[4] [6]), .B1(n_1_737_5619), .B2(
      n_1_737_5369), .ZN(n_1_737_5367));
   INV_X1 i_1_737_6119 (.A(n_1_737_5369), .ZN(n_1_737_5368));
   OAI22_X1 i_1_737_6120 (.A1(n_1_737_5624), .A2(\out_as[4] [5]), .B1(
      n_1_737_5371), .B2(n_1_737_5370), .ZN(n_1_737_5369));
   OAI22_X1 i_1_737_6121 (.A1(\out_bs[4] [4]), .A2(n_1_737_5617), .B1(
      \out_bs[4] [5]), .B2(n_1_737_5618), .ZN(n_1_737_5370));
   AOI222_X1 i_1_737_6122 (.A1(\out_bs[4] [3]), .A2(n_1_737_5616), .B1(
      \out_bs[4] [4]), .B2(n_1_737_5617), .C1(n_1_737_5373), .C2(n_1_737_5372), 
      .ZN(n_1_737_5371));
   AOI22_X1 i_1_737_6123 (.A1(n_1_737_5621), .A2(\out_as[4] [2]), .B1(
      n_1_737_5622), .B2(\out_as[4] [3]), .ZN(n_1_737_5372));
   OAI221_X1 i_1_737_6124 (.A(n_1_737_5374), .B1(n_1_737_5621), .B2(
      \out_as[4] [2]), .C1(n_1_737_5620), .C2(\out_as[4] [1]), .ZN(n_1_737_5373));
   OAI22_X1 i_1_737_6125 (.A1(\out_bs[4] [0]), .A2(n_1_737_5613), .B1(
      \out_bs[4] [1]), .B2(n_1_737_5614), .ZN(n_1_737_5374));
   INV_X1 i_1_737_6126 (.A(n_1_737_5376), .ZN(n_1_737_5375));
   NOR2_X1 i_1_737_6127 (.A1(\out_as[4] [6]), .A2(n_1_737_5377), .ZN(
      n_1_737_5376));
   OR2_X1 i_1_737_6128 (.A1(\out_as[4] [5]), .A2(n_1_737_5378), .ZN(n_1_737_5377));
   OR2_X1 i_1_737_6129 (.A1(\out_as[4] [4]), .A2(n_1_737_5380), .ZN(n_1_737_5378));
   NAND3_X1 i_1_737_6130 (.A1(n_1_737_5617), .A2(n_1_737_5616), .A3(n_1_737_5615), 
      .ZN(n_1_737_5379));
   OR2_X1 i_1_737_6131 (.A1(\out_as[4] [3]), .A2(n_1_737_5389), .ZN(n_1_737_5380));
   NAND2_X1 i_1_737_6132 (.A1(n_1_737_5616), .A2(n_1_737_5615), .ZN(n_1_737_5381));
   OR2_X1 i_1_737_6133 (.A1(\out_as[4] [6]), .A2(n_1_737_5383), .ZN(n_1_737_5382));
   NAND3_X1 i_1_737_6134 (.A1(n_1_737_5618), .A2(n_1_737_5617), .A3(n_1_737_5616), 
      .ZN(n_1_737_5383));
   NAND2_X1 i_1_737_6135 (.A1(n_1_737_5617), .A2(n_1_737_5616), .ZN(n_1_737_5384));
   NAND2_X1 i_1_737_6136 (.A1(n_1_737_5617), .A2(n_1_737_5387), .ZN(n_1_737_5385));
   INV_X1 i_1_737_6137 (.A(n_1_737_5387), .ZN(n_1_737_5386));
   NOR2_X1 i_1_737_6138 (.A1(\out_as[4] [6]), .A2(\out_as[4] [5]), .ZN(
      n_1_737_5387));
   NAND2_X1 i_1_737_6139 (.A1(n_1_737_5618), .A2(n_1_737_5617), .ZN(n_1_737_5388));
   NAND2_X1 i_1_737_6140 (.A1(n_1_737_5615), .A2(n_1_737_5614), .ZN(n_1_737_5389));
   INV_X1 i_1_737_6141 (.A(n_1_737_5391), .ZN(n_1_737_5390));
   NOR2_X1 i_1_737_6142 (.A1(\out_bs[4] [6]), .A2(n_1_737_5400), .ZN(
      n_1_737_5391));
   INV_X1 i_1_737_6143 (.A(n_1_737_5393), .ZN(n_1_737_5392));
   NOR2_X1 i_1_737_6144 (.A1(\out_bs[4] [6]), .A2(\out_bs[4] [5]), .ZN(
      n_1_737_5393));
   INV_X1 i_1_737_6145 (.A(n_1_737_5395), .ZN(n_1_737_5394));
   NOR2_X1 i_1_737_6146 (.A1(n_1_737_5404), .A2(n_1_737_5397), .ZN(n_1_737_5395));
   NOR2_X1 i_1_737_6147 (.A1(n_1_737_5400), .A2(n_1_737_5397), .ZN(n_1_737_5396));
   INV_X1 i_1_737_6148 (.A(n_1_737_5398), .ZN(n_1_737_5397));
   NOR2_X1 i_1_737_6149 (.A1(\out_bs[4] [3]), .A2(\out_bs[4] [2]), .ZN(
      n_1_737_5398));
   NAND2_X1 i_1_737_6150 (.A1(n_1_737_5624), .A2(n_1_737_5403), .ZN(n_1_737_5399));
   INV_X1 i_1_737_6151 (.A(n_1_737_5401), .ZN(n_1_737_5400));
   NOR2_X1 i_1_737_6152 (.A1(\out_bs[4] [5]), .A2(\out_bs[4] [4]), .ZN(
      n_1_737_5401));
   INV_X1 i_1_737_6153 (.A(n_1_737_5403), .ZN(n_1_737_5402));
   NOR2_X1 i_1_737_6154 (.A1(\out_bs[4] [4]), .A2(\out_bs[4] [3]), .ZN(
      n_1_737_5403));
   INV_X1 i_1_737_6155 (.A(n_1_737_5405), .ZN(n_1_737_5404));
   NOR2_X1 i_1_737_6156 (.A1(\out_bs[4] [1]), .A2(\out_bs[4] [0]), .ZN(
      n_1_737_5405));
   INV_X1 i_1_737_6157 (.A(n_1_737_954), .ZN(n_1_737_5406));
   INV_X1 i_1_737_6158 (.A(n_1_737_953), .ZN(n_1_737_5407));
   INV_X1 i_1_737_6159 (.A(n_1_737_951), .ZN(n_746));
   INV_X1 i_1_737_6160 (.A(n_1_737_949), .ZN(n_1_737_5408));
   INV_X1 i_1_737_6161 (.A(n_1_737_947), .ZN(n_1_737_5409));
   INV_X1 i_1_737_6162 (.A(n_1_737_946), .ZN(n_1_737_5410));
   INV_X1 i_1_737_6163 (.A(n_1_737_945), .ZN(n_1_737_5411));
   INV_X1 i_1_737_6164 (.A(n_1_737_942), .ZN(n_1_737_5412));
   INV_X1 i_1_737_6165 (.A(n_1_737_939), .ZN(n_1_737_5413));
   INV_X1 i_1_737_6166 (.A(n_1_737_937), .ZN(n_747));
   INV_X1 i_1_737_6167 (.A(n_1_737_935), .ZN(n_1_737_5414));
   INV_X1 i_1_737_6168 (.A(n_1_737_934), .ZN(n_1_737_5415));
   INV_X1 i_1_737_6169 (.A(n_1_737_933), .ZN(n_1_737_5416));
   INV_X1 i_1_737_6170 (.A(n_1_737_932), .ZN(n_1_737_5417));
   INV_X1 i_1_737_6171 (.A(n_1_737_931), .ZN(n_1_737_5418));
   INV_X1 i_1_737_6172 (.A(n_1_737_930), .ZN(n_748));
   INV_X1 i_1_737_6173 (.A(n_1_737_928), .ZN(n_1_737_5419));
   INV_X1 i_1_737_6174 (.A(n_1_737_927), .ZN(n_1_737_5420));
   INV_X1 i_1_737_6175 (.A(n_1_737_925), .ZN(n_1_737_5421));
   INV_X1 i_1_737_6176 (.A(n_1_737_921), .ZN(n_1_737_5422));
   INV_X1 i_1_737_6177 (.A(n_1_737_920), .ZN(n_1_737_5423));
   INV_X1 i_1_737_6178 (.A(n_1_737_919), .ZN(n_1_737_5424));
   INV_X1 i_1_737_6179 (.A(n_1_737_918), .ZN(n_1_737_5425));
   INV_X1 i_1_737_6180 (.A(n_1_737_915), .ZN(n_1_737_5426));
   INV_X1 i_1_737_6181 (.A(n_1_737_914), .ZN(n_1_737_5427));
   INV_X1 i_1_737_6182 (.A(n_1_737_909), .ZN(n_749));
   INV_X1 i_1_737_6183 (.A(n_1_737_907), .ZN(n_1_737_5428));
   INV_X1 i_1_737_6184 (.A(n_1_737_906), .ZN(n_1_737_5429));
   INV_X1 i_1_737_6185 (.A(n_1_737_905), .ZN(n_1_737_5430));
   INV_X1 i_1_737_6186 (.A(n_1_737_900), .ZN(n_1_737_5431));
   INV_X1 i_1_737_6187 (.A(n_1_737_899), .ZN(n_1_737_5432));
   INV_X1 i_1_737_6188 (.A(n_1_737_897), .ZN(n_1_737_5433));
   INV_X1 i_1_737_6189 (.A(n_1_737_893), .ZN(n_1_737_5434));
   INV_X1 i_1_737_6190 (.A(n_1_737_892), .ZN(n_1_737_5435));
   INV_X1 i_1_737_6191 (.A(n_1_737_891), .ZN(n_1_737_5436));
   INV_X1 i_1_737_6192 (.A(n_1_737_890), .ZN(n_1_737_5437));
   INV_X1 i_1_737_6193 (.A(n_1_737_889), .ZN(n_1_737_5438));
   INV_X1 i_1_737_6194 (.A(n_1_737_886), .ZN(n_1_737_5439));
   INV_X1 i_1_737_6195 (.A(n_1_737_885), .ZN(n_1_737_5440));
   INV_X1 i_1_737_6196 (.A(n_1_737_884), .ZN(n_1_737_5441));
   INV_X1 i_1_737_6197 (.A(n_1_737_883), .ZN(n_1_737_5442));
   INV_X1 i_1_737_6198 (.A(n_1_737_879), .ZN(n_1_737_5443));
   INV_X1 i_1_737_6199 (.A(n_1_737_878), .ZN(n_1_737_5444));
   INV_X1 i_1_737_6200 (.A(n_1_737_877), .ZN(n_1_737_5445));
   INV_X1 i_1_737_6201 (.A(n_1_737_876), .ZN(n_1_737_5446));
   INV_X1 i_1_737_6202 (.A(n_1_737_872), .ZN(n_1_737_5447));
   INV_X1 i_1_737_6203 (.A(n_1_737_871), .ZN(n_1_737_5448));
   INV_X1 i_1_737_6204 (.A(n_1_737_870), .ZN(n_1_737_5449));
   INV_X1 i_1_737_6205 (.A(n_1_737_869), .ZN(n_1_737_5450));
   INV_X1 i_1_737_6206 (.A(n_1_737_865), .ZN(n_1_737_5451));
   INV_X1 i_1_737_6207 (.A(n_1_737_864), .ZN(n_1_737_5452));
   INV_X1 i_1_737_6208 (.A(n_1_737_863), .ZN(n_1_737_5453));
   INV_X1 i_1_737_6209 (.A(n_1_737_862), .ZN(n_1_737_5454));
   INV_X1 i_1_737_6210 (.A(n_1_737_853), .ZN(n_750));
   INV_X1 i_1_737_6211 (.A(n_1_737_851), .ZN(n_1_737_5455));
   INV_X1 i_1_737_6212 (.A(n_1_737_850), .ZN(n_1_737_5456));
   INV_X1 i_1_737_6213 (.A(n_1_737_849), .ZN(n_1_737_5457));
   INV_X1 i_1_737_6214 (.A(n_1_737_846), .ZN(n_751));
   INV_X1 i_1_737_6215 (.A(n_1_737_844), .ZN(n_1_737_5458));
   INV_X1 i_1_737_6216 (.A(n_1_737_843), .ZN(n_1_737_5459));
   INV_X1 i_1_737_6217 (.A(n_1_737_842), .ZN(n_1_737_5460));
   INV_X1 i_1_737_6218 (.A(n_1_737_839), .ZN(n_752));
   INV_X1 i_1_737_6219 (.A(n_1_737_834), .ZN(n_1_737_5461));
   INV_X1 i_1_737_6220 (.A(n_1_737_829), .ZN(n_1_737_5462));
   INV_X1 i_1_737_6221 (.A(n_1_737_827), .ZN(n_1_737_5463));
   INV_X1 i_1_737_6222 (.A(n_1_737_825), .ZN(n_753));
   INV_X1 i_1_737_6223 (.A(n_1_737_823), .ZN(n_1_737_5464));
   INV_X1 i_1_737_6224 (.A(n_1_737_821), .ZN(n_1_737_5465));
   INV_X1 i_1_737_6225 (.A(n_1_737_820), .ZN(n_1_737_5466));
   INV_X1 i_1_737_6226 (.A(n_1_737_819), .ZN(n_1_737_5467));
   INV_X1 i_1_737_6227 (.A(n_1_737_816), .ZN(n_1_737_5468));
   INV_X1 i_1_737_6228 (.A(n_1_737_815), .ZN(n_1_737_5469));
   INV_X1 i_1_737_6229 (.A(n_1_737_814), .ZN(n_1_737_5470));
   INV_X1 i_1_737_6230 (.A(n_1_737_809), .ZN(n_1_737_5471));
   INV_X1 i_1_737_6231 (.A(n_1_737_808), .ZN(n_1_737_5472));
   INV_X1 i_1_737_6232 (.A(n_1_737_807), .ZN(n_1_737_5473));
   INV_X1 i_1_737_6233 (.A(n_1_737_804), .ZN(n_754));
   INV_X1 i_1_737_6234 (.A(n_1_737_803), .ZN(n_1_737_5474));
   INV_X1 i_1_737_6235 (.A(n_1_737_795), .ZN(n_1_737_5475));
   INV_X1 i_1_737_6236 (.A(n_1_737_791), .ZN(n_1_737_5476));
   INV_X1 i_1_737_6237 (.A(n_1_737_788), .ZN(n_1_737_5477));
   INV_X1 i_1_737_6238 (.A(n_1_737_785), .ZN(n_1_737_5478));
   INV_X1 i_1_737_6239 (.A(n_1_737_781), .ZN(n_1_737_5479));
   INV_X1 i_1_737_6240 (.A(n_1_737_780), .ZN(n_1_737_5480));
   INV_X1 i_1_737_6241 (.A(n_1_737_779), .ZN(n_1_737_5481));
   INV_X1 i_1_737_6242 (.A(n_1_737_778), .ZN(n_1_737_5482));
   INV_X1 i_1_737_6243 (.A(n_1_737_773), .ZN(n_1_737_5483));
   INV_X1 i_1_737_6244 (.A(n_1_737_771), .ZN(n_1_737_5484));
   INV_X1 i_1_737_6245 (.A(n_1_737_770), .ZN(n_1_737_5485));
   INV_X1 i_1_737_6246 (.A(n_1_737_767), .ZN(n_1_737_5486));
   INV_X1 i_1_737_6247 (.A(n_1_737_764), .ZN(n_1_737_5487));
   INV_X1 i_1_737_6248 (.A(n_1_737_762), .ZN(n_755));
   INV_X1 i_1_737_6249 (.A(n_1_737_759), .ZN(n_1_737_5488));
   INV_X1 i_1_737_6250 (.A(n_1_737_757), .ZN(n_1_737_5489));
   INV_X1 i_1_737_6251 (.A(n_1_737_753), .ZN(n_1_737_5490));
   INV_X1 i_1_737_6252 (.A(n_1_737_752), .ZN(n_1_737_5491));
   INV_X1 i_1_737_6253 (.A(n_1_737_751), .ZN(n_1_737_5492));
   INV_X1 i_1_737_6254 (.A(n_1_737_750), .ZN(n_1_737_5493));
   INV_X1 i_1_737_6255 (.A(n_1_737_748), .ZN(n_756));
   INV_X1 i_1_737_6256 (.A(n_1_737_747), .ZN(n_1_737_5494));
   INV_X1 i_1_737_6257 (.A(n_1_737_745), .ZN(n_1_737_5495));
   INV_X1 i_1_737_6258 (.A(n_1_737_738), .ZN(n_1_737_5496));
   INV_X1 i_1_737_6259 (.A(n_1_737_736), .ZN(n_1_737_5497));
   INV_X1 i_1_737_6260 (.A(n_1_737_732), .ZN(n_1_737_5498));
   INV_X1 i_1_737_6261 (.A(n_1_737_731), .ZN(n_1_737_5499));
   INV_X1 i_1_737_6262 (.A(n_1_737_729), .ZN(n_1_737_5500));
   INV_X1 i_1_737_6263 (.A(n_1_737_723), .ZN(n_1_737_5501));
   INV_X1 i_1_737_6264 (.A(n_1_737_722), .ZN(n_1_737_5502));
   INV_X1 i_1_737_6265 (.A(n_1_737_717), .ZN(n_1_737_5503));
   INV_X1 i_1_737_6266 (.A(n_1_737_716), .ZN(n_1_737_5504));
   INV_X1 i_1_737_6267 (.A(n_1_737_715), .ZN(n_1_737_5505));
   INV_X1 i_1_737_6268 (.A(n_1_737_713), .ZN(n_757));
   INV_X1 i_1_737_6269 (.A(n_1_737_703), .ZN(n_1_737_5506));
   INV_X1 i_1_737_6270 (.A(n_1_737_701), .ZN(n_1_737_5507));
   INV_X1 i_1_737_6271 (.A(n_1_737_699), .ZN(n_758));
   INV_X1 i_1_737_6272 (.A(n_1_737_697), .ZN(n_1_737_5508));
   INV_X1 i_1_737_6273 (.A(n_1_737_696), .ZN(n_1_737_5509));
   INV_X1 i_1_737_6274 (.A(n_1_737_695), .ZN(n_1_737_5510));
   INV_X1 i_1_737_6275 (.A(n_1_737_690), .ZN(n_1_737_5511));
   INV_X1 i_1_737_6276 (.A(n_1_737_688), .ZN(n_1_737_5512));
   INV_X1 i_1_737_6277 (.A(n_1_737_686), .ZN(n_1_737_5513));
   INV_X1 i_1_737_6278 (.A(n_1_737_685), .ZN(n_759));
   INV_X1 i_1_737_6279 (.A(n_1_737_683), .ZN(n_1_737_5514));
   INV_X1 i_1_737_6280 (.A(n_1_737_682), .ZN(n_1_737_5515));
   INV_X1 i_1_737_6281 (.A(n_1_737_681), .ZN(n_1_737_5516));
   INV_X1 i_1_737_6282 (.A(n_1_737_680), .ZN(n_1_737_5517));
   INV_X1 i_1_737_6283 (.A(n_1_737_678), .ZN(n_760));
   INV_X1 i_1_737_6284 (.A(n_1_737_671), .ZN(n_761));
   INV_X1 i_1_737_6285 (.A(n_1_737_669), .ZN(n_1_737_5518));
   INV_X1 i_1_737_6286 (.A(n_1_737_668), .ZN(n_1_737_5519));
   INV_X1 i_1_737_6287 (.A(n_1_737_667), .ZN(n_1_737_5520));
   INV_X1 i_1_737_6288 (.A(n_1_737_666), .ZN(n_1_737_5521));
   INV_X1 i_1_737_6289 (.A(n_1_737_662), .ZN(n_1_737_5522));
   INV_X1 i_1_737_6290 (.A(n_1_737_661), .ZN(n_1_737_5523));
   INV_X1 i_1_737_6291 (.A(n_1_737_660), .ZN(n_1_737_5524));
   INV_X1 i_1_737_6292 (.A(n_1_737_659), .ZN(n_1_737_5525));
   INV_X1 i_1_737_6293 (.A(n_1_737_657), .ZN(n_762));
   INV_X1 i_1_737_6294 (.A(n_1_737_655), .ZN(n_1_737_5526));
   INV_X1 i_1_737_6295 (.A(n_1_737_654), .ZN(n_1_737_5527));
   INV_X1 i_1_737_6296 (.A(n_1_737_652), .ZN(n_1_737_5528));
   INV_X1 i_1_737_6297 (.A(n_1_737_646), .ZN(n_1_737_5529));
   INV_X1 i_1_737_6298 (.A(n_1_737_645), .ZN(n_1_737_5530));
   INV_X1 i_1_737_6299 (.A(n_1_737_643), .ZN(n_763));
   INV_X1 i_1_737_6300 (.A(n_1_737_641), .ZN(n_1_737_5531));
   INV_X1 i_1_737_6301 (.A(n_1_737_640), .ZN(n_1_737_5532));
   INV_X1 i_1_737_6302 (.A(n_1_737_638), .ZN(n_1_737_5533));
   INV_X1 i_1_737_6303 (.A(n_1_737_634), .ZN(n_1_737_5534));
   INV_X1 i_1_737_6304 (.A(n_1_737_631), .ZN(n_1_737_5535));
   INV_X1 i_1_737_6305 (.A(n_1_737_629), .ZN(n_764));
   INV_X1 i_1_737_6306 (.A(n_1_737_627), .ZN(n_1_737_5536));
   INV_X1 i_1_737_6307 (.A(n_1_737_626), .ZN(n_1_737_5537));
   INV_X1 i_1_737_6308 (.A(n_1_737_625), .ZN(n_1_737_5538));
   INV_X1 i_1_737_6309 (.A(n_1_737_624), .ZN(n_1_737_5539));
   INV_X1 i_1_737_6310 (.A(n_1_737_622), .ZN(n_765));
   INV_X1 i_1_737_6311 (.A(n_1_737_620), .ZN(n_1_737_5540));
   INV_X1 i_1_737_6312 (.A(n_1_737_619), .ZN(n_1_737_5541));
   INV_X1 i_1_737_6313 (.A(n_1_737_618), .ZN(n_1_737_5542));
   INV_X1 i_1_737_6314 (.A(n_1_737_617), .ZN(n_1_737_5543));
   INV_X1 i_1_737_6315 (.A(n_1_737_615), .ZN(n_766));
   INV_X1 i_1_737_6316 (.A(n_1_737_613), .ZN(n_1_737_5544));
   INV_X1 i_1_737_6317 (.A(n_1_737_612), .ZN(n_1_737_5545));
   INV_X1 i_1_737_6318 (.A(n_1_737_610), .ZN(n_1_737_5546));
   INV_X1 i_1_737_6319 (.A(n_1_737_606), .ZN(n_1_737_5547));
   INV_X1 i_1_737_6320 (.A(n_1_737_605), .ZN(n_1_737_5548));
   INV_X1 i_1_737_6321 (.A(n_1_737_604), .ZN(n_1_737_5549));
   INV_X1 i_1_737_6322 (.A(n_1_737_603), .ZN(n_1_737_5550));
   INV_X1 i_1_737_6323 (.A(n_1_737_598), .ZN(n_1_737_5551));
   INV_X1 i_1_737_6324 (.A(n_1_737_592), .ZN(n_1_737_5552));
   INV_X1 i_1_737_6325 (.A(n_1_737_591), .ZN(n_1_737_5553));
   INV_X1 i_1_737_6326 (.A(n_1_737_590), .ZN(n_1_737_5554));
   INV_X1 i_1_737_6327 (.A(n_1_737_587), .ZN(n_767));
   INV_X1 i_1_737_6328 (.A(n_1_737_584), .ZN(n_1_737_5555));
   INV_X1 i_1_737_6329 (.A(n_1_737_583), .ZN(n_1_737_5556));
   INV_X1 i_1_737_6330 (.A(n_1_737_582), .ZN(n_1_737_5557));
   INV_X1 i_1_737_6331 (.A(n_1_737_577), .ZN(n_1_737_5558));
   INV_X1 i_1_737_6332 (.A(n_1_737_575), .ZN(n_1_737_5559));
   INV_X1 i_1_737_6333 (.A(n_1_737_571), .ZN(n_1_737_5560));
   INV_X1 i_1_737_6334 (.A(n_1_737_570), .ZN(n_1_737_5561));
   INV_X1 i_1_737_6335 (.A(n_1_737_568), .ZN(n_1_737_5562));
   INV_X1 i_1_737_6336 (.A(n_1_737_564), .ZN(n_1_737_5563));
   INV_X1 i_1_737_6337 (.A(n_1_737_563), .ZN(n_1_737_5564));
   INV_X1 i_1_737_6338 (.A(n_1_737_557), .ZN(n_1_737_5565));
   INV_X1 i_1_737_6339 (.A(n_1_737_556), .ZN(n_1_737_5566));
   INV_X1 i_1_737_6340 (.A(n_1_737_555), .ZN(n_1_737_5567));
   INV_X1 i_1_737_6341 (.A(n_1_737_554), .ZN(n_1_737_5568));
   INV_X1 i_1_737_6342 (.A(n_1_737_552), .ZN(n_768));
   INV_X1 i_1_737_6343 (.A(n_1_737_550), .ZN(n_1_737_5569));
   INV_X1 i_1_737_6344 (.A(n_1_737_548), .ZN(n_1_737_5570));
   INV_X1 i_1_737_6345 (.A(n_1_737_547), .ZN(n_1_737_5571));
   INV_X1 i_1_737_6346 (.A(n_1_737_546), .ZN(n_1_737_5572));
   INV_X1 i_1_737_6347 (.A(n_1_737_545), .ZN(n_769));
   INV_X1 i_1_737_6348 (.A(n_1_737_542), .ZN(n_1_737_5573));
   INV_X1 i_1_737_6349 (.A(n_1_737_541), .ZN(n_1_737_5574));
   INV_X1 i_1_737_6350 (.A(n_1_737_540), .ZN(n_1_737_5575));
   INV_X1 i_1_737_6351 (.A(n_1_737_536), .ZN(n_1_737_5576));
   INV_X1 i_1_737_6352 (.A(n_1_737_535), .ZN(n_1_737_5577));
   INV_X1 i_1_737_6353 (.A(n_1_737_534), .ZN(n_1_737_5578));
   INV_X1 i_1_737_6354 (.A(n_1_737_532), .ZN(n_1_737_5579));
   INV_X1 i_1_737_6355 (.A(n_1_737_531), .ZN(n_770));
   INV_X1 i_1_737_6356 (.A(n_1_737_529), .ZN(n_1_737_5580));
   INV_X1 i_1_737_6357 (.A(n_1_737_528), .ZN(n_1_737_5581));
   INV_X1 i_1_737_6358 (.A(n_1_737_526), .ZN(n_1_737_5582));
   INV_X1 i_1_737_6359 (.A(n_1_737_522), .ZN(n_1_737_5583));
   INV_X1 i_1_737_6360 (.A(n_1_737_521), .ZN(n_1_737_5584));
   INV_X1 i_1_737_6361 (.A(n_1_737_520), .ZN(n_1_737_5585));
   INV_X1 i_1_737_6362 (.A(n_1_737_519), .ZN(n_1_737_5586));
   INV_X1 i_1_737_6363 (.A(n_1_737_192), .ZN(n_1_737_5587));
   INV_X1 i_1_737_6364 (.A(n_1_737_190), .ZN(n_1_737_5588));
   INV_X1 i_1_737_6365 (.A(n_1_737_183), .ZN(n_1_737_5589));
   INV_X1 i_1_737_6366 (.A(n_1_737_155), .ZN(n_1_737_5590));
   INV_X1 i_1_737_6367 (.A(n_1_737_143), .ZN(n_1_737_5591));
   INV_X1 i_1_737_6368 (.A(n_1_737_141), .ZN(n_1_737_5592));
   INV_X1 i_1_737_6369 (.A(n_1_737_134), .ZN(n_1_737_5593));
   INV_X1 i_1_737_6370 (.A(n_1_737_118), .ZN(n_771));
   INV_X1 i_1_737_6371 (.A(n_1_737_112), .ZN(n_772));
   INV_X1 i_1_737_6372 (.A(n_1_737_107), .ZN(n_773));
   INV_X1 i_1_737_6373 (.A(n_1_737_102), .ZN(n_774));
   INV_X1 i_1_737_6374 (.A(n_1_737_98), .ZN(n_775));
   INV_X1 i_1_737_6375 (.A(n_1_737_94), .ZN(n_776));
   INV_X1 i_1_737_6376 (.A(n_1_737_90), .ZN(n_777));
   INV_X1 i_1_737_6377 (.A(n_1_737_86), .ZN(n_778));
   INV_X1 i_1_737_6378 (.A(n_1_737_83), .ZN(n_779));
   INV_X1 i_1_737_6380 (.A(n_1_737_77), .ZN(n_780));
   INV_X1 i_1_737_6381 (.A(n_1_737_74), .ZN(n_781));
   INV_X1 i_1_737_6382 (.A(n_1_737_71), .ZN(n_782));
   INV_X1 i_1_737_6383 (.A(n_1_737_68), .ZN(n_783));
   INV_X1 i_1_737_6384 (.A(n_1_737_65), .ZN(n_784));
   INV_X1 i_1_737_6385 (.A(n_1_737_62), .ZN(n_785));
   INV_X1 i_1_737_6386 (.A(n_1_737_60), .ZN(n_786));
   INV_X1 i_1_737_6387 (.A(n_1_737_58), .ZN(n_787));
   INV_X1 i_1_737_6388 (.A(n_1_737_56), .ZN(n_788));
   INV_X1 i_1_737_6389 (.A(n_1_737_54), .ZN(n_789));
   INV_X1 i_1_737_6390 (.A(n_1_737_52), .ZN(n_790));
   INV_X1 i_1_737_6391 (.A(n_1_737_50), .ZN(n_791));
   INV_X1 i_1_737_6392 (.A(n_1_737_48), .ZN(n_792));
   INV_X1 i_1_737_6393 (.A(n_1_737_46), .ZN(n_793));
   INV_X1 i_1_737_6395 (.A(n_1_737_42), .ZN(n_794));
   INV_X1 i_1_737_6396 (.A(n_1_737_40), .ZN(n_795));
   INV_X1 i_1_737_6397 (.A(n_1_737_38), .ZN(n_796));
   INV_X1 i_1_737_6398 (.A(n_1_737_36), .ZN(n_797));
   INV_X1 i_1_737_6399 (.A(n_1_737_34), .ZN(n_798));
   INV_X1 i_1_737_6400 (.A(n_1_737_32), .ZN(n_799));
   INV_X1 i_1_737_6401 (.A(n_1_737_30), .ZN(n_800));
   INV_X1 i_1_737_6402 (.A(n_1_737_29), .ZN(n_801));
   INV_X1 i_1_737_6403 (.A(n_1_737_28), .ZN(n_802));
   INV_X1 i_1_737_6404 (.A(n_1_737_27), .ZN(n_803));
   INV_X1 i_1_737_6405 (.A(n_1_737_26), .ZN(n_804));
   INV_X1 i_1_737_6406 (.A(n_1_737_25), .ZN(n_805));
   INV_X1 i_1_737_6407 (.A(n_1_737_24), .ZN(n_806));
   INV_X1 i_1_737_6408 (.A(n_1_737_23), .ZN(n_807));
   INV_X1 i_1_737_6409 (.A(n_1_737_22), .ZN(n_808));
   INV_X1 i_1_737_6410 (.A(n_1_737_21), .ZN(n_809));
   INV_X1 i_1_737_6411 (.A(n_1_737_20), .ZN(n_810));
   INV_X1 i_1_737_6412 (.A(n_1_737_19), .ZN(n_811));
   INV_X1 i_1_737_6413 (.A(n_1_737_18), .ZN(n_812));
   INV_X1 i_1_737_6414 (.A(n_1_737_17), .ZN(n_813));
   INV_X1 i_1_737_6415 (.A(n_1_737_16), .ZN(n_814));
   INV_X1 i_1_737_6416 (.A(n_1_737_15), .ZN(n_815));
   INV_X1 i_1_737_6417 (.A(n_1_737_14), .ZN(n_816));
   INV_X1 i_1_737_6418 (.A(n_1_737_13), .ZN(n_817));
   INV_X1 i_1_737_6419 (.A(n_1_737_12), .ZN(n_818));
   INV_X1 i_1_737_6420 (.A(n_1_737_11), .ZN(n_819));
   INV_X1 i_1_737_6421 (.A(n_1_737_10), .ZN(n_820));
   INV_X1 i_1_737_6422 (.A(n_1_737_9), .ZN(n_821));
   INV_X1 i_1_737_6423 (.A(n_1_737_8), .ZN(n_822));
   INV_X1 i_1_737_6424 (.A(n_1_737_7), .ZN(n_823));
   INV_X1 i_1_737_6425 (.A(n_1_737_6), .ZN(n_824));
   INV_X1 i_1_737_6426 (.A(n_1_737_5), .ZN(n_825));
   INV_X1 i_1_737_6427 (.A(n_1_737_4), .ZN(n_826));
   INV_X1 i_1_737_6428 (.A(n_1_737_3), .ZN(n_827));
   INV_X1 i_1_737_6429 (.A(n_1_737_2), .ZN(n_828));
   INV_X1 i_1_737_6430 (.A(n_1_737_1), .ZN(n_829));
   INV_X1 i_1_737_6431 (.A(n_1_737_0), .ZN(n_830));
   INV_X1 i_1_737_6432 (.A(n_952), .ZN(n_1_737_5594));
   INV_X1 i_1_737_6433 (.A(in_data[4]), .ZN(n_1_737_5595));
   INV_X1 i_1_737_6435 (.A(in_data[12]), .ZN(n_1_737_5597));
   INV_X1 i_1_737_6436 (.A(in_data[16]), .ZN(n_1_737_5598));
   INV_X1 i_1_737_6437 (.A(in_data[20]), .ZN(n_1_737_5599));
   INV_X1 i_1_737_6438 (.A(in_data[24]), .ZN(n_1_737_5600));
   INV_X1 i_1_737_6439 (.A(in_data[28]), .ZN(n_1_737_5601));
   INV_X1 i_1_737_6441 (.A(n_851), .ZN(n_1_737_5603));
   INV_X1 i_1_737_6442 (.A(n_847), .ZN(n_1_737_5604));
   INV_X1 i_1_737_6443 (.A(\out_bs[6] [4]), .ZN(n_1_737_5605));
   INV_X1 i_1_737_6444 (.A(\out_bs[6] [5]), .ZN(n_1_737_5606));
   INV_X1 i_1_737_6445 (.A(\out_bs[6] [6]), .ZN(n_1_737_5607));
   INV_X1 i_1_737_6446 (.A(\out_as[7] [6]), .ZN(n_831));
   INV_X1 i_1_737_6447 (.A(n_849), .ZN(n_1_737_5608));
   INV_X1 i_1_737_6448 (.A(n_846), .ZN(n_1_737_5609));
   INV_X1 i_1_737_6449 (.A(n_848), .ZN(n_1_737_5610));
   INV_X1 i_1_737_6450 (.A(n_845), .ZN(n_1_737_5611));
   INV_X1 i_1_737_6451 (.A(n_844), .ZN(n_1_737_5612));
   INV_X1 i_1_737_6452 (.A(\out_as[4] [0]), .ZN(n_1_737_5613));
   INV_X1 i_1_737_6453 (.A(\out_as[4] [1]), .ZN(n_1_737_5614));
   INV_X1 i_1_737_6454 (.A(\out_as[4] [2]), .ZN(n_1_737_5615));
   INV_X1 i_1_737_6455 (.A(\out_as[4] [3]), .ZN(n_1_737_5616));
   INV_X1 i_1_737_6456 (.A(\out_as[4] [4]), .ZN(n_1_737_5617));
   INV_X1 i_1_737_6457 (.A(\out_as[4] [5]), .ZN(n_1_737_5618));
   INV_X1 i_1_737_6458 (.A(\out_as[4] [6]), .ZN(n_1_737_5619));
   INV_X1 i_1_737_6459 (.A(\out_bs[4] [1]), .ZN(n_1_737_5620));
   INV_X1 i_1_737_6460 (.A(\out_bs[4] [2]), .ZN(n_1_737_5621));
   INV_X1 i_1_737_6461 (.A(\out_bs[4] [3]), .ZN(n_1_737_5622));
   INV_X1 i_1_737_6462 (.A(\out_bs[4] [4]), .ZN(n_1_737_5623));
   INV_X1 i_1_737_6463 (.A(\out_bs[4] [5]), .ZN(n_1_737_5624));
   INV_X1 i_1_737_6464 (.A(\out_bs[4] [6]), .ZN(n_1_737_5625));
   INV_X1 i_1_737_6465 (.A(\out_as[3] [1]), .ZN(n_1_737_5626));
   INV_X1 i_1_737_6466 (.A(\out_as[3] [2]), .ZN(n_1_737_5627));
   INV_X1 i_1_737_6467 (.A(\out_as[3] [3]), .ZN(n_1_737_5628));
   INV_X1 i_1_737_6468 (.A(\out_as[3] [4]), .ZN(n_1_737_5629));
   INV_X1 i_1_737_6469 (.A(\out_as[3] [5]), .ZN(n_1_737_5630));
   INV_X1 i_1_737_6470 (.A(\out_as[3] [6]), .ZN(n_1_737_5631));
   INV_X1 i_1_737_6471 (.A(\out_bs[3] [0]), .ZN(n_1_737_5632));
   INV_X1 i_1_737_6472 (.A(\out_bs[3] [1]), .ZN(n_1_737_5633));
   INV_X1 i_1_737_6473 (.A(\out_bs[3] [2]), .ZN(n_1_737_5634));
   INV_X1 i_1_737_6474 (.A(\out_bs[3] [3]), .ZN(n_1_737_5635));
   INV_X1 i_1_737_6475 (.A(\out_bs[3] [4]), .ZN(n_1_737_5636));
   INV_X1 i_1_737_6476 (.A(\out_bs[3] [5]), .ZN(n_1_737_5637));
   INV_X1 i_1_737_6477 (.A(\out_bs[3] [6]), .ZN(n_1_737_5638));
   INV_X1 i_1_737_6478 (.A(\out_as[2] [1]), .ZN(n_1_737_5639));
   INV_X1 i_1_737_6479 (.A(\out_as[2] [2]), .ZN(n_1_737_5640));
   INV_X1 i_1_737_6480 (.A(\out_as[2] [3]), .ZN(n_1_737_5641));
   INV_X1 i_1_737_6481 (.A(\out_as[2] [4]), .ZN(n_1_737_5642));
   INV_X1 i_1_737_6482 (.A(\out_as[2] [5]), .ZN(n_1_737_5643));
   INV_X1 i_1_737_6483 (.A(\out_as[2] [6]), .ZN(n_1_737_5644));
   INV_X1 i_1_737_6484 (.A(\out_bs[2] [0]), .ZN(n_1_737_5645));
   INV_X1 i_1_737_6485 (.A(\out_bs[2] [1]), .ZN(n_1_737_5646));
   INV_X1 i_1_737_6486 (.A(\out_bs[2] [2]), .ZN(n_1_737_5647));
   INV_X1 i_1_737_6487 (.A(\out_bs[2] [3]), .ZN(n_1_737_5648));
   INV_X1 i_1_737_6488 (.A(\out_bs[2] [4]), .ZN(n_1_737_5649));
   INV_X1 i_1_737_6489 (.A(\out_bs[2] [5]), .ZN(n_1_737_5650));
   INV_X1 i_1_737_6490 (.A(\out_bs[2] [6]), .ZN(n_1_737_5651));
   INV_X1 i_1_737_6491 (.A(\out_as[1] [0]), .ZN(n_1_737_5652));
   INV_X1 i_1_737_6492 (.A(\out_as[1] [1]), .ZN(n_1_737_5653));
   INV_X1 i_1_737_6493 (.A(\out_as[1] [2]), .ZN(n_1_737_5654));
   INV_X1 i_1_737_6494 (.A(\out_as[1] [3]), .ZN(n_1_737_5655));
   INV_X1 i_1_737_6495 (.A(\out_as[1] [4]), .ZN(n_1_737_5656));
   INV_X1 i_1_737_6496 (.A(\out_as[1] [5]), .ZN(n_1_737_5657));
   INV_X1 i_1_737_6497 (.A(\out_as[1] [6]), .ZN(n_1_737_5658));
   INV_X1 i_1_737_6498 (.A(\out_bs[1] [1]), .ZN(n_1_737_5659));
   INV_X1 i_1_737_6499 (.A(\out_bs[1] [2]), .ZN(n_1_737_5660));
   INV_X1 i_1_737_6500 (.A(\out_bs[1] [3]), .ZN(n_1_737_5661));
   INV_X1 i_1_737_6501 (.A(\out_bs[1] [4]), .ZN(n_1_737_5662));
   INV_X1 i_1_737_6502 (.A(\out_bs[1] [5]), .ZN(n_1_737_5663));
   INV_X1 i_1_737_6503 (.A(\out_bs[1] [6]), .ZN(n_1_737_5664));
   INV_X1 i_1_737_6504 (.A(\out_bs[0] [0]), .ZN(n_1_737_5665));
   INV_X1 i_1_737_6505 (.A(\out_bs[0] [1]), .ZN(n_1_737_5666));
   INV_X1 i_1_737_6506 (.A(\out_bs[0] [2]), .ZN(n_1_737_5667));
   INV_X1 i_1_737_6507 (.A(\out_bs[0] [3]), .ZN(n_1_737_5668));
   INV_X1 i_1_737_6508 (.A(\out_bs[0] [4]), .ZN(n_1_737_5669));
   INV_X1 i_1_737_6509 (.A(\out_bs[0] [5]), .ZN(n_1_737_5670));
   INV_X1 i_1_737_6510 (.A(\out_bs[0] [6]), .ZN(n_1_737_5671));
   INV_X1 i_1_737_6511 (.A(\out_as[0] [0]), .ZN(n_1_737_5672));
   INV_X1 i_1_737_6512 (.A(\out_as[0] [1]), .ZN(n_1_737_5673));
   INV_X1 i_1_737_6513 (.A(\out_as[0] [2]), .ZN(n_1_737_5674));
   INV_X1 i_1_737_6514 (.A(\out_as[0] [3]), .ZN(n_1_737_5675));
   INV_X1 i_1_737_6515 (.A(\out_as[0] [4]), .ZN(n_1_737_5676));
   INV_X1 i_1_737_6516 (.A(\out_as[0] [5]), .ZN(n_1_737_5677));
   INV_X1 i_1_737_6517 (.A(\out_as[0] [6]), .ZN(n_1_737_5678));
   OAI21_X1 i_1_737_6518 (.A(\out_bs[3] [5]), .B1(n_1_737_4427), .B2(
      n_1_737_4381), .ZN(n_1_737_5679));
   OAI21_X1 i_1_737_6519 (.A(\out_bs[2] [5]), .B1(n_1_737_4416), .B2(
      n_1_737_4387), .ZN(n_1_737_5680));
   NOR2_X1 i_1_737_1980 (.A1(n_844), .A2(n_845), .ZN(n_1_737_1870));
   NOR2_X1 i_1_737_1981 (.A1(n_1_737_5610), .A2(n_1_737_5609), .ZN(n_1_737_1871));
   INV_X1 i_1_737_1982 (.A(n_1_737_1871), .ZN(n_1_737_1874));
   NAND2_X1 i_1_737_1985 (.A1(n_1_737_1870), .A2(n_1_737_1874), .ZN(n_1_737_1875));
   INV_X1 i_1_737_1986 (.A(n_1_737_1875), .ZN(n_1_737_4402));
   INV_X1 i_1_737_2098 (.A(n_1_737_1870), .ZN(n_1_737_5181));
   INV_X1 i_1_737_2099 (.A(in_data[8]), .ZN(n_1_737_5596));
   INV_X1 i_1_737_2100 (.A(n_1_737_1974), .ZN(n_1_737_1973));
   NOR2_X1 i_1_737_2101 (.A1(n_1_737_5612), .A2(n_1_737_5611), .ZN(n_1_737_1969));
   NOR2_X1 i_1_737_2103 (.A1(n_1_737_4614), .A2(n_1_737_5610), .ZN(n_1_737_1979));
   INV_X1 i_1_737_2106 (.A(n_1089), .ZN(n_1_737_4400));
   AND2_X1 i_1_737_2108 (.A1(n_1_737_1969), .A2(n_1_737_1979), .ZN(n_1_737_5681));
   NOR2_X1 i_1_737_2109 (.A1(n_1_737_4400), .A2(n_1_737_5681), .ZN(n_1_737_1970));
   NOR2_X1 i_1_737_3495 (.A1(n_1_737_5608), .A2(n_1_737_5183), .ZN(n_1_737_5682));
   INV_X1 i_1_737_4641 (.A(n_1_737_5168), .ZN(n_1_737_5683));
   NAND2_X1 i_1_737_4987 (.A1(n_848), .A2(n_1_737_5682), .ZN(n_1_737_5684));
   NAND2_X1 i_1_737_4988 (.A1(n_1_737_1874), .A2(n_1_737_5684), .ZN(n_1_737_5685));
   NOR2_X1 i_1_737_4989 (.A1(n_1_737_5683), .A2(n_1_737_236), .ZN(n_1_737_5686));
   NOR4_X1 i_1_737_4990 (.A1(n_844), .A2(n_845), .A3(n_1_737_5685), .A4(
      n_1_737_5686), .ZN(n_1_737_5687));
   INV_X1 i_1_737_4991 (.A(n_1_737_5687), .ZN(n_832));
   OAI21_X1 i_1_737_4993 (.A(n_1_737_4454), .B1(n_1_737_5366), .B2(n_1_737_4455), 
      .ZN(n_1_737_5688));
   NOR3_X1 i_1_737_5043 (.A1(n_844), .A2(n_845), .A3(n_1_737_5685), .ZN(
      n_1_737_5689));
   NOR3_X1 i_1_737_5618 (.A1(n_1_737_5689), .A2(n_1_737_5683), .A3(n_1_737_236), 
      .ZN(n_1_737_5690));
   NOR2_X1 i_1_737_5809 (.A1(n_1089), .A2(n_1_737_5687), .ZN(n_1_737_5691));
   AOI211_X1 i_1_737_5817 (.A(n_1_737_1872), .B(n_1_737_5688), .C1(n_1_737_4417), 
      .C2(n_1_737_5598), .ZN(n_1_737_5692));
   AND2_X1 i_1_737_5819 (.A1(n_1_737_5688), .A2(in_data[12]), .ZN(n_1_737_5693));
   NOR4_X1 i_1_737_5917 (.A1(n_1_737_5691), .A2(n_1_737_5692), .A3(n_1_737_5690), 
      .A4(n_1_737_5693), .ZN(n_1_737_5694));
   INV_X1 i_1_737_5931 (.A(n_1_737_5691), .ZN(n_1_737_5695));
   INV_X1 i_1_737_5932 (.A(n_1_737_5690), .ZN(n_1_737_5696));
   AOI21_X1 i_1_737_6088 (.A(in_data[8]), .B1(n_1_737_5695), .B2(n_1_737_5696), 
      .ZN(n_1_737_5697));
   NOR2_X1 i_1_737_6379 (.A1(n_1_737_5694), .A2(n_1_737_5697), .ZN(n_833));
   OAI21_X1 i_1_737_6394 (.A(n_1_737_5190), .B1(n_1_737_5191), .B2(n_1_737_3150), 
      .ZN(n_1_737_5698));
   OAI21_X1 i_1_737_6434 (.A(n_1_737_5236), .B1(n_1_737_5237), .B2(n_1_737_3160), 
      .ZN(n_1_737_5699));
   INV_X1 i_1_737_6440 (.A(n_1_737_1972), .ZN(n_1_737_1971));
   OAI21_X1 i_1_737_6520 (.A(n_1_737_5338), .B1(\out_as[0] [6]), .B2(
      n_1_737_5339), .ZN(n_1_737_5700));
   NOR4_X1 i_1_737_6521 (.A1(n_1_737_4400), .A2(n_1_737_5698), .A3(n_1_737_5699), 
      .A4(n_1_737_5681), .ZN(n_1_737_5701));
   INV_X1 i_1_737_6522 (.A(n_1_737_5700), .ZN(n_1_737_5702));
   NOR2_X1 i_1_737_6523 (.A1(n_1_737_5338), .A2(n_1_737_3163), .ZN(n_1_737_5703));
   NOR4_X1 i_1_737_6524 (.A1(n_1_737_1974), .A2(n_1_737_1972), .A3(n_1_737_5702), 
      .A4(n_1_737_5703), .ZN(n_1_737_5704));
   NAND2_X1 i_1_737_6525 (.A1(n_1_737_5701), .A2(n_1_737_5704), .ZN(n_834));
   INV_X1 i_1_737_6526 (.A(n_1_737_80), .ZN(n_1_737_5705));
   OR2_X1 i_1_737_6527 (.A1(n_955), .A2(n_1_737_5705), .ZN(n_835));
   INV_X1 i_1_737_6528 (.A(n_1_737_44), .ZN(n_1_737_5706));
   OR2_X1 i_1_737_6529 (.A1(n_962), .A2(n_1_737_5706), .ZN(n_836));
   OR2_X1 i_1_737_6530 (.A1(\out_bs[7] [6]), .A2(n_970), .ZN(n_837));
   BUF_X1 i_1_737_6531 (.A(n_1_737_1870), .Z(n_1_737_5182));
   BUF_X1 i_1_737_6532 (.A(n_1_737_1875), .Z(n_1_737_4401));
   BUF_X1 i_1_737_6533 (.A(n_1_737_1871), .Z(n_1_737_4404));
   BUF_X1 i_1_737_6534 (.A(n_1_737_1969), .Z(n_1_737_3110));
   BUF_X1 i_1_737_6535 (.A(n_1_737_1979), .Z(n_1_737_4092));
   BUF_X1 i_1_737_6536 (.A(n_1_737_4400), .Z(n_1_737_5602));
   BUF_X1 i_1_737_6537 (.A(n_1_737_5682), .Z(n_1_737_4965));
   BUF_X1 i_1_737_6538 (.A(n_1_737_5683), .Z(n_1_737_5167));
   BUF_X1 i_1_737_6539 (.A(n_1_737_5688), .Z(n_1_737_4453));
   BUF_X1 i_1_737_6540 (.A(n_1_737_5690), .Z(n_838));
   BUF_X1 i_1_737_6541 (.A(n_1_737_5698), .Z(n_1_737_1978));
   BUF_X1 i_1_737_6542 (.A(n_1_737_5699), .Z(n_1_737_1976));
   BUF_X1 i_1_737_6543 (.A(n_1_737_5700), .Z(n_1_737_5337));
   BUF_X1 i_1_737_6544 (.A(n_1_737_5705), .Z(n_839));
   BUF_X1 i_1_737_6545 (.A(n_1_737_5706), .Z(n_840));
   OAI21_X1 i_4_1_0 (.A(n_4_1_0), .B1(n_952), .B2(n_4_1_1), .ZN(n_841));
   AOI21_X1 i_4_1_1 (.A(n_4_0), .B1(n_952), .B2(n_4_1), .ZN(n_4_1_0));
   INV_X1 i_4_1_2 (.A(n_4_2), .ZN(n_4_1_1));
   OAI21_X1 i_4_513_0 (.A(n_4_513_0), .B1(n_4_513_3), .B2(n_4_513_1), .ZN(n_842));
   NAND2_X1 i_4_513_1 (.A1(n_128), .A2(n_4_513_1), .ZN(n_4_513_0));
   OAI22_X1 i_4_513_2 (.A1(n_952), .A2(n_4_2), .B1(n_4_513_2), .B2(n_4_1), 
      .ZN(n_4_513_1));
   INV_X1 i_4_513_3 (.A(n_952), .ZN(n_4_513_2));
   INV_X1 i_4_513_4 (.A(in_data[4]), .ZN(n_4_513_3));
   OAI21_X1 i_4_54_0 (.A(n_4_54_0), .B1(n_1011), .B2(n_4_54_1), .ZN(n_4_0));
   AOI21_X1 i_4_54_1 (.A(n_745), .B1(n_1011), .B2(n_743), .ZN(n_4_54_0));
   INV_X1 i_4_54_2 (.A(n_744), .ZN(n_4_54_1));
   AND2_X1 i_4_56_0 (.A1(n_739), .A2(n_4_3), .ZN(n_4_1));
   OR2_X1 i_4_57_0 (.A1(n_4_3), .A2(n_739), .ZN(n_4_2));
   datapath__1_13511 i_4_55 (.to_int5359({1'b0, n_843, n_1312, n_850, n_847, 
      n_851, n_1311, \out_bs[6] [0]}), .p_0(n_4_3));
   BUF_X1 rt_shieldBuf (.A(\out_bs[6] [6]), .Z(n_843));
   BUF_X1 rt_shieldBuf__0 (.A(\out_bs[5] [6]), .Z(n_844));
   BUF_X1 rt_shieldBuf__1 (.A(\out_bs[5] [5]), .Z(n_845));
   BUF_X1 rt_shieldBuf__2 (.A(\out_bs[5] [3]), .Z(n_846));
   BUF_X1 rt_shieldBuf__3 (.A(\out_bs[6] [3]), .Z(n_847));
   BUF_X1 rt_shieldBuf__4 (.A(\out_bs[5] [4]), .Z(n_848));
   BUF_X1 rt_shieldBuf__5 (.A(\out_bs[5] [2]), .Z(n_849));
   BUF_X1 rt_shieldBuf__6 (.A(\out_bs[6] [4]), .Z(n_850));
   BUF_X1 rt_shieldBuf__7 (.A(\out_bs[6] [2]), .Z(n_851));
   datapath__1_7666 i_0_0 (.to_int6126({uc_0, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_2));
   AND2_X1 i_0_1_0 (.A1(n_0), .A2(n_0_2), .ZN(n_0_129));
   OR2_X1 i_0_2_0 (.A1(n_0_2), .A2(n_0), .ZN(n_0_390));
   datapath__1_7740 i_0_3 (.to_int6126({uc_1, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_5));
   datapath__1_18134 i_0_4 (.to_int6126({1'b0, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_0));
   datapath__1_14001 i_0_5 (.to_int6126({uc_2, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_711));
   datapath__1_13985 i_0_6 (.to_int6126({uc_3, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_701));
   datapath__1_13961 i_0_7 (.to_int6126({uc_4, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_688));
   datapath__1_13953 i_0_8 (.to_int6126({uc_5, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_683));
   datapath__1_13945 i_0_9 (.to_int6126({uc_6, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_677));
   datapath__1_13937 i_0_10 (.to_int6126({uc_7, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_672));
   datapath__1_13929 i_0_11 (.to_int6126({uc_8, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_667));
   datapath__1_13913 i_0_12 (.to_int6126({uc_9, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_657));
   datapath__1_13905 i_0_13 (.to_int6126({uc_10, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_651));
   datapath__1_13897 i_0_14 (.to_int6126({uc_11, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_645));
   datapath__1_13889 i_0_15 (.to_int6126({uc_12, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_639));
   datapath__1_13881 i_0_16 (.to_int6126({uc_13, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_633));
   datapath__1_13873 i_0_17 (.to_int6126({uc_14, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_627));
   datapath__1_13865 i_0_18 (.to_int6126({uc_15, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_621));
   datapath__1_13857 i_0_19 (.to_int6126({uc_16, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_615));
   datapath__1_13849 i_0_20 (.to_int6126({uc_17, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_609));
   datapath__1_13841 i_0_21 (.to_int6126({uc_18, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_603));
   datapath__1_13833 i_0_22 (.to_int6126({uc_19, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_597));
   datapath__1_13825 i_0_23 (.to_int6126({uc_20, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_592));
   datapath__1_13817 i_0_24 (.to_int6126({uc_21, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_586));
   datapath__1_13809 i_0_25 (.to_int6126({1'b0, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_580));
   datapath__1_13801 i_0_26 (.to_int6126({1'b0, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_574));
   datapath__1_13793 i_0_27 (.to_int6126({uc_22, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_568));
   datapath__1_13785 i_0_28 (.to_int6126({uc_23, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_562));
   datapath__1_13777 i_0_29 (.to_int6126({uc_24, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_556));
   datapath__1_13769 i_0_30 (.to_int6126({uc_25, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_550));
   datapath__1_13762 i_0_31 (.to_int6126({uc_26, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_545));
   datapath__1_13754 i_0_32 (.to_int6126({uc_27, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_541));
   datapath__1_13746 i_0_33 (.to_int6126({uc_28, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_535));
   datapath__1_13738 i_0_34 (.to_int6126({uc_29, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_529));
   datapath__1_13730 i_0_35 (.to_int6126({1'b0, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_523));
   datapath__1_13722 i_0_36 (.to_int6126({1'b0, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_517));
   datapath__1_13714 i_0_37 (.to_int6126({uc_30, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_511));
   datapath__1_13706 i_0_38 (.to_int6126({uc_31, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_505));
   datapath__1_13698 i_0_39 (.to_int6126({1'b0, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_499));
   datapath__1_13690 i_0_40 (.to_int6126({uc_32, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_493));
   datapath__1_13682 i_0_41 (.to_int6126({1'b0, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_487));
   datapath__1_13674 i_0_42 (.to_int6126({1'b0, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_481));
   datapath__1_13666 i_0_43 (.to_int6126({uc_33, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_475));
   datapath__1_13658 i_0_44 (.to_int6126({uc_34, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_469));
   datapath__1_13650 i_0_45 (.to_int6126({uc_35, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_463));
   datapath__1_13642 i_0_46 (.to_int6126({uc_36, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_457));
   datapath__1_13634 i_0_47 (.to_int6126({uc_37, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_452));
   datapath__1_13626 i_0_48 (.to_int6126({uc_38, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_449));
   datapath__1_13618 i_0_49 (.to_int6126({uc_39, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_443));
   datapath__1_13610 i_0_50 (.to_int6126({uc_40, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_437));
   datapath__1_13602 i_0_51 (.to_int6126({uc_41, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_432));
   datapath__1_13594 i_0_52 (.to_int6126({uc_42, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_426));
   datapath__1_13586 i_0_53 (.to_int6126({uc_43, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_420));
   datapath__1_13578 i_0_54 (.to_int6126({uc_44, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_414));
   datapath__1_13562 i_0_55 (.to_int6126({uc_45, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_408));
   datapath__1_13538 i_0_56 (.to_int6126({uc_46, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 
      \out_bs[7] [0]}), .p_0(n_0_403));
   datapath__1_13997 i_0_57 (.to_int6126({uc_47, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], uc_48}), 
      .p_0(n_0_708));
   datapath__1_13949 i_0_58 (.to_int6126({uc_49, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], uc_50}), 
      .p_0(n_0_680));
   datapath__1_13901 i_0_59 (.to_int6126({uc_51, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], uc_52}), 
      .p_0(n_0_648));
   datapath__1_13885 i_0_60 (.to_int6126({uc_53, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], uc_54}), 
      .p_0(n_0_636));
   datapath__1_13869 i_0_61 (.to_int6126({uc_55, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], uc_56}), 
      .p_0(n_0_624));
   datapath__1_13853 i_0_62 (.to_int6126({1'b0, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 1'b0}), 
      .p_0(n_0_612));
   datapath__1_13837 i_0_63 (.to_int6126({1'b0, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 1'b0}), 
      .p_0(n_0_600));
   datapath__1_13821 i_0_64 (.to_int6126({uc_57, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], uc_58}), 
      .p_0(n_0_589));
   datapath__1_13805 i_0_65 (.to_int6126({uc_59, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], uc_60}), 
      .p_0(n_0_577));
   datapath__1_13789 i_0_66 (.to_int6126({uc_61, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], uc_62}), 
      .p_0(n_0_565));
   datapath__1_13773 i_0_67 (.to_int6126({uc_63, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], uc_64}), 
      .p_0(n_0_553));
   datapath__1_13758 i_0_68 (.to_int6126({uc_65, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], uc_66}), 
      .p_0(n_0_544));
   datapath__1_13742 i_0_69 (.to_int6126({1'b0, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 1'b0}), 
      .p_0(n_0_532));
   datapath__1_13726 i_0_70 (.to_int6126({uc_67, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], uc_68}), 
      .p_0(n_0_520));
   datapath__1_13710 i_0_71 (.to_int6126({uc_69, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], uc_70}), 
      .p_0(n_0_508));
   datapath__1_13694 i_0_72 (.to_int6126({1'b0, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 1'b0}), 
      .p_0(n_0_496));
   datapath__1_13678 i_0_73 (.to_int6126({1'b0, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], 1'b0}), 
      .p_0(n_0_484));
   datapath__1_13662 i_0_74 (.to_int6126({uc_71, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], uc_72}), 
      .p_0(n_0_472));
   datapath__1_13646 i_0_75 (.to_int6126({uc_73, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], uc_74}), 
      .p_0(n_0_460));
   datapath__1_13614 i_0_76 (.to_int6126({uc_75, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], uc_76}), 
      .p_0(n_0_440));
   datapath__1_13598 i_0_77 (.to_int6126({uc_77, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], uc_78}), 
      .p_0(n_0_429));
   datapath__1_13582 i_0_78 (.to_int6126({uc_79, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], uc_80}), 
      .p_0(n_0_417));
   datapath__1_13566 i_0_79 (.to_int6126({uc_81, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], uc_82}), 
      .p_0(n_0_411));
   datapath__1_13550 i_0_80 (.to_int6126({uc_83, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], uc_84}), 
      .p_0(n_0_405));
   datapath__1_13534 i_0_81 (.to_int6126({uc_85, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], uc_86}), 
      .p_0(n_0_400));
   datapath__1_13519 i_0_82 (.to_int6126({uc_87, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], \out_bs[7] [1], uc_88}), 
      .p_0(n_0_392));
   datapath__1_13909 i_0_83 (.to_int6126({uc_89, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], uc_90, uc_91}), .p_0(
      n_0_654));
   datapath__1_13877 i_0_84 (.to_int6126({uc_92, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], uc_93, uc_94}), .p_0(
      n_0_630));
   datapath__1_13845 i_0_85 (.to_int6126({uc_95, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], uc_96, uc_97}), .p_0(
      n_0_606));
   datapath__1_13813 i_0_86 (.to_int6126({uc_98, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], uc_99, uc_100}), .p_0(
      n_0_583));
   datapath__1_13781 i_0_87 (.to_int6126({uc_101, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], uc_102, uc_103}), .p_0(
      n_0_559));
   datapath__1_13750 i_0_88 (.to_int6126({uc_104, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], uc_105, uc_106}), .p_0(
      n_0_538));
   datapath__1_13718 i_0_89 (.to_int6126({uc_107, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], uc_108, uc_109}), .p_0(
      n_0_514));
   datapath__1_13686 i_0_90 (.to_int6126({uc_110, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], uc_111, uc_112}), .p_0(
      n_0_490));
   datapath__1_13654 i_0_91 (.to_int6126({uc_113, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], uc_114, uc_115}), .p_0(
      n_0_466));
   datapath__1_13622 i_0_92 (.to_int6126({uc_116, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], uc_117, uc_118}), .p_0(
      n_0_446));
   datapath__1_13590 i_0_93 (.to_int6126({uc_119, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], uc_120, uc_121}), .p_0(
      n_0_423));
   datapath__1_13558 i_0_94 (.to_int6126({uc_122, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], uc_123, uc_124}), .p_0(
      n_852));
   datapath__1_13526 i_0_95 (.to_int6126({uc_125, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], uc_126, uc_127}), .p_0(
      n_0_397));
   datapath__1_13925 i_0_96 (.to_int6126({uc_128, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], uc_129, uc_130, uc_131}), .p_0(n_0_664));
   datapath__1_13861 i_0_97 (.to_int6126({1'b0, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], 1'b0, 1'b0, 1'b0}), .p_0(n_0_618));
   datapath__1_13797 i_0_98 (.to_int6126({1'b0, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], 1'b0, 1'b0, 1'b0}), .p_0(n_0_571));
   datapath__1_13734 i_0_99 (.to_int6126({uc_132, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], uc_133, uc_134, uc_135}), .p_0(n_0_526));
   datapath__1_13670 i_0_100 (.to_int6126({1'b0, \out_bs[7] [6], \out_bs[7] [5], 
      \out_bs[7] [4], \out_bs[7] [3], 1'b0, 1'b0, 1'b0}), .p_0(n_0_478));
   datapath__1_13606 i_0_101 (.to_int6126({uc_136, \out_bs[7] [6], 
      \out_bs[7] [5], \out_bs[7] [4], \out_bs[7] [3], uc_137, uc_138, uc_139}), 
      .p_0(n_853));
   datapath__1_13542 i_0_102 (.to_int6126({uc_140, \out_bs[7] [6], 
      \out_bs[7] [5], \out_bs[7] [4], \out_bs[7] [3], uc_141, uc_142, uc_143}), 
      .p_0(n_0_404));
   datapath__1_13702 i_0_103 (.to_int6126({uc_144, \out_bs[7] [6], 
      \out_bs[7] [5], \out_bs[7] [4], uc_145, uc_146, uc_147, uc_148}), .p_0(
      n_0_502));
   datapath__1_13893 i_0_104 (.to_int6126({1'b0, \out_bs[7] [6], \out_bs[7] [5], 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0}), .p_0(n_0_642));
   AND2_X1 i_0_105_0 (.A1(n_970), .A2(\out_bs[7] [6]), .ZN(n_0_1));
   INV_X1 i_0_106_0 (.A(n_0_106_0), .ZN(n_0_128));
   OAI21_X1 i_0_106_1 (.A(n_0_106_1), .B1(n_842), .B2(n_0_129), .ZN(n_0_106_0));
   NAND2_X1 i_0_106_2 (.A1(n_0_129), .A2(n_0_106_2), .ZN(n_0_106_1));
   INV_X1 i_0_106_3 (.A(in_data[0]), .ZN(n_0_106_2));
   OR2_X1 i_0_107_0 (.A1(n_1213), .A2(n_132), .ZN(n_0_131));
   OR2_X1 i_0_107_4 (.A1(n_1266), .A2(n_0_78), .ZN(n_0_137));
   OR2_X1 i_0_107_5 (.A1(n_1265), .A2(n_0_125), .ZN(n_0_138));
   OR2_X1 i_0_107_6 (.A1(n_1264), .A2(n_0_127), .ZN(n_0_139));
   OR2_X1 i_0_107_11 (.A1(n_1261), .A2(n_0_76), .ZN(n_0_145));
   OR2_X1 i_0_107_14 (.A1(n_1258), .A2(n_0_75), .ZN(n_0_149));
   OR2_X1 i_0_107_15 (.A1(n_1257), .A2(n_0_52), .ZN(n_0_150));
   OR2_X1 i_0_107_16 (.A1(n_1256), .A2(n_0_90), .ZN(n_0_151));
   OR2_X1 i_0_107_18 (.A1(n_1255), .A2(n_0_74), .ZN(n_0_153));
   OR2_X1 i_0_107_19 (.A1(n_1254), .A2(n_0_50), .ZN(n_0_154));
   OR2_X1 i_0_107_20 (.A1(n_1253), .A2(n_1309), .ZN(n_0_155));
   OR2_X1 i_0_107_22 (.A1(n_1021), .A2(n_0_73), .ZN(n_0_157));
   OR2_X1 i_0_107_26 (.A1(n_1250), .A2(n_0_46), .ZN(n_0_162));
   OR2_X1 i_0_107_31 (.A1(n_1249), .A2(n_0_43), .ZN(n_0_168));
   OR2_X1 i_0_107_32 (.A1(n_1248), .A2(n_0_71), .ZN(n_0_169));
   OR2_X1 i_0_107_33 (.A1(n_1029), .A2(n_0_97), .ZN(n_0_171));
   OR2_X1 i_0_107_34 (.A1(n_1030), .A2(n_0_41), .ZN(n_0_172));
   OR2_X1 i_0_107_35 (.A1(n_1031), .A2(n_0_70), .ZN(n_0_173));
   OR2_X1 i_0_107_36 (.A1(n_1032), .A2(n_0_40), .ZN(n_0_174));
   OR2_X1 i_0_107_37 (.A1(n_1246), .A2(n_0_87), .ZN(n_0_175));
   OR2_X1 i_0_107_38 (.A1(n_1033), .A2(n_0_39), .ZN(n_0_176));
   OR2_X1 i_0_107_39 (.A1(n_1034), .A2(n_0_69), .ZN(n_0_177));
   OR2_X1 i_0_107_40 (.A1(n_1035), .A2(n_0_38), .ZN(n_0_178));
   OR2_X1 i_0_107_43 (.A1(n_1245), .A2(n_0_36), .ZN(n_0_182));
   OR2_X1 i_0_107_44 (.A1(n_1039), .A2(n_0_86), .ZN(n_0_183));
   OR2_X1 i_0_107_45 (.A1(n_1040), .A2(n_0_35), .ZN(n_0_184));
   OR2_X1 i_0_107_46 (.A1(n_1244), .A2(n_0_67), .ZN(n_0_185));
   OR2_X1 i_0_107_47 (.A1(n_1041), .A2(n_0_34), .ZN(n_0_186));
   OR2_X1 i_0_107_48 (.A1(n_1042), .A2(n_0_96), .ZN(n_0_187));
   OR2_X1 i_0_107_49 (.A1(n_1243), .A2(n_0_33), .ZN(n_0_188));
   OR2_X1 i_0_107_50 (.A1(n_1043), .A2(n_0_66), .ZN(n_0_189));
   OR2_X1 i_0_107_51 (.A1(n_1242), .A2(n_0_32), .ZN(n_0_190));
   OR2_X1 i_0_107_53 (.A1(n_1241), .A2(n_0_31), .ZN(n_0_192));
   OR2_X1 i_0_107_54 (.A1(n_1240), .A2(n_0_126), .ZN(n_0_193));
   OR2_X1 i_0_107_55 (.A1(n_1239), .A2(n_0_30), .ZN(n_0_194));
   OR2_X1 i_0_107_59 (.A1(n_1047), .A2(n_0_84), .ZN(n_0_199));
   OR2_X1 i_0_107_63 (.A1(n_1051), .A2(n_0_95), .ZN(n_0_203));
   OR2_X1 i_0_107_66 (.A1(n_1054), .A2(n_0_24), .ZN(n_0_206));
   OR2_X1 i_0_107_69 (.A1(n_1236), .A2(n_0_62), .ZN(n_0_209));
   OR2_X1 i_0_107_70 (.A1(n_1235), .A2(n_0_22), .ZN(n_0_210));
   OR2_X1 i_0_107_71 (.A1(n_1057), .A2(n_0_117), .ZN(n_0_211));
   OR2_X1 i_0_107_72 (.A1(n_1234), .A2(n_0_21), .ZN(n_0_212));
   OR2_X1 i_0_107_73 (.A1(n_1058), .A2(n_0_61), .ZN(n_0_213));
   OR2_X1 i_0_107_74 (.A1(n_1233), .A2(n_0_20), .ZN(n_0_214));
   OR2_X1 i_0_107_75 (.A1(n_1232), .A2(n_0_82), .ZN(n_0_215));
   OR2_X1 i_0_107_76 (.A1(n_1231), .A2(n_0_19), .ZN(n_0_216));
   OR2_X1 i_0_107_78 (.A1(n_1060), .A2(n_0_18), .ZN(n_0_218));
   OR2_X1 i_0_107_79 (.A1(n_1061), .A2(n_0_94), .ZN(n_0_219));
   OR2_X1 i_0_107_80 (.A1(n_1062), .A2(n_0_17), .ZN(n_0_220));
   OR2_X1 i_0_107_86 (.A1(n_1228), .A2(n_0_99), .ZN(n_0_227));
   OR2_X1 i_0_107_89 (.A1(n_1227), .A2(n_0_12), .ZN(n_0_230));
   OR2_X1 i_0_107_92 (.A1(n_1071), .A2(n_0_111), .ZN(n_0_233));
   OR2_X1 i_0_107_93 (.A1(n_1226), .A2(n_0_106), .ZN(n_0_234));
   OR2_X1 i_0_107_95 (.A1(n_1224), .A2(n_0_10), .ZN(n_0_236));
   OR2_X1 i_0_107_98 (.A1(n_1222), .A2(n_0_114), .ZN(n_0_239));
   OR2_X1 i_0_107_101 (.A1(n_1221), .A2(n_0_116), .ZN(n_0_243));
   OR2_X1 i_0_107_102 (.A1(n_1220), .A2(n_0_6), .ZN(n_0_244));
   OR2_X1 i_0_107_103 (.A1(n_1219), .A2(n_0_109), .ZN(n_0_245));
   OR2_X1 i_0_107_104 (.A1(n_1076), .A2(n_0_105), .ZN(n_0_246));
   OR2_X1 i_0_107_105 (.A1(n_1218), .A2(n_0_113), .ZN(n_0_247));
   OR2_X1 i_0_107_107 (.A1(n_1078), .A2(n_0_108), .ZN(n_0_249));
   OR2_X1 i_0_107_110 (.A1(n_1216), .A2(n_0_112), .ZN(n_0_255));
   NAND2_X1 i_0_107_117 (.A1(n_0_107_1), .A2(n_0_107_0), .ZN(n_0_143));
   INV_X1 i_0_107_118 (.A(n_1016), .ZN(n_0_107_0));
   INV_X1 i_0_107_119 (.A(n_0_91), .ZN(n_0_107_1));
   OR2_X1 i_0_107_1 (.A1(n_0_129), .A2(n_841), .ZN(n_0_132));
   OR2_X1 i_0_107_2 (.A1(n_0_79), .A2(n_1012), .ZN(n_0_133));
   OR2_X1 i_0_107_3 (.A1(n_0_130), .A2(n_1013), .ZN(n_0_134));
   OR2_X1 i_0_107_7 (.A1(n_0_92), .A2(n_1014), .ZN(n_0_135));
   OR2_X1 i_0_107_8 (.A1(n_1275), .A2(n_1267), .ZN(n_0_136));
   OR2_X1 i_0_107_9 (.A1(n_1278), .A2(n_1263), .ZN(n_0_140));
   OR2_X1 i_0_107_10 (.A1(n_0_77), .A2(n_1015), .ZN(n_0_141));
   OR2_X1 i_0_107_12 (.A1(n_1281), .A2(n_1262), .ZN(n_0_142));
   OR2_X1 i_0_107_13 (.A1(n_0_54), .A2(n_1017), .ZN(n_0_144));
   OR2_X1 i_0_107_17 (.A1(n_1289), .A2(n_1260), .ZN(n_0_146));
   OR2_X1 i_0_107_21 (.A1(n_1310), .A2(n_1259), .ZN(n_0_147));
   OR2_X1 i_0_107_23 (.A1(n_0_53), .A2(n_1018), .ZN(n_0_148));
   OR2_X1 i_0_107_24 (.A1(n_0_51), .A2(n_1019), .ZN(n_0_152));
   OR2_X1 i_0_107_25 (.A1(n_0_49), .A2(n_1020), .ZN(n_0_156));
   OR2_X1 i_0_107_27 (.A1(n_0_48), .A2(n_1022), .ZN(n_0_158));
   OR2_X1 i_0_107_28 (.A1(n_0_89), .A2(n_1252), .ZN(n_0_159));
   OR2_X1 i_0_107_29 (.A1(n_0_47), .A2(n_1023), .ZN(n_0_160));
   OR2_X1 i_0_107_30 (.A1(n_1287), .A2(n_1251), .ZN(n_0_161));
   OR2_X1 i_0_107_41 (.A1(n_0_118), .A2(n_1024), .ZN(n_0_163));
   OR2_X1 i_0_107_42 (.A1(n_0_45), .A2(n_1025), .ZN(n_0_164));
   OR2_X1 i_0_107_52 (.A1(n_0_72), .A2(n_1026), .ZN(n_0_165));
   OR2_X1 i_0_107_56 (.A1(n_0_44), .A2(n_1027), .ZN(n_0_166));
   OR2_X1 i_0_107_57 (.A1(n_0_88), .A2(n_1028), .ZN(n_0_167));
   OR2_X1 i_0_107_58 (.A1(n_0_42), .A2(n_1247), .ZN(n_0_170));
   OR2_X1 i_0_107_60 (.A1(n_0_98), .A2(n_1036), .ZN(n_0_179));
   OR2_X1 i_0_107_61 (.A1(n_0_37), .A2(n_1037), .ZN(n_0_180));
   OR2_X1 i_0_107_62 (.A1(n_0_68), .A2(n_1038), .ZN(n_0_181));
   OR2_X1 i_0_107_64 (.A1(n_0_85), .A2(n_1044), .ZN(n_0_191));
   OR2_X1 i_0_107_65 (.A1(n_0_1), .A2(n_1238), .ZN(n_0_195));
   OR2_X1 i_0_107_67 (.A1(n_0_29), .A2(n_1237), .ZN(n_0_196));
   OR2_X1 i_0_107_68 (.A1(n_0_65), .A2(n_1045), .ZN(n_0_197));
   OR2_X1 i_0_107_77 (.A1(n_0_28), .A2(n_1046), .ZN(n_0_198));
   OR2_X1 i_0_107_81 (.A1(n_0_27), .A2(n_1048), .ZN(n_0_200));
   OR2_X1 i_0_107_82 (.A1(n_0_64), .A2(n_1049), .ZN(n_0_201));
   OR2_X1 i_0_107_83 (.A1(n_0_26), .A2(n_1050), .ZN(n_0_202));
   OR2_X1 i_0_107_84 (.A1(n_0_25), .A2(n_1052), .ZN(n_0_204));
   OR2_X1 i_0_107_85 (.A1(n_0_63), .A2(n_1053), .ZN(n_0_205));
   OR2_X1 i_0_107_87 (.A1(n_0_83), .A2(n_1055), .ZN(n_0_207));
   OR2_X1 i_0_107_88 (.A1(n_0_23), .A2(n_1056), .ZN(n_0_208));
   OR2_X1 i_0_107_90 (.A1(n_0_60), .A2(n_1059), .ZN(n_0_217));
   OR2_X1 i_0_107_91 (.A1(n_0_59), .A2(n_1063), .ZN(n_0_221));
   OR2_X1 i_0_107_94 (.A1(n_0_16), .A2(n_1064), .ZN(n_0_222));
   OR2_X1 i_0_107_96 (.A1(n_0_81), .A2(n_1230), .ZN(n_0_223));
   OR2_X1 i_0_107_97 (.A1(n_0_15), .A2(n_1065), .ZN(n_0_224));
   OR2_X1 i_0_107_99 (.A1(n_0_58), .A2(n_1066), .ZN(n_0_225));
   OR2_X1 i_0_107_100 (.A1(n_0_14), .A2(n_1229), .ZN(n_0_226));
   OR2_X1 i_0_107_106 (.A1(n_0_13), .A2(n_1067), .ZN(n_0_228));
   OR2_X1 i_0_107_108 (.A1(n_0_57), .A2(n_1068), .ZN(n_0_229));
   OR2_X1 i_0_107_109 (.A1(n_0_80), .A2(n_1069), .ZN(n_0_231));
   OR2_X1 i_0_107_111 (.A1(n_0_11), .A2(n_1070), .ZN(n_0_232));
   OR2_X1 i_0_107_112 (.A1(n_0_93), .A2(n_1225), .ZN(n_0_235));
   OR2_X1 i_0_107_113 (.A1(n_0_110), .A2(n_1223), .ZN(n_0_237));
   OR2_X1 i_0_107_114 (.A1(n_0_9), .A2(n_1072), .ZN(n_0_238));
   OR2_X1 i_0_107_115 (.A1(n_0_8), .A2(n_1073), .ZN(n_0_240));
   OR2_X1 i_0_107_116 (.A1(n_0_56), .A2(n_1074), .ZN(n_0_241));
   OR2_X1 i_0_107_120 (.A1(n_0_7), .A2(n_1075), .ZN(n_0_242));
   OR2_X1 i_0_107_121 (.A1(n_0_104), .A2(n_1077), .ZN(n_0_248));
   OR2_X1 i_0_107_122 (.A1(n_0_4), .A2(n_1079), .ZN(n_0_250));
   OR2_X1 i_0_107_123 (.A1(n_0_115), .A2(n_1217), .ZN(n_0_251));
   OR2_X1 i_0_107_124 (.A1(n_0_103), .A2(n_1080), .ZN(n_0_252));
   OR2_X1 i_0_107_125 (.A1(n_0_55), .A2(n_1081), .ZN(n_0_253));
   OR2_X1 i_0_107_126 (.A1(n_0_3), .A2(n_1082), .ZN(n_0_254));
   OR2_X1 i_0_107_127 (.A1(n_0_102), .A2(n_1083), .ZN(n_0_256));
   OR2_X1 i_0_107_128 (.A1(n_0_107), .A2(n_1215), .ZN(n_0_257));
   OR2_X1 i_0_107_129 (.A1(n_0_0), .A2(n_1214), .ZN(n_0_258));
   INV_X1 i_0_108_0 (.A(n_0_108_0), .ZN(n_0_259));
   OAI21_X1 i_0_108_1 (.A(n_0_108_1), .B1(n_842), .B2(n_0_390), .ZN(n_0_108_0));
   NAND2_X1 i_0_108_2 (.A1(n_0_390), .A2(n_0_108_2), .ZN(n_0_108_1));
   INV_X1 i_0_108_3 (.A(in_data[0]), .ZN(n_0_108_2));
   OR2_X1 i_0_109_0 (.A1(n_841), .A2(n_0_390), .ZN(n_0_260));
   AND2_X1 i_0_110_0 (.A1(n_0_5), .A2(n_1), .ZN(n_0_130));
   OR2_X1 i_0_111_0 (.A1(n_0_5), .A2(n_1), .ZN(n_0_395));
   INV_X1 i_0_112_0 (.A(n_0_0), .ZN(n_0_112_0));
   AOI22_X1 i_0_112_1 (.A1(n_0_112_0), .A2(n_2), .B1(in_data[0]), .B2(n_0_0), 
      .ZN(n_0_112_1));
   INV_X1 i_0_112_2 (.A(n_0_112_1), .ZN(n_0_261));
   AND2_X1 i_0_113_0 (.A1(n_774), .A2(n_0_711), .ZN(n_0_3));
   OR2_X1 i_0_114_0 (.A1(n_0_711), .A2(n_774), .ZN(n_0_712));
   AND2_X1 i_0_115_0 (.A1(n_778), .A2(n_0_701), .ZN(n_0_4));
   OR2_X1 i_0_116_0 (.A1(n_0_701), .A2(n_778), .ZN(n_0_702));
   AND2_X1 i_0_117_0 (.A1(n_783), .A2(n_0_688), .ZN(n_0_6));
   OR2_X1 i_0_118_0 (.A1(n_0_688), .A2(n_783), .ZN(n_0_689));
   AND2_X1 i_0_119_0 (.A1(n_785), .A2(n_0_683), .ZN(n_0_7));
   OR2_X1 i_0_120_0 (.A1(n_0_683), .A2(n_785), .ZN(n_0_684));
   AND2_X1 i_0_121_0 (.A1(n_787), .A2(n_0_677), .ZN(n_0_8));
   OR2_X1 i_0_122_0 (.A1(n_0_677), .A2(n_787), .ZN(n_0_678));
   AND2_X1 i_0_123_0 (.A1(n_789), .A2(n_0_672), .ZN(n_0_9));
   OR2_X1 i_0_124_0 (.A1(n_0_672), .A2(n_789), .ZN(n_0_673));
   AND2_X1 i_0_125_0 (.A1(n_791), .A2(n_0_667), .ZN(n_0_10));
   OR2_X1 i_0_126_0 (.A1(n_0_667), .A2(n_791), .ZN(n_0_668));
   AND2_X1 i_0_127_0 (.A1(n_794), .A2(n_0_657), .ZN(n_0_11));
   OR2_X1 i_0_128_0 (.A1(n_0_657), .A2(n_794), .ZN(n_0_658));
   AND2_X1 i_0_129_0 (.A1(n_796), .A2(n_0_651), .ZN(n_0_12));
   OR2_X1 i_0_130_0 (.A1(n_0_651), .A2(n_796), .ZN(n_0_652));
   AND2_X1 i_0_131_0 (.A1(n_798), .A2(n_0_645), .ZN(n_0_13));
   OR2_X1 i_0_132_0 (.A1(n_0_645), .A2(n_798), .ZN(n_0_646));
   AND2_X1 i_0_133_0 (.A1(n_800), .A2(n_0_639), .ZN(n_0_14));
   OR2_X1 i_0_134_0 (.A1(n_0_639), .A2(n_800), .ZN(n_0_640));
   AND2_X1 i_0_135_0 (.A1(n_802), .A2(n_0_633), .ZN(n_0_15));
   OR2_X1 i_0_136_0 (.A1(n_0_633), .A2(n_802), .ZN(n_0_634));
   AND2_X1 i_0_137_0 (.A1(n_804), .A2(n_0_627), .ZN(n_0_16));
   OR2_X1 i_0_138_0 (.A1(n_0_627), .A2(n_804), .ZN(n_0_628));
   AND2_X1 i_0_139_0 (.A1(n_806), .A2(n_0_621), .ZN(n_0_17));
   OR2_X1 i_0_140_0 (.A1(n_0_621), .A2(n_806), .ZN(n_0_622));
   AND2_X1 i_0_141_0 (.A1(n_808), .A2(n_0_615), .ZN(n_0_18));
   OR2_X1 i_0_142_0 (.A1(n_0_615), .A2(n_808), .ZN(n_0_616));
   AND2_X1 i_0_143_0 (.A1(n_810), .A2(n_0_609), .ZN(n_0_19));
   OR2_X1 i_0_144_0 (.A1(n_0_609), .A2(n_810), .ZN(n_0_610));
   AND2_X1 i_0_145_0 (.A1(n_812), .A2(n_0_603), .ZN(n_0_20));
   OR2_X1 i_0_146_0 (.A1(n_0_603), .A2(n_812), .ZN(n_0_604));
   AND2_X1 i_0_147_0 (.A1(n_814), .A2(n_0_597), .ZN(n_0_21));
   OR2_X1 i_0_148_0 (.A1(n_0_597), .A2(n_814), .ZN(n_0_598));
   AND2_X1 i_0_149_0 (.A1(n_816), .A2(n_0_592), .ZN(n_0_22));
   OR2_X1 i_0_150_0 (.A1(n_0_592), .A2(n_816), .ZN(n_0_593));
   AND2_X1 i_0_151_0 (.A1(n_818), .A2(n_0_586), .ZN(n_0_23));
   OR2_X1 i_0_152_0 (.A1(n_0_586), .A2(n_818), .ZN(n_0_587));
   AND2_X1 i_0_153_0 (.A1(n_820), .A2(n_0_580), .ZN(n_0_24));
   OR2_X1 i_0_154_0 (.A1(n_0_580), .A2(n_820), .ZN(n_0_581));
   AND2_X1 i_0_155_0 (.A1(n_822), .A2(n_0_574), .ZN(n_0_25));
   OR2_X1 i_0_156_0 (.A1(n_0_574), .A2(n_822), .ZN(n_0_575));
   AND2_X1 i_0_157_0 (.A1(n_824), .A2(n_0_568), .ZN(n_0_26));
   OR2_X1 i_0_158_0 (.A1(n_0_568), .A2(n_824), .ZN(n_0_569));
   AND2_X1 i_0_159_0 (.A1(n_826), .A2(n_0_562), .ZN(n_0_27));
   OR2_X1 i_0_160_0 (.A1(n_0_562), .A2(n_826), .ZN(n_0_563));
   AND2_X1 i_0_161_0 (.A1(n_828), .A2(n_0_556), .ZN(n_0_28));
   OR2_X1 i_0_162_0 (.A1(n_0_556), .A2(n_828), .ZN(n_0_557));
   AND2_X1 i_0_163_0 (.A1(n_830), .A2(n_0_550), .ZN(n_0_29));
   OR2_X1 i_0_164_0 (.A1(n_0_550), .A2(n_830), .ZN(n_0_551));
   AND2_X1 i_0_165_0 (.A1(n_831), .A2(n_0_545), .ZN(n_0_30));
   OR2_X1 i_0_166_0 (.A1(n_0_545), .A2(n_831), .ZN(n_0_546));
   AND2_X1 i_0_167_0 (.A1(n_679), .A2(n_0_541), .ZN(n_0_31));
   OR2_X1 i_0_168_0 (.A1(n_0_541), .A2(n_679), .ZN(n_0_542));
   AND2_X1 i_0_169_0 (.A1(n_681), .A2(n_0_535), .ZN(n_0_32));
   OR2_X1 i_0_170_0 (.A1(n_0_535), .A2(n_681), .ZN(n_0_536));
   AND2_X1 i_0_171_0 (.A1(n_683), .A2(n_0_529), .ZN(n_0_33));
   OR2_X1 i_0_172_0 (.A1(n_0_529), .A2(n_683), .ZN(n_0_530));
   AND2_X1 i_0_173_0 (.A1(n_685), .A2(n_0_523), .ZN(n_0_34));
   OR2_X1 i_0_174_0 (.A1(n_0_523), .A2(n_685), .ZN(n_0_524));
   AND2_X1 i_0_175_0 (.A1(n_687), .A2(n_0_517), .ZN(n_0_35));
   OR2_X1 i_0_176_0 (.A1(n_0_517), .A2(n_687), .ZN(n_0_518));
   AND2_X1 i_0_177_0 (.A1(n_689), .A2(n_0_511), .ZN(n_0_36));
   OR2_X1 i_0_178_0 (.A1(n_0_511), .A2(n_689), .ZN(n_0_512));
   AND2_X1 i_0_179_0 (.A1(n_691), .A2(n_0_505), .ZN(n_0_37));
   OR2_X1 i_0_180_0 (.A1(n_0_505), .A2(n_691), .ZN(n_0_506));
   AND2_X1 i_0_181_0 (.A1(n_693), .A2(n_0_499), .ZN(n_0_38));
   OR2_X1 i_0_182_0 (.A1(n_0_499), .A2(n_693), .ZN(n_0_500));
   AND2_X1 i_0_183_0 (.A1(n_695), .A2(n_0_493), .ZN(n_0_39));
   OR2_X1 i_0_184_0 (.A1(n_0_493), .A2(n_695), .ZN(n_0_494));
   AND2_X1 i_0_185_0 (.A1(n_697), .A2(n_0_487), .ZN(n_0_40));
   OR2_X1 i_0_186_0 (.A1(n_0_487), .A2(n_697), .ZN(n_0_488));
   AND2_X1 i_0_187_0 (.A1(n_699), .A2(n_0_481), .ZN(n_0_41));
   OR2_X1 i_0_188_0 (.A1(n_0_481), .A2(n_699), .ZN(n_0_482));
   AND2_X1 i_0_189_0 (.A1(n_0_475), .A2(n_701), .ZN(n_0_42));
   OR2_X1 i_0_190_0 (.A1(n_0_475), .A2(n_701), .ZN(n_0_476));
   AND2_X1 i_0_191_0 (.A1(n_703), .A2(n_0_469), .ZN(n_0_43));
   OR2_X1 i_0_192_0 (.A1(n_0_469), .A2(n_703), .ZN(n_0_470));
   AND2_X1 i_0_193_0 (.A1(n_705), .A2(n_0_463), .ZN(n_0_44));
   NAND2_X1 i_0_194_0 (.A1(n_0_194_0), .A2(n_0_194_1), .ZN(n_0_464));
   INV_X1 i_0_194_1 (.A(n_0_463), .ZN(n_0_194_0));
   INV_X1 i_0_194_2 (.A(n_705), .ZN(n_0_194_1));
   AND2_X1 i_0_195_0 (.A1(n_0_457), .A2(n_707), .ZN(n_0_45));
   NAND2_X1 i_0_196_0 (.A1(n_0_196_0), .A2(n_0_196_1), .ZN(n_0_458));
   INV_X1 i_0_196_1 (.A(n_0_457), .ZN(n_0_196_0));
   INV_X1 i_0_196_2 (.A(n_707), .ZN(n_0_196_1));
   AND2_X1 i_0_197_0 (.A1(n_738), .A2(n_0_452), .ZN(n_0_46));
   OR2_X1 i_0_198_0 (.A1(n_0_452), .A2(n_738), .ZN(n_0_453));
   AND2_X1 i_0_199_0 (.A1(n_711), .A2(n_0_449), .ZN(n_0_47));
   OR2_X1 i_0_200_0 (.A1(n_0_449), .A2(n_711), .ZN(n_0_450));
   AND2_X1 i_0_201_0 (.A1(n_713), .A2(n_0_443), .ZN(n_0_48));
   OR2_X1 i_0_202_0 (.A1(n_0_443), .A2(n_713), .ZN(n_0_444));
   AND2_X1 i_0_203_0 (.A1(n_715), .A2(n_0_437), .ZN(n_0_49));
   OR2_X1 i_0_204_0 (.A1(n_0_437), .A2(n_715), .ZN(n_0_438));
   AND2_X1 i_0_205_0 (.A1(n_717), .A2(n_0_432), .ZN(n_0_50));
   OR2_X1 i_0_206_0 (.A1(n_0_432), .A2(n_717), .ZN(n_0_433));
   AND2_X1 i_0_207_0 (.A1(n_719), .A2(n_0_426), .ZN(n_0_51));
   OR2_X1 i_0_208_0 (.A1(n_0_426), .A2(n_719), .ZN(n_0_427));
   AND2_X1 i_0_209_0 (.A1(n_721), .A2(n_0_420), .ZN(n_0_52));
   OR2_X1 i_0_210_0 (.A1(n_0_420), .A2(n_721), .ZN(n_0_421));
   AND2_X1 i_0_211_0 (.A1(n_723), .A2(n_0_414), .ZN(n_0_53));
   OR2_X1 i_0_212_0 (.A1(n_0_414), .A2(n_723), .ZN(n_0_415));
   AND2_X1 i_0_213_0 (.A1(n_726), .A2(n_0_408), .ZN(n_0_54));
   NAND2_X1 i_0_214_0 (.A1(n_0_214_0), .A2(n_0_214_1), .ZN(n_0_409));
   INV_X1 i_0_214_1 (.A(n_0_408), .ZN(n_0_214_0));
   INV_X1 i_0_214_2 (.A(n_726), .ZN(n_0_214_1));
   OR2_X1 i_0_215_0 (.A1(n_0_403), .A2(n_735), .ZN(n_854));
   AND2_X1 i_0_216_0 (.A1(n_775), .A2(n_0_708), .ZN(n_0_55));
   OR2_X1 i_0_217_0 (.A1(n_0_708), .A2(n_775), .ZN(n_0_709));
   AND2_X1 i_0_218_0 (.A1(n_786), .A2(n_0_680), .ZN(n_0_56));
   OR2_X1 i_0_219_0 (.A1(n_0_680), .A2(n_786), .ZN(n_0_681));
   AND2_X1 i_0_220_0 (.A1(n_797), .A2(n_0_648), .ZN(n_0_57));
   OR2_X1 i_0_221_0 (.A1(n_0_648), .A2(n_797), .ZN(n_0_649));
   AND2_X1 i_0_222_0 (.A1(n_801), .A2(n_0_636), .ZN(n_0_58));
   OR2_X1 i_0_223_0 (.A1(n_0_636), .A2(n_801), .ZN(n_0_637));
   AND2_X1 i_0_224_0 (.A1(n_805), .A2(n_0_624), .ZN(n_0_59));
   OR2_X1 i_0_225_0 (.A1(n_0_624), .A2(n_805), .ZN(n_0_625));
   AND2_X1 i_0_226_0 (.A1(n_809), .A2(n_0_612), .ZN(n_0_60));
   OR2_X1 i_0_227_0 (.A1(n_0_612), .A2(n_809), .ZN(n_0_613));
   AND2_X1 i_0_228_0 (.A1(n_813), .A2(n_0_600), .ZN(n_0_61));
   OR2_X1 i_0_229_0 (.A1(n_0_600), .A2(n_813), .ZN(n_0_601));
   AND2_X1 i_0_230_0 (.A1(n_817), .A2(n_0_589), .ZN(n_0_62));
   OR2_X1 i_0_231_0 (.A1(n_0_589), .A2(n_817), .ZN(n_0_590));
   AND2_X1 i_0_232_0 (.A1(n_821), .A2(n_0_577), .ZN(n_0_63));
   OR2_X1 i_0_233_0 (.A1(n_0_577), .A2(n_821), .ZN(n_0_578));
   AND2_X1 i_0_234_0 (.A1(n_825), .A2(n_0_565), .ZN(n_0_64));
   OR2_X1 i_0_235_0 (.A1(n_0_565), .A2(n_825), .ZN(n_0_566));
   AND2_X1 i_0_236_0 (.A1(n_829), .A2(n_0_553), .ZN(n_0_65));
   OR2_X1 i_0_237_0 (.A1(n_0_553), .A2(n_829), .ZN(n_0_554));
   OR2_X1 i_0_238_0 (.A1(n_0_544), .A2(n_678), .ZN(n_855));
   AND2_X1 i_0_239_0 (.A1(n_682), .A2(n_0_532), .ZN(n_0_66));
   OR2_X1 i_0_240_0 (.A1(n_0_532), .A2(n_682), .ZN(n_0_533));
   AND2_X1 i_0_241_0 (.A1(n_686), .A2(n_0_520), .ZN(n_0_67));
   OR2_X1 i_0_242_0 (.A1(n_0_520), .A2(n_686), .ZN(n_0_521));
   AND2_X1 i_0_243_0 (.A1(n_690), .A2(n_0_508), .ZN(n_0_68));
   OR2_X1 i_0_244_0 (.A1(n_0_508), .A2(n_690), .ZN(n_0_509));
   AND2_X1 i_0_245_0 (.A1(n_694), .A2(n_0_496), .ZN(n_0_69));
   OR2_X1 i_0_246_0 (.A1(n_0_496), .A2(n_694), .ZN(n_0_497));
   AND2_X1 i_0_247_0 (.A1(n_698), .A2(n_0_484), .ZN(n_0_70));
   OR2_X1 i_0_248_0 (.A1(n_0_484), .A2(n_698), .ZN(n_0_485));
   AND2_X1 i_0_249_0 (.A1(n_702), .A2(n_0_472), .ZN(n_0_71));
   OR2_X1 i_0_250_0 (.A1(n_0_472), .A2(n_702), .ZN(n_0_473));
   AND2_X1 i_0_251_0 (.A1(n_0_460), .A2(n_706), .ZN(n_0_72));
   NAND2_X1 i_0_252_0 (.A1(n_0_252_0), .A2(n_0_252_1), .ZN(n_0_461));
   INV_X1 i_0_252_1 (.A(n_0_460), .ZN(n_0_252_0));
   INV_X1 i_0_252_2 (.A(n_706), .ZN(n_0_252_1));
   AND2_X1 i_0_253_0 (.A1(n_714), .A2(n_0_440), .ZN(n_0_73));
   OR2_X1 i_0_254_0 (.A1(n_0_440), .A2(n_714), .ZN(n_0_441));
   AND2_X1 i_0_255_0 (.A1(n_718), .A2(n_0_429), .ZN(n_0_74));
   OR2_X1 i_0_256_0 (.A1(n_0_429), .A2(n_718), .ZN(n_0_430));
   AND2_X1 i_0_257_0 (.A1(n_722), .A2(n_0_417), .ZN(n_0_75));
   OR2_X1 i_0_258_0 (.A1(n_0_417), .A2(n_722), .ZN(n_0_418));
   AND2_X1 i_0_259_0 (.A1(n_725), .A2(n_0_411), .ZN(n_0_76));
   OR2_X1 i_0_260_0 (.A1(n_0_411), .A2(n_725), .ZN(n_0_412));
   AND2_X1 i_0_261_0 (.A1(n_729), .A2(n_0_405), .ZN(n_0_77));
   NAND2_X1 i_0_262_0 (.A1(n_0_262_0), .A2(n_0_262_1), .ZN(n_0_406));
   INV_X1 i_0_262_1 (.A(n_0_405), .ZN(n_0_262_0));
   INV_X1 i_0_262_2 (.A(n_729), .ZN(n_0_262_1));
   AND2_X1 i_0_263_0 (.A1(n_732), .A2(n_0_400), .ZN(n_0_78));
   OR2_X1 i_0_264_0 (.A1(n_0_400), .A2(n_732), .ZN(n_0_401));
   AND2_X1 i_0_265_0 (.A1(n_736), .A2(n_0_392), .ZN(n_0_79));
   OR2_X1 i_0_266_0 (.A1(n_0_392), .A2(n_736), .ZN(n_0_393));
   AND2_X1 i_0_267_0 (.A1(n_795), .A2(n_0_654), .ZN(n_0_80));
   OR2_X1 i_0_268_0 (.A1(n_0_654), .A2(n_795), .ZN(n_0_655));
   AND2_X1 i_0_269_0 (.A1(n_803), .A2(n_0_630), .ZN(n_0_81));
   OR2_X1 i_0_270_0 (.A1(n_0_630), .A2(n_803), .ZN(n_0_631));
   AND2_X1 i_0_271_0 (.A1(n_811), .A2(n_0_606), .ZN(n_0_82));
   OR2_X1 i_0_272_0 (.A1(n_0_606), .A2(n_811), .ZN(n_0_607));
   AND2_X1 i_0_273_0 (.A1(n_819), .A2(n_0_583), .ZN(n_0_83));
   OR2_X1 i_0_274_0 (.A1(n_0_583), .A2(n_819), .ZN(n_0_584));
   AND2_X1 i_0_275_0 (.A1(n_827), .A2(n_0_559), .ZN(n_0_84));
   OR2_X1 i_0_276_0 (.A1(n_0_559), .A2(n_827), .ZN(n_0_560));
   AND2_X1 i_0_277_0 (.A1(n_680), .A2(n_0_538), .ZN(n_0_85));
   NAND2_X1 i_0_278_0 (.A1(n_0_278_0), .A2(n_0_278_1), .ZN(n_0_539));
   INV_X1 i_0_278_1 (.A(n_0_538), .ZN(n_0_278_0));
   INV_X1 i_0_278_2 (.A(n_680), .ZN(n_0_278_1));
   AND2_X1 i_0_279_0 (.A1(n_688), .A2(n_0_514), .ZN(n_0_86));
   OR2_X1 i_0_280_0 (.A1(n_0_514), .A2(n_688), .ZN(n_0_515));
   AND2_X1 i_0_281_0 (.A1(n_696), .A2(n_0_490), .ZN(n_0_87));
   OR2_X1 i_0_282_0 (.A1(n_0_490), .A2(n_696), .ZN(n_0_491));
   AND2_X1 i_0_283_0 (.A1(n_704), .A2(n_0_466), .ZN(n_0_88));
   NAND2_X1 i_0_284_0 (.A1(n_0_284_0), .A2(n_0_284_1), .ZN(n_0_467));
   INV_X1 i_0_284_1 (.A(n_0_466), .ZN(n_0_284_0));
   INV_X1 i_0_284_2 (.A(n_704), .ZN(n_0_284_1));
   AND2_X1 i_0_285_0 (.A1(n_712), .A2(n_0_446), .ZN(n_0_89));
   OR2_X1 i_0_286_0 (.A1(n_0_446), .A2(n_712), .ZN(n_0_447));
   AND2_X1 i_0_287_0 (.A1(n_720), .A2(n_0_423), .ZN(n_0_90));
   OR2_X1 i_0_288_0 (.A1(n_0_423), .A2(n_720), .ZN(n_0_424));
   AND2_X1 i_0_289_0 (.A1(n_727), .A2(n_852), .ZN(n_0_91));
   AND2_X1 i_0_290_0 (.A1(n_734), .A2(n_0_397), .ZN(n_0_92));
   OR2_X1 i_0_291_0 (.A1(n_0_397), .A2(n_734), .ZN(n_0_398));
   AND2_X1 i_0_292_0 (.A1(n_792), .A2(n_0_664), .ZN(n_0_93));
   OR2_X1 i_0_293_0 (.A1(n_0_664), .A2(n_792), .ZN(n_0_665));
   AND2_X1 i_0_294_0 (.A1(n_807), .A2(n_0_618), .ZN(n_0_94));
   OR2_X1 i_0_295_0 (.A1(n_0_618), .A2(n_807), .ZN(n_0_619));
   AND2_X1 i_0_296_0 (.A1(n_823), .A2(n_0_571), .ZN(n_0_95));
   OR2_X1 i_0_297_0 (.A1(n_0_571), .A2(n_823), .ZN(n_0_572));
   AND2_X1 i_0_298_0 (.A1(n_684), .A2(n_0_526), .ZN(n_0_96));
   OR2_X1 i_0_299_0 (.A1(n_0_526), .A2(n_684), .ZN(n_0_527));
   AND2_X1 i_0_300_0 (.A1(n_700), .A2(n_0_478), .ZN(n_0_97));
   OR2_X1 i_0_301_0 (.A1(n_0_478), .A2(n_700), .ZN(n_0_479));
   OR2_X1 i_0_302_0 (.A1(n_853), .A2(n_716), .ZN(n_0_435));
   OR2_X1 i_0_303_0 (.A1(n_0_404), .A2(n_731), .ZN(n_856));
   AND2_X1 i_0_304_0 (.A1(n_692), .A2(n_0_502), .ZN(n_0_98));
   NAND2_X1 i_0_305_0 (.A1(n_0_305_0), .A2(n_0_305_1), .ZN(n_0_503));
   INV_X1 i_0_305_1 (.A(n_0_502), .ZN(n_0_305_0));
   INV_X1 i_0_305_2 (.A(n_692), .ZN(n_0_305_1));
   AND2_X1 i_0_306_0 (.A1(n_799), .A2(n_0_642), .ZN(n_0_99));
   OR2_X1 i_0_307_0 (.A1(n_0_642), .A2(n_799), .ZN(n_0_643));
   INV_X1 i_0_308_0 (.A(n_0_1), .ZN(n_0_308_0));
   AOI22_X1 i_0_308_1 (.A1(n_0_308_0), .A2(n_0_120), .B1(in_data[0]), .B2(n_0_1), 
      .ZN(n_0_308_1));
   INV_X1 i_0_308_2 (.A(n_0_308_1), .ZN(n_0_262));
   OAI21_X1 i_0_309_0 (.A(n_0_309_0), .B1(n_0_309_1), .B2(n_0_393), .ZN(n_0_263));
   NAND2_X1 i_0_309_1 (.A1(n_0_393), .A2(in_data[0]), .ZN(n_0_309_0));
   INV_X1 i_0_309_2 (.A(n_1091), .ZN(n_0_309_1));
   INV_X1 i_0_310_0 (.A(n_0_310_0), .ZN(n_0_264));
   OAI21_X1 i_0_310_1 (.A(n_0_310_1), .B1(n_0_119), .B2(n_0_395), .ZN(n_0_310_0));
   NAND2_X1 i_0_310_2 (.A1(n_0_395), .A2(n_0_310_2), .ZN(n_0_310_1));
   INV_X1 i_0_310_3 (.A(in_data[0]), .ZN(n_0_310_2));
   INV_X1 i_0_311_0 (.A(n_0_311_0), .ZN(n_0_265));
   OAI21_X1 i_0_311_1 (.A(n_0_311_1), .B1(n_1092), .B2(n_0_398), .ZN(n_0_311_0));
   NAND2_X1 i_0_311_2 (.A1(n_0_398), .A2(n_0_311_2), .ZN(n_0_311_1));
   INV_X1 i_0_311_3 (.A(in_data[0]), .ZN(n_0_311_2));
   INV_X1 i_0_312_0 (.A(n_0_312_0), .ZN(n_0_266));
   OAI21_X1 i_0_312_1 (.A(n_0_312_1), .B1(n_1093), .B2(n_0_401), .ZN(n_0_312_0));
   NAND2_X1 i_0_312_2 (.A1(n_0_401), .A2(n_0_312_2), .ZN(n_0_312_1));
   INV_X1 i_0_312_3 (.A(in_data[0]), .ZN(n_0_312_2));
   INV_X1 i_0_313_0 (.A(n_0_313_0), .ZN(n_0_267));
   OAI21_X1 i_0_313_1 (.A(n_0_313_1), .B1(n_1094), .B2(n_854), .ZN(n_0_313_0));
   NAND2_X1 i_0_313_2 (.A1(n_854), .A2(n_0_313_2), .ZN(n_0_313_1));
   INV_X1 i_0_313_3 (.A(in_data[0]), .ZN(n_0_313_2));
   INV_X1 i_0_314_0 (.A(n_0_314_0), .ZN(n_0_268));
   OAI21_X1 i_0_314_1 (.A(n_0_314_1), .B1(n_1095), .B2(n_856), .ZN(n_0_314_0));
   NAND2_X1 i_0_314_2 (.A1(n_856), .A2(n_0_314_2), .ZN(n_0_314_1));
   INV_X1 i_0_314_3 (.A(in_data[0]), .ZN(n_0_314_2));
   OAI21_X1 i_0_315_0 (.A(n_0_315_0), .B1(n_0_315_1), .B2(n_0_406), .ZN(n_0_269));
   NAND2_X1 i_0_315_1 (.A1(n_0_406), .A2(in_data[0]), .ZN(n_0_315_0));
   INV_X1 i_0_315_2 (.A(n_1096), .ZN(n_0_315_1));
   OAI21_X1 i_0_316_0 (.A(n_0_316_0), .B1(n_0_316_1), .B2(n_0_409), .ZN(n_0_270));
   NAND2_X1 i_0_316_1 (.A1(n_0_409), .A2(in_data[0]), .ZN(n_0_316_0));
   INV_X1 i_0_316_2 (.A(n_1097), .ZN(n_0_316_1));
   INV_X1 i_0_317_0 (.A(n_0_317_0), .ZN(n_0_271));
   OAI21_X1 i_0_317_1 (.A(n_0_317_1), .B1(n_0_895), .B2(n_0_412), .ZN(n_0_317_0));
   NAND2_X1 i_0_317_2 (.A1(n_0_412), .A2(n_0_317_2), .ZN(n_0_317_1));
   INV_X1 i_0_317_3 (.A(in_data[0]), .ZN(n_0_317_2));
   INV_X1 i_0_318_0 (.A(n_0_318_0), .ZN(n_0_272));
   OAI21_X1 i_0_318_1 (.A(n_0_318_1), .B1(n_1189), .B2(n_0_415), .ZN(n_0_318_0));
   NAND2_X1 i_0_318_2 (.A1(n_0_415), .A2(n_0_318_2), .ZN(n_0_318_1));
   INV_X1 i_0_318_3 (.A(in_data[0]), .ZN(n_0_318_2));
   INV_X1 i_0_319_0 (.A(n_0_319_0), .ZN(n_0_273));
   OAI21_X1 i_0_319_1 (.A(n_0_319_1), .B1(n_1098), .B2(n_0_418), .ZN(n_0_319_0));
   NAND2_X1 i_0_319_2 (.A1(n_0_418), .A2(n_0_319_2), .ZN(n_0_319_1));
   INV_X1 i_0_319_3 (.A(in_data[0]), .ZN(n_0_319_2));
   INV_X1 i_0_320_0 (.A(n_0_320_0), .ZN(n_0_274));
   OAI21_X1 i_0_320_1 (.A(n_0_320_1), .B1(n_1099), .B2(n_0_421), .ZN(n_0_320_0));
   NAND2_X1 i_0_320_2 (.A1(n_0_421), .A2(n_0_320_2), .ZN(n_0_320_1));
   INV_X1 i_0_320_3 (.A(in_data[0]), .ZN(n_0_320_2));
   INV_X1 i_0_321_0 (.A(n_0_321_0), .ZN(n_0_275));
   OAI21_X1 i_0_321_1 (.A(n_0_321_1), .B1(n_1100), .B2(n_0_424), .ZN(n_0_321_0));
   NAND2_X1 i_0_321_2 (.A1(n_0_424), .A2(n_0_321_2), .ZN(n_0_321_1));
   INV_X1 i_0_321_3 (.A(in_data[0]), .ZN(n_0_321_2));
   INV_X1 i_0_322_0 (.A(n_0_322_0), .ZN(n_0_276));
   OAI21_X1 i_0_322_1 (.A(n_0_322_1), .B1(n_1101), .B2(n_0_427), .ZN(n_0_322_0));
   NAND2_X1 i_0_322_2 (.A1(n_0_427), .A2(n_0_322_2), .ZN(n_0_322_1));
   INV_X1 i_0_322_3 (.A(in_data[0]), .ZN(n_0_322_2));
   INV_X1 i_0_323_0 (.A(n_0_323_0), .ZN(n_0_277));
   OAI21_X1 i_0_323_1 (.A(n_0_323_1), .B1(n_1102), .B2(n_0_430), .ZN(n_0_323_0));
   NAND2_X1 i_0_323_2 (.A1(n_0_430), .A2(n_0_323_2), .ZN(n_0_323_1));
   INV_X1 i_0_323_3 (.A(in_data[0]), .ZN(n_0_323_2));
   INV_X1 i_0_324_0 (.A(n_0_324_0), .ZN(n_0_278));
   OAI21_X1 i_0_324_1 (.A(n_0_324_1), .B1(n_1103), .B2(n_0_433), .ZN(n_0_324_0));
   NAND2_X1 i_0_324_2 (.A1(n_0_433), .A2(n_0_324_2), .ZN(n_0_324_1));
   INV_X1 i_0_324_3 (.A(in_data[0]), .ZN(n_0_324_2));
   INV_X1 i_0_325_0 (.A(n_0_325_0), .ZN(n_0_279));
   OAI21_X1 i_0_325_1 (.A(n_0_325_1), .B1(n_1188), .B2(n_0_435), .ZN(n_0_325_0));
   NAND2_X1 i_0_325_2 (.A1(n_0_435), .A2(n_0_325_2), .ZN(n_0_325_1));
   INV_X1 i_0_325_3 (.A(in_data[0]), .ZN(n_0_325_2));
   OAI21_X1 i_0_326_0 (.A(n_0_326_0), .B1(n_0_326_1), .B2(n_0_438), .ZN(n_0_280));
   NAND2_X1 i_0_326_1 (.A1(n_0_438), .A2(in_data[0]), .ZN(n_0_326_0));
   INV_X1 i_0_326_2 (.A(n_1104), .ZN(n_0_326_1));
   INV_X1 i_0_327_0 (.A(n_0_327_0), .ZN(n_0_281));
   OAI21_X1 i_0_327_1 (.A(n_0_327_1), .B1(n_1187), .B2(n_0_441), .ZN(n_0_327_0));
   NAND2_X1 i_0_327_2 (.A1(n_0_441), .A2(n_0_327_2), .ZN(n_0_327_1));
   INV_X1 i_0_327_3 (.A(in_data[0]), .ZN(n_0_327_2));
   INV_X1 i_0_328_0 (.A(n_0_328_0), .ZN(n_0_282));
   OAI21_X1 i_0_328_1 (.A(n_0_328_1), .B1(n_1105), .B2(n_0_444), .ZN(n_0_328_0));
   NAND2_X1 i_0_328_2 (.A1(n_0_444), .A2(n_0_328_2), .ZN(n_0_328_1));
   INV_X1 i_0_328_3 (.A(in_data[0]), .ZN(n_0_328_2));
   OAI21_X1 i_0_329_0 (.A(n_0_329_0), .B1(n_0_329_1), .B2(n_0_447), .ZN(n_0_283));
   NAND2_X1 i_0_329_1 (.A1(n_0_447), .A2(in_data[0]), .ZN(n_0_329_0));
   INV_X1 i_0_329_2 (.A(n_0_896), .ZN(n_0_329_1));
   INV_X1 i_0_330_0 (.A(n_0_330_0), .ZN(n_0_284));
   OAI21_X1 i_0_330_1 (.A(n_0_330_1), .B1(n_1186), .B2(n_0_450), .ZN(n_0_330_0));
   NAND2_X1 i_0_330_2 (.A1(n_0_450), .A2(n_0_330_2), .ZN(n_0_330_1));
   INV_X1 i_0_330_3 (.A(in_data[0]), .ZN(n_0_330_2));
   INV_X1 i_0_331_0 (.A(n_0_331_0), .ZN(n_0_285));
   OAI21_X1 i_0_331_1 (.A(n_0_331_1), .B1(n_1106), .B2(n_0_453), .ZN(n_0_331_0));
   NAND2_X1 i_0_331_2 (.A1(n_0_453), .A2(n_0_331_2), .ZN(n_0_331_1));
   INV_X1 i_0_331_3 (.A(in_data[0]), .ZN(n_0_331_2));
   INV_X1 i_0_332_0 (.A(n_0_332_0), .ZN(n_0_286));
   OAI21_X1 i_0_332_1 (.A(n_0_332_1), .B1(n_1107), .B2(n_708), .ZN(n_0_332_0));
   NAND2_X1 i_0_332_2 (.A1(n_708), .A2(n_0_332_2), .ZN(n_0_332_1));
   INV_X1 i_0_332_3 (.A(in_data[0]), .ZN(n_0_332_2));
   OAI21_X1 i_0_333_0 (.A(n_0_333_0), .B1(n_0_333_1), .B2(n_0_458), .ZN(n_0_287));
   NAND2_X1 i_0_333_1 (.A1(n_0_458), .A2(in_data[0]), .ZN(n_0_333_0));
   INV_X1 i_0_333_2 (.A(n_1108), .ZN(n_0_333_1));
   OAI21_X1 i_0_334_0 (.A(n_0_334_0), .B1(n_0_334_1), .B2(n_0_461), .ZN(n_0_288));
   NAND2_X1 i_0_334_1 (.A1(n_0_461), .A2(in_data[0]), .ZN(n_0_334_0));
   INV_X1 i_0_334_2 (.A(n_1109), .ZN(n_0_334_1));
   OAI21_X1 i_0_335_0 (.A(n_0_335_0), .B1(n_0_335_1), .B2(n_0_464), .ZN(n_0_289));
   NAND2_X1 i_0_335_1 (.A1(n_0_464), .A2(in_data[0]), .ZN(n_0_335_0));
   INV_X1 i_0_335_2 (.A(n_0_124), .ZN(n_0_335_1));
   OAI21_X1 i_0_336_0 (.A(n_0_336_0), .B1(n_0_336_1), .B2(n_0_467), .ZN(n_0_290));
   NAND2_X1 i_0_336_1 (.A1(n_0_467), .A2(in_data[0]), .ZN(n_0_336_0));
   INV_X1 i_0_336_2 (.A(n_0_123), .ZN(n_0_336_1));
   INV_X1 i_0_337_0 (.A(n_0_337_0), .ZN(n_0_291));
   OAI21_X1 i_0_337_1 (.A(n_0_337_1), .B1(n_1185), .B2(n_0_470), .ZN(n_0_337_0));
   NAND2_X1 i_0_337_2 (.A1(n_0_470), .A2(n_0_337_2), .ZN(n_0_337_1));
   INV_X1 i_0_337_3 (.A(in_data[0]), .ZN(n_0_337_2));
   INV_X1 i_0_338_0 (.A(n_0_338_0), .ZN(n_0_292));
   OAI21_X1 i_0_338_1 (.A(n_0_338_1), .B1(n_1110), .B2(n_0_473), .ZN(n_0_338_0));
   NAND2_X1 i_0_338_2 (.A1(n_0_473), .A2(n_0_338_2), .ZN(n_0_338_1));
   INV_X1 i_0_338_3 (.A(in_data[0]), .ZN(n_0_338_2));
   OAI21_X1 i_0_339_0 (.A(n_0_339_0), .B1(n_0_339_1), .B2(n_0_476), .ZN(n_0_293));
   NAND2_X1 i_0_339_1 (.A1(n_0_476), .A2(in_data[0]), .ZN(n_0_339_0));
   INV_X1 i_0_339_2 (.A(n_0_100), .ZN(n_0_339_1));
   INV_X1 i_0_340_0 (.A(n_0_479), .ZN(n_0_340_0));
   AOI22_X1 i_0_340_1 (.A1(n_0_340_0), .A2(n_1184), .B1(in_data[0]), .B2(n_0_479), 
      .ZN(n_0_340_1));
   INV_X1 i_0_340_2 (.A(n_0_340_1), .ZN(n_0_294));
   INV_X1 i_0_341_0 (.A(n_0_482), .ZN(n_0_341_0));
   AOI22_X1 i_0_341_1 (.A1(n_0_341_0), .A2(n_1111), .B1(in_data[0]), .B2(n_0_482), 
      .ZN(n_0_341_1));
   INV_X1 i_0_341_2 (.A(n_0_341_1), .ZN(n_0_295));
   INV_X1 i_0_342_0 (.A(n_0_485), .ZN(n_0_342_0));
   AOI22_X1 i_0_342_1 (.A1(n_0_342_0), .A2(n_1112), .B1(in_data[0]), .B2(n_0_485), 
      .ZN(n_0_342_1));
   INV_X1 i_0_342_2 (.A(n_0_342_1), .ZN(n_0_296));
   INV_X1 i_0_343_0 (.A(n_0_488), .ZN(n_0_343_0));
   AOI22_X1 i_0_343_1 (.A1(n_0_343_0), .A2(n_1113), .B1(in_data[0]), .B2(n_0_488), 
      .ZN(n_0_343_1));
   INV_X1 i_0_343_2 (.A(n_0_343_1), .ZN(n_0_297));
   INV_X1 i_0_344_0 (.A(n_0_344_0), .ZN(n_0_298));
   OAI21_X1 i_0_344_1 (.A(n_0_344_1), .B1(n_1183), .B2(n_0_491), .ZN(n_0_344_0));
   NAND2_X1 i_0_344_2 (.A1(n_0_491), .A2(n_0_344_2), .ZN(n_0_344_1));
   INV_X1 i_0_344_3 (.A(in_data[0]), .ZN(n_0_344_2));
   INV_X1 i_0_345_0 (.A(n_0_494), .ZN(n_0_345_0));
   AOI22_X1 i_0_345_1 (.A1(n_0_345_0), .A2(n_1182), .B1(in_data[0]), .B2(n_0_494), 
      .ZN(n_0_345_1));
   INV_X1 i_0_345_2 (.A(n_0_345_1), .ZN(n_0_299));
   INV_X1 i_0_346_0 (.A(n_0_497), .ZN(n_0_346_0));
   AOI22_X1 i_0_346_1 (.A1(n_0_346_0), .A2(n_1181), .B1(in_data[0]), .B2(n_0_497), 
      .ZN(n_0_346_1));
   INV_X1 i_0_346_2 (.A(n_0_346_1), .ZN(n_0_300));
   INV_X1 i_0_347_0 (.A(n_0_500), .ZN(n_0_347_0));
   AOI22_X1 i_0_347_1 (.A1(n_0_347_0), .A2(n_1180), .B1(in_data[0]), .B2(n_0_500), 
      .ZN(n_0_347_1));
   INV_X1 i_0_347_2 (.A(n_0_347_1), .ZN(n_0_301));
   OAI21_X1 i_0_348_0 (.A(n_0_348_0), .B1(n_0_348_1), .B2(n_0_503), .ZN(n_0_302));
   NAND2_X1 i_0_348_1 (.A1(n_0_503), .A2(in_data[0]), .ZN(n_0_348_0));
   INV_X1 i_0_348_2 (.A(n_0_897), .ZN(n_0_348_1));
   INV_X1 i_0_349_0 (.A(n_0_349_0), .ZN(n_0_303));
   OAI21_X1 i_0_349_1 (.A(n_0_349_1), .B1(n_0_101), .B2(n_0_506), .ZN(n_0_349_0));
   NAND2_X1 i_0_349_2 (.A1(n_0_506), .A2(n_0_349_2), .ZN(n_0_349_1));
   INV_X1 i_0_349_3 (.A(in_data[0]), .ZN(n_0_349_2));
   INV_X1 i_0_350_0 (.A(n_0_350_0), .ZN(n_0_304));
   OAI21_X1 i_0_350_1 (.A(n_0_350_1), .B1(n_1114), .B2(n_0_509), .ZN(n_0_350_0));
   NAND2_X1 i_0_350_2 (.A1(n_0_509), .A2(n_0_350_2), .ZN(n_0_350_1));
   INV_X1 i_0_350_3 (.A(in_data[0]), .ZN(n_0_350_2));
   INV_X1 i_0_351_0 (.A(n_0_351_0), .ZN(n_0_305));
   OAI21_X1 i_0_351_1 (.A(n_0_351_1), .B1(n_1115), .B2(n_0_512), .ZN(n_0_351_0));
   NAND2_X1 i_0_351_2 (.A1(n_0_512), .A2(n_0_351_2), .ZN(n_0_351_1));
   INV_X1 i_0_351_3 (.A(in_data[0]), .ZN(n_0_351_2));
   INV_X1 i_0_352_0 (.A(n_0_515), .ZN(n_0_352_0));
   AOI22_X1 i_0_352_1 (.A1(n_0_352_0), .A2(n_1116), .B1(in_data[0]), .B2(n_0_515), 
      .ZN(n_0_352_1));
   INV_X1 i_0_352_2 (.A(n_0_352_1), .ZN(n_0_306));
   INV_X1 i_0_353_0 (.A(n_0_518), .ZN(n_0_353_0));
   AOI22_X1 i_0_353_1 (.A1(n_0_353_0), .A2(n_1117), .B1(in_data[0]), .B2(n_0_518), 
      .ZN(n_0_353_1));
   INV_X1 i_0_353_2 (.A(n_0_353_1), .ZN(n_0_307));
   INV_X1 i_0_354_0 (.A(n_0_354_0), .ZN(n_0_308));
   OAI21_X1 i_0_354_1 (.A(n_0_354_1), .B1(n_1118), .B2(n_0_521), .ZN(n_0_354_0));
   NAND2_X1 i_0_354_2 (.A1(n_0_521), .A2(n_0_354_2), .ZN(n_0_354_1));
   INV_X1 i_0_354_3 (.A(in_data[0]), .ZN(n_0_354_2));
   INV_X1 i_0_355_0 (.A(n_0_524), .ZN(n_0_355_0));
   AOI22_X1 i_0_355_1 (.A1(n_0_355_0), .A2(n_1119), .B1(in_data[0]), .B2(n_0_524), 
      .ZN(n_0_355_1));
   INV_X1 i_0_355_2 (.A(n_0_355_1), .ZN(n_0_309));
   INV_X1 i_0_356_0 (.A(n_0_527), .ZN(n_0_356_0));
   AOI22_X1 i_0_356_1 (.A1(n_0_356_0), .A2(n_1120), .B1(in_data[0]), .B2(n_0_527), 
      .ZN(n_0_356_1));
   INV_X1 i_0_356_2 (.A(n_0_356_1), .ZN(n_0_310));
   INV_X1 i_0_357_0 (.A(n_0_357_0), .ZN(n_0_311));
   OAI21_X1 i_0_357_1 (.A(n_0_357_1), .B1(n_1121), .B2(n_0_530), .ZN(n_0_357_0));
   NAND2_X1 i_0_357_2 (.A1(n_0_530), .A2(n_0_357_2), .ZN(n_0_357_1));
   INV_X1 i_0_357_3 (.A(in_data[0]), .ZN(n_0_357_2));
   INV_X1 i_0_358_0 (.A(n_0_533), .ZN(n_0_358_0));
   AOI22_X1 i_0_358_1 (.A1(n_0_358_0), .A2(n_1122), .B1(in_data[0]), .B2(n_0_533), 
      .ZN(n_0_358_1));
   INV_X1 i_0_358_2 (.A(n_0_358_1), .ZN(n_0_312));
   INV_X1 i_0_359_0 (.A(n_0_359_0), .ZN(n_0_313));
   OAI21_X1 i_0_359_1 (.A(n_0_359_1), .B1(n_1123), .B2(n_0_536), .ZN(n_0_359_0));
   NAND2_X1 i_0_359_2 (.A1(n_0_536), .A2(n_0_359_2), .ZN(n_0_359_1));
   INV_X1 i_0_359_3 (.A(in_data[0]), .ZN(n_0_359_2));
   OAI21_X1 i_0_360_0 (.A(n_0_360_0), .B1(n_0_360_1), .B2(n_0_539), .ZN(n_0_314));
   NAND2_X1 i_0_360_1 (.A1(n_0_539), .A2(in_data[0]), .ZN(n_0_360_0));
   INV_X1 i_0_360_2 (.A(n_0_122), .ZN(n_0_360_1));
   INV_X1 i_0_361_0 (.A(n_0_361_0), .ZN(n_0_315));
   OAI21_X1 i_0_361_1 (.A(n_0_361_1), .B1(n_1124), .B2(n_0_542), .ZN(n_0_361_0));
   NAND2_X1 i_0_361_2 (.A1(n_0_542), .A2(n_0_361_2), .ZN(n_0_361_1));
   INV_X1 i_0_361_3 (.A(in_data[0]), .ZN(n_0_361_2));
   INV_X1 i_0_362_0 (.A(n_0_362_0), .ZN(n_0_316));
   OAI21_X1 i_0_362_1 (.A(n_0_362_1), .B1(n_1125), .B2(n_855), .ZN(n_0_362_0));
   NAND2_X1 i_0_362_2 (.A1(n_855), .A2(n_0_362_2), .ZN(n_0_362_1));
   INV_X1 i_0_362_3 (.A(in_data[0]), .ZN(n_0_362_2));
   INV_X1 i_0_363_0 (.A(n_0_363_0), .ZN(n_0_317));
   OAI21_X1 i_0_363_1 (.A(n_0_363_1), .B1(n_1179), .B2(n_0_546), .ZN(n_0_363_0));
   NAND2_X1 i_0_363_2 (.A1(n_0_546), .A2(n_0_363_2), .ZN(n_0_363_1));
   INV_X1 i_0_363_3 (.A(in_data[0]), .ZN(n_0_363_2));
   INV_X1 i_0_364_0 (.A(n_0_364_0), .ZN(n_0_318));
   OAI21_X1 i_0_364_1 (.A(n_0_364_1), .B1(n_0_120), .B2(n_837), .ZN(n_0_364_0));
   NAND2_X1 i_0_364_2 (.A1(n_837), .A2(n_0_364_2), .ZN(n_0_364_1));
   INV_X1 i_0_364_3 (.A(in_data[0]), .ZN(n_0_364_2));
   INV_X1 i_0_365_0 (.A(n_0_551), .ZN(n_0_365_0));
   AOI22_X1 i_0_365_1 (.A1(n_0_365_0), .A2(n_1126), .B1(in_data[0]), .B2(n_0_551), 
      .ZN(n_0_365_1));
   INV_X1 i_0_365_2 (.A(n_0_365_1), .ZN(n_0_319));
   INV_X1 i_0_366_0 (.A(n_0_366_0), .ZN(n_0_320));
   OAI21_X1 i_0_366_1 (.A(n_0_366_1), .B1(n_1127), .B2(n_0_554), .ZN(n_0_366_0));
   NAND2_X1 i_0_366_2 (.A1(n_0_554), .A2(n_0_366_2), .ZN(n_0_366_1));
   INV_X1 i_0_366_3 (.A(in_data[0]), .ZN(n_0_366_2));
   INV_X1 i_0_367_0 (.A(n_0_557), .ZN(n_0_367_0));
   AOI22_X1 i_0_367_1 (.A1(n_0_367_0), .A2(n_1128), .B1(in_data[0]), .B2(n_0_557), 
      .ZN(n_0_367_1));
   INV_X1 i_0_367_2 (.A(n_0_367_1), .ZN(n_0_321));
   INV_X1 i_0_368_0 (.A(n_0_368_0), .ZN(n_0_322));
   OAI21_X1 i_0_368_1 (.A(n_0_368_1), .B1(n_1178), .B2(n_0_560), .ZN(n_0_368_0));
   NAND2_X1 i_0_368_2 (.A1(n_0_560), .A2(n_0_368_2), .ZN(n_0_368_1));
   INV_X1 i_0_368_3 (.A(in_data[0]), .ZN(n_0_368_2));
   INV_X1 i_0_369_0 (.A(n_0_563), .ZN(n_0_369_0));
   AOI22_X1 i_0_369_1 (.A1(n_0_369_0), .A2(n_1129), .B1(in_data[0]), .B2(n_0_563), 
      .ZN(n_0_369_1));
   INV_X1 i_0_369_2 (.A(n_0_369_1), .ZN(n_0_323));
   INV_X1 i_0_370_0 (.A(n_0_566), .ZN(n_0_370_0));
   AOI22_X1 i_0_370_1 (.A1(n_0_370_0), .A2(n_1130), .B1(in_data[0]), .B2(n_0_566), 
      .ZN(n_0_370_1));
   INV_X1 i_0_370_2 (.A(n_0_370_1), .ZN(n_0_324));
   INV_X1 i_0_371_0 (.A(n_0_569), .ZN(n_0_371_0));
   AOI22_X1 i_0_371_1 (.A1(n_0_371_0), .A2(n_1131), .B1(in_data[0]), .B2(n_0_569), 
      .ZN(n_0_371_1));
   INV_X1 i_0_371_2 (.A(n_0_371_1), .ZN(n_0_325));
   INV_X1 i_0_372_0 (.A(n_0_572), .ZN(n_0_372_0));
   AOI22_X1 i_0_372_1 (.A1(n_0_372_0), .A2(n_1132), .B1(in_data[0]), .B2(n_0_572), 
      .ZN(n_0_372_1));
   INV_X1 i_0_372_2 (.A(n_0_372_1), .ZN(n_0_326));
   INV_X1 i_0_373_0 (.A(n_0_575), .ZN(n_0_373_0));
   AOI22_X1 i_0_373_1 (.A1(n_0_373_0), .A2(n_1133), .B1(in_data[0]), .B2(n_0_575), 
      .ZN(n_0_373_1));
   INV_X1 i_0_373_2 (.A(n_0_373_1), .ZN(n_0_327));
   INV_X1 i_0_374_0 (.A(n_0_578), .ZN(n_0_374_0));
   AOI22_X1 i_0_374_1 (.A1(n_0_374_0), .A2(n_1134), .B1(in_data[0]), .B2(n_0_578), 
      .ZN(n_0_374_1));
   INV_X1 i_0_374_2 (.A(n_0_374_1), .ZN(n_0_328));
   INV_X1 i_0_375_0 (.A(n_0_581), .ZN(n_0_375_0));
   AOI22_X1 i_0_375_1 (.A1(n_0_375_0), .A2(n_1135), .B1(in_data[0]), .B2(n_0_581), 
      .ZN(n_0_375_1));
   INV_X1 i_0_375_2 (.A(n_0_375_1), .ZN(n_0_329));
   INV_X1 i_0_376_0 (.A(n_0_376_0), .ZN(n_0_330));
   OAI21_X1 i_0_376_1 (.A(n_0_376_1), .B1(n_1177), .B2(n_0_584), .ZN(n_0_376_0));
   NAND2_X1 i_0_376_2 (.A1(n_0_584), .A2(n_0_376_2), .ZN(n_0_376_1));
   INV_X1 i_0_376_3 (.A(in_data[0]), .ZN(n_0_376_2));
   INV_X1 i_0_377_0 (.A(n_0_587), .ZN(n_0_377_0));
   AOI22_X1 i_0_377_1 (.A1(n_0_377_0), .A2(n_1136), .B1(in_data[0]), .B2(n_0_587), 
      .ZN(n_0_377_1));
   INV_X1 i_0_377_2 (.A(n_0_377_1), .ZN(n_0_331));
   INV_X1 i_0_378_0 (.A(n_0_378_0), .ZN(n_0_332));
   OAI21_X1 i_0_378_1 (.A(n_0_378_1), .B1(n_1137), .B2(n_0_590), .ZN(n_0_378_0));
   NAND2_X1 i_0_378_2 (.A1(n_0_590), .A2(n_0_378_2), .ZN(n_0_378_1));
   INV_X1 i_0_378_3 (.A(in_data[0]), .ZN(n_0_378_2));
   INV_X1 i_0_379_0 (.A(n_0_379_0), .ZN(n_0_333));
   OAI21_X1 i_0_379_1 (.A(n_0_379_1), .B1(n_1138), .B2(n_0_593), .ZN(n_0_379_0));
   NAND2_X1 i_0_379_2 (.A1(n_0_593), .A2(n_0_379_2), .ZN(n_0_379_1));
   INV_X1 i_0_379_3 (.A(in_data[0]), .ZN(n_0_379_2));
   OAI21_X1 i_0_380_0 (.A(n_0_380_0), .B1(n_0_380_1), .B2(n_677), .ZN(n_0_334));
   NAND2_X1 i_0_380_1 (.A1(n_677), .A2(in_data[0]), .ZN(n_0_380_0));
   INV_X1 i_0_380_2 (.A(n_1139), .ZN(n_0_380_1));
   INV_X1 i_0_381_0 (.A(n_0_381_0), .ZN(n_0_335));
   OAI21_X1 i_0_381_1 (.A(n_0_381_1), .B1(n_1140), .B2(n_0_598), .ZN(n_0_381_0));
   NAND2_X1 i_0_381_2 (.A1(n_0_598), .A2(n_0_381_2), .ZN(n_0_381_1));
   INV_X1 i_0_381_3 (.A(in_data[0]), .ZN(n_0_381_2));
   INV_X1 i_0_382_0 (.A(n_0_601), .ZN(n_0_382_0));
   AOI22_X1 i_0_382_1 (.A1(n_0_382_0), .A2(n_1141), .B1(in_data[0]), .B2(n_0_601), 
      .ZN(n_0_382_1));
   INV_X1 i_0_382_2 (.A(n_0_382_1), .ZN(n_0_336));
   INV_X1 i_0_383_0 (.A(n_0_383_0), .ZN(n_0_337));
   OAI21_X1 i_0_383_1 (.A(n_0_383_1), .B1(n_1142), .B2(n_0_604), .ZN(n_0_383_0));
   NAND2_X1 i_0_383_2 (.A1(n_0_604), .A2(n_0_383_2), .ZN(n_0_383_1));
   INV_X1 i_0_383_3 (.A(in_data[0]), .ZN(n_0_383_2));
   INV_X1 i_0_384_0 (.A(n_0_384_0), .ZN(n_0_338));
   OAI21_X1 i_0_384_1 (.A(n_0_384_1), .B1(n_1143), .B2(n_0_607), .ZN(n_0_384_0));
   NAND2_X1 i_0_384_2 (.A1(n_0_607), .A2(n_0_384_2), .ZN(n_0_384_1));
   INV_X1 i_0_384_3 (.A(in_data[0]), .ZN(n_0_384_2));
   INV_X1 i_0_385_0 (.A(n_0_385_0), .ZN(n_0_339));
   OAI21_X1 i_0_385_1 (.A(n_0_385_1), .B1(n_1144), .B2(n_0_610), .ZN(n_0_385_0));
   NAND2_X1 i_0_385_2 (.A1(n_0_610), .A2(n_0_385_2), .ZN(n_0_385_1));
   INV_X1 i_0_385_3 (.A(in_data[0]), .ZN(n_0_385_2));
   INV_X1 i_0_386_0 (.A(n_0_613), .ZN(n_0_386_0));
   AOI22_X1 i_0_386_1 (.A1(n_0_386_0), .A2(n_1145), .B1(in_data[0]), .B2(n_0_613), 
      .ZN(n_0_386_1));
   INV_X1 i_0_386_2 (.A(n_0_386_1), .ZN(n_0_340));
   INV_X1 i_0_387_0 (.A(n_0_387_0), .ZN(n_0_341));
   OAI21_X1 i_0_387_1 (.A(n_0_387_1), .B1(n_1146), .B2(n_0_616), .ZN(n_0_387_0));
   NAND2_X1 i_0_387_2 (.A1(n_0_616), .A2(n_0_387_2), .ZN(n_0_387_1));
   INV_X1 i_0_387_3 (.A(in_data[0]), .ZN(n_0_387_2));
   INV_X1 i_0_388_0 (.A(n_0_619), .ZN(n_0_388_0));
   AOI22_X1 i_0_388_1 (.A1(n_0_388_0), .A2(n_1147), .B1(in_data[0]), .B2(n_0_619), 
      .ZN(n_0_388_1));
   INV_X1 i_0_388_2 (.A(n_0_388_1), .ZN(n_0_342));
   INV_X1 i_0_389_0 (.A(n_0_389_0), .ZN(n_0_343));
   OAI21_X1 i_0_389_1 (.A(n_0_389_1), .B1(n_1148), .B2(n_0_622), .ZN(n_0_389_0));
   NAND2_X1 i_0_389_2 (.A1(n_0_622), .A2(n_0_389_2), .ZN(n_0_389_1));
   INV_X1 i_0_389_3 (.A(in_data[0]), .ZN(n_0_389_2));
   INV_X1 i_0_390_0 (.A(n_0_390_0), .ZN(n_0_344));
   OAI21_X1 i_0_390_1 (.A(n_0_390_1), .B1(n_1176), .B2(n_0_625), .ZN(n_0_390_0));
   NAND2_X1 i_0_390_2 (.A1(n_0_625), .A2(n_0_390_2), .ZN(n_0_390_1));
   INV_X1 i_0_390_3 (.A(in_data[0]), .ZN(n_0_390_2));
   OAI21_X1 i_0_391_0 (.A(n_0_391_0), .B1(n_0_391_1), .B2(n_0_628), .ZN(n_0_345));
   NAND2_X1 i_0_391_1 (.A1(n_0_628), .A2(in_data[0]), .ZN(n_0_391_0));
   INV_X1 i_0_391_2 (.A(n_0_898), .ZN(n_0_391_1));
   INV_X1 i_0_392_0 (.A(n_0_392_0), .ZN(n_0_346));
   OAI21_X1 i_0_392_1 (.A(n_0_392_1), .B1(n_1149), .B2(n_0_631), .ZN(n_0_392_0));
   NAND2_X1 i_0_392_2 (.A1(n_0_631), .A2(n_0_392_2), .ZN(n_0_392_1));
   INV_X1 i_0_392_3 (.A(in_data[0]), .ZN(n_0_392_2));
   INV_X1 i_0_393_0 (.A(n_0_393_0), .ZN(n_0_347));
   OAI21_X1 i_0_393_1 (.A(n_0_393_1), .B1(n_1175), .B2(n_0_634), .ZN(n_0_393_0));
   NAND2_X1 i_0_393_2 (.A1(n_0_634), .A2(n_0_393_2), .ZN(n_0_393_1));
   INV_X1 i_0_393_3 (.A(in_data[0]), .ZN(n_0_393_2));
   INV_X1 i_0_394_0 (.A(n_0_394_0), .ZN(n_0_348));
   OAI21_X1 i_0_394_1 (.A(n_0_394_1), .B1(n_1150), .B2(n_0_637), .ZN(n_0_394_0));
   NAND2_X1 i_0_394_2 (.A1(n_0_637), .A2(n_0_394_2), .ZN(n_0_394_1));
   INV_X1 i_0_394_3 (.A(in_data[0]), .ZN(n_0_394_2));
   INV_X1 i_0_395_0 (.A(n_0_395_0), .ZN(n_0_349));
   OAI21_X1 i_0_395_1 (.A(n_0_395_1), .B1(n_0_121), .B2(n_0_640), .ZN(n_0_395_0));
   NAND2_X1 i_0_395_2 (.A1(n_0_640), .A2(n_0_395_2), .ZN(n_0_395_1));
   INV_X1 i_0_395_3 (.A(in_data[0]), .ZN(n_0_395_2));
   INV_X1 i_0_396_0 (.A(n_0_643), .ZN(n_0_396_0));
   AOI22_X1 i_0_396_1 (.A1(n_0_396_0), .A2(n_1174), .B1(in_data[0]), .B2(n_0_643), 
      .ZN(n_0_396_1));
   INV_X1 i_0_396_2 (.A(n_0_396_1), .ZN(n_0_350));
   INV_X1 i_0_397_0 (.A(n_0_397_0), .ZN(n_0_351));
   OAI21_X1 i_0_397_1 (.A(n_0_397_1), .B1(n_1151), .B2(n_0_646), .ZN(n_0_397_0));
   NAND2_X1 i_0_397_2 (.A1(n_0_646), .A2(n_0_397_2), .ZN(n_0_397_1));
   INV_X1 i_0_397_3 (.A(in_data[0]), .ZN(n_0_397_2));
   INV_X1 i_0_398_0 (.A(n_0_398_0), .ZN(n_0_352));
   OAI21_X1 i_0_398_1 (.A(n_0_398_1), .B1(n_1173), .B2(n_0_649), .ZN(n_0_398_0));
   NAND2_X1 i_0_398_2 (.A1(n_0_649), .A2(n_0_398_2), .ZN(n_0_398_1));
   INV_X1 i_0_398_3 (.A(in_data[0]), .ZN(n_0_398_2));
   INV_X1 i_0_399_0 (.A(n_0_399_0), .ZN(n_0_353));
   OAI21_X1 i_0_399_1 (.A(n_0_399_1), .B1(n_1152), .B2(n_0_652), .ZN(n_0_399_0));
   NAND2_X1 i_0_399_2 (.A1(n_0_652), .A2(n_0_399_2), .ZN(n_0_399_1));
   INV_X1 i_0_399_3 (.A(in_data[0]), .ZN(n_0_399_2));
   INV_X1 i_0_400_0 (.A(n_0_400_0), .ZN(n_0_354));
   OAI21_X1 i_0_400_1 (.A(n_0_400_1), .B1(n_1172), .B2(n_0_655), .ZN(n_0_400_0));
   NAND2_X1 i_0_400_2 (.A1(n_0_655), .A2(n_0_400_2), .ZN(n_0_400_1));
   INV_X1 i_0_400_3 (.A(in_data[0]), .ZN(n_0_400_2));
   INV_X1 i_0_401_0 (.A(n_0_658), .ZN(n_0_401_0));
   AOI22_X1 i_0_401_1 (.A1(n_0_401_0), .A2(n_1153), .B1(in_data[0]), .B2(n_0_658), 
      .ZN(n_0_401_1));
   INV_X1 i_0_401_2 (.A(n_0_401_1), .ZN(n_0_355));
   INV_X1 i_0_402_0 (.A(n_0_402_0), .ZN(n_0_356));
   OAI21_X1 i_0_402_1 (.A(n_0_402_1), .B1(n_1154), .B2(n_836), .ZN(n_0_402_0));
   NAND2_X1 i_0_402_2 (.A1(n_836), .A2(n_0_402_2), .ZN(n_0_402_1));
   INV_X1 i_0_402_3 (.A(in_data[0]), .ZN(n_0_402_2));
   INV_X1 i_0_403_0 (.A(n_0_403_0), .ZN(n_0_357));
   OAI21_X1 i_0_403_1 (.A(n_0_403_1), .B1(n_1155), .B2(n_676), .ZN(n_0_403_0));
   NAND2_X1 i_0_403_2 (.A1(n_676), .A2(n_0_403_2), .ZN(n_0_403_1));
   INV_X1 i_0_403_3 (.A(in_data[0]), .ZN(n_0_403_2));
   INV_X1 i_0_404_0 (.A(n_0_404_0), .ZN(n_0_358));
   OAI21_X1 i_0_404_1 (.A(n_0_404_1), .B1(n_1171), .B2(n_0_665), .ZN(n_0_404_0));
   NAND2_X1 i_0_404_2 (.A1(n_0_665), .A2(n_0_404_2), .ZN(n_0_404_1));
   INV_X1 i_0_404_3 (.A(in_data[0]), .ZN(n_0_404_2));
   INV_X1 i_0_405_0 (.A(n_0_405_0), .ZN(n_0_359));
   OAI21_X1 i_0_405_1 (.A(n_0_405_1), .B1(n_1156), .B2(n_0_668), .ZN(n_0_405_0));
   NAND2_X1 i_0_405_2 (.A1(n_0_668), .A2(n_0_405_2), .ZN(n_0_405_1));
   INV_X1 i_0_405_3 (.A(in_data[0]), .ZN(n_0_405_2));
   INV_X1 i_0_406_0 (.A(n_0_406_0), .ZN(n_0_360));
   OAI21_X1 i_0_406_1 (.A(n_0_406_1), .B1(n_1157), .B2(n_675), .ZN(n_0_406_0));
   NAND2_X1 i_0_406_2 (.A1(n_675), .A2(n_0_406_2), .ZN(n_0_406_1));
   INV_X1 i_0_406_3 (.A(in_data[0]), .ZN(n_0_406_2));
   INV_X1 i_0_407_0 (.A(n_0_407_0), .ZN(n_0_361));
   OAI21_X1 i_0_407_1 (.A(n_0_407_1), .B1(n_1084), .B2(n_0_673), .ZN(n_0_407_0));
   NAND2_X1 i_0_407_2 (.A1(n_0_673), .A2(n_0_407_2), .ZN(n_0_407_1));
   INV_X1 i_0_407_3 (.A(in_data[0]), .ZN(n_0_407_2));
   INV_X1 i_0_408_0 (.A(n_0_408_0), .ZN(n_0_362));
   OAI21_X1 i_0_408_1 (.A(n_0_408_1), .B1(n_1158), .B2(n_674), .ZN(n_0_408_0));
   NAND2_X1 i_0_408_2 (.A1(n_674), .A2(n_0_408_2), .ZN(n_0_408_1));
   INV_X1 i_0_408_3 (.A(in_data[0]), .ZN(n_0_408_2));
   INV_X1 i_0_409_0 (.A(n_0_409_0), .ZN(n_0_363));
   OAI21_X1 i_0_409_1 (.A(n_0_409_1), .B1(n_0_899), .B2(n_0_678), .ZN(n_0_409_0));
   NAND2_X1 i_0_409_2 (.A1(n_0_678), .A2(n_0_409_2), .ZN(n_0_409_1));
   INV_X1 i_0_409_3 (.A(in_data[0]), .ZN(n_0_409_2));
   INV_X1 i_0_410_0 (.A(n_0_410_0), .ZN(n_0_364));
   OAI21_X1 i_0_410_1 (.A(n_0_410_1), .B1(n_1085), .B2(n_0_681), .ZN(n_0_410_0));
   NAND2_X1 i_0_410_2 (.A1(n_0_681), .A2(n_0_410_2), .ZN(n_0_410_1));
   INV_X1 i_0_410_3 (.A(in_data[0]), .ZN(n_0_410_2));
   INV_X1 i_0_411_0 (.A(n_0_411_0), .ZN(n_0_365));
   OAI21_X1 i_0_411_1 (.A(n_0_411_1), .B1(n_1086), .B2(n_0_684), .ZN(n_0_411_0));
   NAND2_X1 i_0_411_2 (.A1(n_0_684), .A2(n_0_411_2), .ZN(n_0_411_1));
   INV_X1 i_0_411_3 (.A(in_data[0]), .ZN(n_0_411_2));
   INV_X1 i_0_412_0 (.A(n_0_412_0), .ZN(n_0_366));
   OAI21_X1 i_0_412_1 (.A(n_0_412_1), .B1(n_1159), .B2(n_673), .ZN(n_0_412_0));
   NAND2_X1 i_0_412_2 (.A1(n_673), .A2(n_0_412_2), .ZN(n_0_412_1));
   INV_X1 i_0_412_3 (.A(in_data[0]), .ZN(n_0_412_2));
   INV_X1 i_0_413_0 (.A(n_0_413_0), .ZN(n_0_367));
   OAI21_X1 i_0_413_1 (.A(n_0_413_1), .B1(n_1160), .B2(n_0_689), .ZN(n_0_413_0));
   NAND2_X1 i_0_413_2 (.A1(n_0_689), .A2(n_0_413_2), .ZN(n_0_413_1));
   INV_X1 i_0_413_3 (.A(in_data[0]), .ZN(n_0_413_2));
   INV_X1 i_0_414_0 (.A(n_0_414_0), .ZN(n_0_368));
   OAI21_X1 i_0_414_1 (.A(n_0_414_1), .B1(n_1161), .B2(n_672), .ZN(n_0_414_0));
   NAND2_X1 i_0_414_2 (.A1(n_672), .A2(n_0_414_2), .ZN(n_0_414_1));
   INV_X1 i_0_414_3 (.A(in_data[0]), .ZN(n_0_414_2));
   INV_X1 i_0_415_0 (.A(n_0_415_0), .ZN(n_0_369));
   OAI21_X1 i_0_415_1 (.A(n_0_415_1), .B1(n_1162), .B2(n_671), .ZN(n_0_415_0));
   NAND2_X1 i_0_415_2 (.A1(n_671), .A2(n_0_415_2), .ZN(n_0_415_1));
   INV_X1 i_0_415_3 (.A(in_data[0]), .ZN(n_0_415_2));
   INV_X1 i_0_416_0 (.A(n_0_416_0), .ZN(n_0_370));
   OAI21_X1 i_0_416_1 (.A(n_0_416_1), .B1(n_1163), .B2(n_670), .ZN(n_0_416_0));
   NAND2_X1 i_0_416_2 (.A1(n_670), .A2(n_0_416_2), .ZN(n_0_416_1));
   INV_X1 i_0_416_3 (.A(in_data[0]), .ZN(n_0_416_2));
   OAI21_X1 i_0_417_0 (.A(n_0_417_0), .B1(n_0_417_1), .B2(n_835), .ZN(n_0_371));
   NAND2_X1 i_0_417_1 (.A1(n_835), .A2(in_data[0]), .ZN(n_0_417_0));
   INV_X1 i_0_417_2 (.A(n_1164), .ZN(n_0_417_1));
   INV_X1 i_0_418_0 (.A(n_0_418_0), .ZN(n_0_372));
   OAI21_X1 i_0_418_1 (.A(n_0_418_1), .B1(n_1165), .B2(n_669), .ZN(n_0_418_0));
   NAND2_X1 i_0_418_2 (.A1(n_669), .A2(n_0_418_2), .ZN(n_0_418_1));
   INV_X1 i_0_418_3 (.A(in_data[0]), .ZN(n_0_418_2));
   INV_X1 i_0_419_0 (.A(n_0_419_0), .ZN(n_0_373));
   OAI21_X1 i_0_419_1 (.A(n_0_419_1), .B1(n_1087), .B2(n_0_702), .ZN(n_0_419_0));
   NAND2_X1 i_0_419_2 (.A1(n_0_702), .A2(n_0_419_2), .ZN(n_0_419_1));
   INV_X1 i_0_419_3 (.A(in_data[0]), .ZN(n_0_419_2));
   INV_X1 i_0_420_0 (.A(n_668), .ZN(n_0_420_0));
   AOI22_X1 i_0_420_1 (.A1(n_0_420_0), .A2(n_1166), .B1(in_data[0]), .B2(n_668), 
      .ZN(n_0_420_1));
   INV_X1 i_0_420_2 (.A(n_0_420_1), .ZN(n_0_374));
   INV_X1 i_0_421_0 (.A(n_667), .ZN(n_0_421_0));
   AOI22_X1 i_0_421_1 (.A1(n_0_421_0), .A2(n_1167), .B1(in_data[0]), .B2(n_667), 
      .ZN(n_0_421_1));
   INV_X1 i_0_421_2 (.A(n_0_421_1), .ZN(n_0_375));
   INV_X1 i_0_422_0 (.A(n_0_422_0), .ZN(n_0_376));
   OAI21_X1 i_0_422_1 (.A(n_0_422_1), .B1(n_0_900), .B2(n_0_709), .ZN(n_0_422_0));
   NAND2_X1 i_0_422_2 (.A1(n_0_709), .A2(n_0_422_2), .ZN(n_0_422_1));
   INV_X1 i_0_422_3 (.A(in_data[0]), .ZN(n_0_422_2));
   INV_X1 i_0_423_0 (.A(n_0_423_0), .ZN(n_0_377));
   OAI21_X1 i_0_423_1 (.A(n_0_423_1), .B1(n_0_901), .B2(n_0_712), .ZN(n_0_423_0));
   NAND2_X1 i_0_423_2 (.A1(n_0_712), .A2(n_0_423_2), .ZN(n_0_423_1));
   INV_X1 i_0_423_3 (.A(in_data[0]), .ZN(n_0_423_2));
   INV_X1 i_0_424_0 (.A(n_0_424_0), .ZN(n_0_378));
   OAI21_X1 i_0_424_1 (.A(n_0_424_1), .B1(n_1168), .B2(n_666), .ZN(n_0_424_0));
   NAND2_X1 i_0_424_2 (.A1(n_666), .A2(n_0_424_2), .ZN(n_0_424_1));
   INV_X1 i_0_424_3 (.A(in_data[0]), .ZN(n_0_424_2));
   INV_X1 i_0_425_0 (.A(n_0_425_0), .ZN(n_0_379));
   OAI21_X1 i_0_425_1 (.A(n_0_425_1), .B1(n_1169), .B2(n_665), .ZN(n_0_425_0));
   NAND2_X1 i_0_425_2 (.A1(n_665), .A2(n_0_425_2), .ZN(n_0_425_1));
   INV_X1 i_0_425_3 (.A(in_data[0]), .ZN(n_0_425_2));
   INV_X1 i_0_426_0 (.A(n_0_426_0), .ZN(n_0_380));
   OAI21_X1 i_0_426_1 (.A(n_0_426_1), .B1(n_1170), .B2(n_664), .ZN(n_0_426_0));
   NAND2_X1 i_0_426_2 (.A1(n_664), .A2(n_0_426_2), .ZN(n_0_426_1));
   INV_X1 i_0_426_3 (.A(in_data[0]), .ZN(n_0_426_2));
   INV_X1 i_0_427_0 (.A(n_0_427_0), .ZN(n_0_381));
   OAI21_X1 i_0_427_1 (.A(n_0_427_1), .B1(n_1091), .B2(n_0_79), .ZN(n_0_427_0));
   NAND2_X1 i_0_427_2 (.A1(n_0_79), .A2(n_0_427_2), .ZN(n_0_427_1));
   INV_X1 i_0_427_3 (.A(in_data[0]), .ZN(n_0_427_2));
   INV_X1 i_0_428_0 (.A(n_0_428_0), .ZN(n_0_382));
   OAI21_X1 i_0_428_1 (.A(n_0_428_1), .B1(n_1092), .B2(n_0_92), .ZN(n_0_428_0));
   NAND2_X1 i_0_428_2 (.A1(n_0_92), .A2(n_0_428_2), .ZN(n_0_428_1));
   INV_X1 i_0_428_3 (.A(in_data[0]), .ZN(n_0_428_2));
   INV_X1 i_0_429_0 (.A(n_0_78), .ZN(n_0_429_0));
   AOI22_X1 i_0_429_1 (.A1(n_0_429_0), .A2(n_1093), .B1(in_data[0]), .B2(n_0_78), 
      .ZN(n_0_429_1));
   INV_X1 i_0_429_2 (.A(n_0_429_1), .ZN(n_0_383));
   INV_X1 i_0_430_0 (.A(n_0_430_0), .ZN(n_0_384));
   OAI21_X1 i_0_430_1 (.A(n_0_430_1), .B1(n_1096), .B2(n_0_77), .ZN(n_0_430_0));
   NAND2_X1 i_0_430_2 (.A1(n_0_77), .A2(n_0_430_2), .ZN(n_0_430_1));
   INV_X1 i_0_430_3 (.A(in_data[0]), .ZN(n_0_430_2));
   OAI21_X1 i_0_431_0 (.A(n_0_431_0), .B1(n_0_431_1), .B2(n_0_91), .ZN(n_0_385));
   NAND2_X1 i_0_431_1 (.A1(n_0_91), .A2(in_data[0]), .ZN(n_0_431_0));
   INV_X1 i_0_431_2 (.A(n_974), .ZN(n_0_431_1));
   INV_X1 i_0_432_0 (.A(n_0_432_0), .ZN(n_0_386));
   OAI21_X1 i_0_432_1 (.A(n_0_432_1), .B1(n_1097), .B2(n_0_54), .ZN(n_0_432_0));
   NAND2_X1 i_0_432_2 (.A1(n_0_54), .A2(n_0_432_2), .ZN(n_0_432_1));
   INV_X1 i_0_432_3 (.A(in_data[0]), .ZN(n_0_432_2));
   INV_X1 i_0_433_0 (.A(n_0_433_0), .ZN(n_0_387));
   OAI21_X1 i_0_433_1 (.A(n_0_433_1), .B1(n_1098), .B2(n_0_75), .ZN(n_0_433_0));
   NAND2_X1 i_0_433_2 (.A1(n_0_75), .A2(n_0_433_2), .ZN(n_0_433_1));
   INV_X1 i_0_433_3 (.A(in_data[0]), .ZN(n_0_433_2));
   INV_X1 i_0_434_0 (.A(n_0_434_0), .ZN(n_0_388));
   OAI21_X1 i_0_434_1 (.A(n_0_434_1), .B1(n_1099), .B2(n_0_52), .ZN(n_0_434_0));
   NAND2_X1 i_0_434_2 (.A1(n_0_52), .A2(n_0_434_2), .ZN(n_0_434_1));
   INV_X1 i_0_434_3 (.A(in_data[0]), .ZN(n_0_434_2));
   INV_X1 i_0_435_0 (.A(n_0_90), .ZN(n_0_435_0));
   AOI22_X1 i_0_435_1 (.A1(n_0_435_0), .A2(n_1100), .B1(in_data[0]), .B2(n_0_90), 
      .ZN(n_0_435_1));
   INV_X1 i_0_435_2 (.A(n_0_435_1), .ZN(n_0_389));
   INV_X1 i_0_436_0 (.A(n_0_51), .ZN(n_0_436_0));
   AOI22_X1 i_0_436_1 (.A1(n_0_436_0), .A2(n_1101), .B1(in_data[0]), .B2(n_0_51), 
      .ZN(n_0_436_1));
   INV_X1 i_0_436_2 (.A(n_0_436_1), .ZN(n_0_391));
   INV_X1 i_0_437_0 (.A(n_0_437_0), .ZN(n_0_394));
   OAI21_X1 i_0_437_1 (.A(n_0_437_1), .B1(n_1102), .B2(n_0_74), .ZN(n_0_437_0));
   NAND2_X1 i_0_437_2 (.A1(n_0_74), .A2(n_0_437_2), .ZN(n_0_437_1));
   INV_X1 i_0_437_3 (.A(in_data[0]), .ZN(n_0_437_2));
   INV_X1 i_0_438_0 (.A(n_0_50), .ZN(n_0_438_0));
   AOI22_X1 i_0_438_1 (.A1(n_0_438_0), .A2(n_1103), .B1(in_data[0]), .B2(n_0_50), 
      .ZN(n_0_438_1));
   INV_X1 i_0_438_2 (.A(n_0_438_1), .ZN(n_0_396));
   INV_X1 i_0_439_0 (.A(n_0_439_0), .ZN(n_0_399));
   OAI21_X1 i_0_439_1 (.A(n_0_439_1), .B1(n_1104), .B2(n_0_49), .ZN(n_0_439_0));
   NAND2_X1 i_0_439_2 (.A1(n_0_49), .A2(n_0_439_2), .ZN(n_0_439_1));
   INV_X1 i_0_439_3 (.A(in_data[0]), .ZN(n_0_439_2));
   INV_X1 i_0_440_0 (.A(n_0_48), .ZN(n_0_440_0));
   AOI22_X1 i_0_440_1 (.A1(n_0_440_0), .A2(n_1105), .B1(in_data[0]), .B2(n_0_48), 
      .ZN(n_0_440_1));
   INV_X1 i_0_440_2 (.A(n_0_440_1), .ZN(n_0_402));
   INV_X1 i_0_441_0 (.A(n_0_441_0), .ZN(n_0_407));
   OAI21_X1 i_0_441_1 (.A(n_0_441_1), .B1(n_1106), .B2(n_0_46), .ZN(n_0_441_0));
   NAND2_X1 i_0_441_2 (.A1(n_0_46), .A2(n_0_441_2), .ZN(n_0_441_1));
   INV_X1 i_0_441_3 (.A(in_data[0]), .ZN(n_0_441_2));
   INV_X1 i_0_442_0 (.A(n_0_118), .ZN(n_0_442_0));
   AOI22_X1 i_0_442_1 (.A1(n_0_442_0), .A2(n_1107), .B1(in_data[0]), .B2(n_0_118), 
      .ZN(n_0_442_1));
   INV_X1 i_0_442_2 (.A(n_0_442_1), .ZN(n_0_410));
   OAI21_X1 i_0_443_0 (.A(n_0_443_0), .B1(n_0_443_1), .B2(n_0_45), .ZN(n_0_413));
   NAND2_X1 i_0_443_1 (.A1(n_0_45), .A2(in_data[0]), .ZN(n_0_443_0));
   INV_X1 i_0_443_2 (.A(n_1108), .ZN(n_0_443_1));
   OAI21_X1 i_0_444_0 (.A(n_0_444_0), .B1(n_0_444_1), .B2(n_0_72), .ZN(n_0_416));
   NAND2_X1 i_0_444_1 (.A1(n_0_72), .A2(in_data[0]), .ZN(n_0_444_0));
   INV_X1 i_0_444_2 (.A(n_1109), .ZN(n_0_444_1));
   OAI21_X1 i_0_445_0 (.A(n_0_445_0), .B1(n_0_445_1), .B2(n_0_44), .ZN(n_0_419));
   NAND2_X1 i_0_445_1 (.A1(n_0_44), .A2(in_data[0]), .ZN(n_0_445_0));
   INV_X1 i_0_445_2 (.A(n_0_124), .ZN(n_0_445_1));
   OAI21_X1 i_0_446_0 (.A(n_0_446_0), .B1(n_0_446_1), .B2(n_0_88), .ZN(n_0_422));
   NAND2_X1 i_0_446_1 (.A1(n_0_88), .A2(in_data[0]), .ZN(n_0_446_0));
   INV_X1 i_0_446_2 (.A(n_0_123), .ZN(n_0_446_1));
   INV_X1 i_0_447_0 (.A(n_0_71), .ZN(n_0_447_0));
   AOI22_X1 i_0_447_1 (.A1(n_0_447_0), .A2(n_1110), .B1(in_data[0]), .B2(n_0_71), 
      .ZN(n_0_447_1));
   INV_X1 i_0_447_2 (.A(n_0_447_1), .ZN(n_0_425));
   INV_X1 i_0_448_0 (.A(n_0_448_0), .ZN(n_0_428));
   OAI21_X1 i_0_448_1 (.A(n_0_448_1), .B1(n_0_100), .B2(n_0_42), .ZN(n_0_448_0));
   NAND2_X1 i_0_448_2 (.A1(n_0_42), .A2(n_0_448_2), .ZN(n_0_448_1));
   INV_X1 i_0_448_3 (.A(in_data[0]), .ZN(n_0_448_2));
   INV_X1 i_0_449_0 (.A(n_0_41), .ZN(n_0_449_0));
   AOI22_X1 i_0_449_1 (.A1(n_0_449_0), .A2(n_1111), .B1(in_data[0]), .B2(n_0_41), 
      .ZN(n_0_449_1));
   INV_X1 i_0_449_2 (.A(n_0_449_1), .ZN(n_0_431));
   INV_X1 i_0_450_0 (.A(n_0_70), .ZN(n_0_450_0));
   AOI22_X1 i_0_450_1 (.A1(n_0_450_0), .A2(n_1112), .B1(in_data[0]), .B2(n_0_70), 
      .ZN(n_0_450_1));
   INV_X1 i_0_450_2 (.A(n_0_450_1), .ZN(n_0_434));
   INV_X1 i_0_451_0 (.A(n_0_40), .ZN(n_0_451_0));
   AOI22_X1 i_0_451_1 (.A1(n_0_451_0), .A2(n_1113), .B1(in_data[0]), .B2(n_0_40), 
      .ZN(n_0_451_1));
   INV_X1 i_0_451_2 (.A(n_0_451_1), .ZN(n_0_436));
   INV_X1 i_0_452_0 (.A(n_0_37), .ZN(n_0_452_0));
   AOI22_X1 i_0_452_1 (.A1(n_0_452_0), .A2(n_0_101), .B1(in_data[0]), .B2(n_0_37), 
      .ZN(n_0_452_1));
   INV_X1 i_0_452_2 (.A(n_0_452_1), .ZN(n_0_439));
   INV_X1 i_0_453_0 (.A(n_0_68), .ZN(n_0_453_0));
   AOI22_X1 i_0_453_1 (.A1(n_0_453_0), .A2(n_1114), .B1(in_data[0]), .B2(n_0_68), 
      .ZN(n_0_453_1));
   INV_X1 i_0_453_2 (.A(n_0_453_1), .ZN(n_0_442));
   INV_X1 i_0_454_0 (.A(n_0_36), .ZN(n_0_454_0));
   AOI22_X1 i_0_454_1 (.A1(n_0_454_0), .A2(n_1115), .B1(in_data[0]), .B2(n_0_36), 
      .ZN(n_0_454_1));
   INV_X1 i_0_454_2 (.A(n_0_454_1), .ZN(n_0_445));
   INV_X1 i_0_455_0 (.A(n_0_86), .ZN(n_0_455_0));
   AOI22_X1 i_0_455_1 (.A1(n_0_455_0), .A2(n_1116), .B1(in_data[0]), .B2(n_0_86), 
      .ZN(n_0_455_1));
   INV_X1 i_0_455_2 (.A(n_0_455_1), .ZN(n_0_448));
   INV_X1 i_0_456_0 (.A(n_0_35), .ZN(n_0_456_0));
   AOI22_X1 i_0_456_1 (.A1(n_0_456_0), .A2(n_1117), .B1(in_data[0]), .B2(n_0_35), 
      .ZN(n_0_456_1));
   INV_X1 i_0_456_2 (.A(n_0_456_1), .ZN(n_0_451));
   INV_X1 i_0_457_0 (.A(n_0_67), .ZN(n_0_457_0));
   AOI22_X1 i_0_457_1 (.A1(n_0_457_0), .A2(n_1118), .B1(in_data[0]), .B2(n_0_67), 
      .ZN(n_0_457_1));
   INV_X1 i_0_457_2 (.A(n_0_457_1), .ZN(n_0_454));
   INV_X1 i_0_458_0 (.A(n_0_34), .ZN(n_0_458_0));
   AOI22_X1 i_0_458_1 (.A1(n_0_458_0), .A2(n_1119), .B1(in_data[0]), .B2(n_0_34), 
      .ZN(n_0_458_1));
   INV_X1 i_0_458_2 (.A(n_0_458_1), .ZN(n_0_455));
   INV_X1 i_0_459_0 (.A(n_0_96), .ZN(n_0_459_0));
   AOI22_X1 i_0_459_1 (.A1(n_0_459_0), .A2(n_1120), .B1(in_data[0]), .B2(n_0_96), 
      .ZN(n_0_459_1));
   INV_X1 i_0_459_2 (.A(n_0_459_1), .ZN(n_0_456));
   INV_X1 i_0_460_0 (.A(n_0_33), .ZN(n_0_460_0));
   AOI22_X1 i_0_460_1 (.A1(n_0_460_0), .A2(n_1121), .B1(in_data[0]), .B2(n_0_33), 
      .ZN(n_0_460_1));
   INV_X1 i_0_460_2 (.A(n_0_460_1), .ZN(n_0_459));
   INV_X1 i_0_461_0 (.A(n_0_66), .ZN(n_0_461_0));
   AOI22_X1 i_0_461_1 (.A1(n_0_461_0), .A2(n_1122), .B1(in_data[0]), .B2(n_0_66), 
      .ZN(n_0_461_1));
   INV_X1 i_0_461_2 (.A(n_0_461_1), .ZN(n_0_462));
   INV_X1 i_0_462_0 (.A(n_0_32), .ZN(n_0_462_0));
   AOI22_X1 i_0_462_1 (.A1(n_0_462_0), .A2(n_1123), .B1(in_data[0]), .B2(n_0_32), 
      .ZN(n_0_462_1));
   INV_X1 i_0_462_2 (.A(n_0_462_1), .ZN(n_0_465));
   OAI21_X1 i_0_463_0 (.A(n_0_463_0), .B1(n_0_463_1), .B2(n_0_85), .ZN(n_0_468));
   NAND2_X1 i_0_463_1 (.A1(n_0_85), .A2(in_data[0]), .ZN(n_0_463_0));
   INV_X1 i_0_463_2 (.A(n_0_122), .ZN(n_0_463_1));
   INV_X1 i_0_464_0 (.A(n_0_31), .ZN(n_0_464_0));
   AOI22_X1 i_0_464_1 (.A1(n_0_464_0), .A2(n_1124), .B1(in_data[0]), .B2(n_0_31), 
      .ZN(n_0_464_1));
   INV_X1 i_0_464_2 (.A(n_0_464_1), .ZN(n_0_471));
   INV_X1 i_0_465_0 (.A(n_0_465_0), .ZN(n_0_474));
   OAI21_X1 i_0_465_1 (.A(n_0_465_1), .B1(n_1126), .B2(n_0_29), .ZN(n_0_465_0));
   NAND2_X1 i_0_465_2 (.A1(n_0_29), .A2(n_0_465_2), .ZN(n_0_465_1));
   INV_X1 i_0_465_3 (.A(in_data[0]), .ZN(n_0_465_2));
   INV_X1 i_0_466_0 (.A(n_0_466_0), .ZN(n_0_477));
   OAI21_X1 i_0_466_1 (.A(n_0_466_1), .B1(n_1127), .B2(n_0_65), .ZN(n_0_466_0));
   NAND2_X1 i_0_466_2 (.A1(n_0_65), .A2(n_0_466_2), .ZN(n_0_466_1));
   INV_X1 i_0_466_3 (.A(in_data[0]), .ZN(n_0_466_2));
   INV_X1 i_0_467_0 (.A(n_0_467_0), .ZN(n_0_480));
   OAI21_X1 i_0_467_1 (.A(n_0_467_1), .B1(n_1128), .B2(n_0_28), .ZN(n_0_467_0));
   NAND2_X1 i_0_467_2 (.A1(n_0_28), .A2(n_0_467_2), .ZN(n_0_467_1));
   INV_X1 i_0_467_3 (.A(in_data[0]), .ZN(n_0_467_2));
   INV_X1 i_0_468_0 (.A(n_0_468_0), .ZN(n_0_483));
   OAI21_X1 i_0_468_1 (.A(n_0_468_1), .B1(n_1129), .B2(n_0_27), .ZN(n_0_468_0));
   NAND2_X1 i_0_468_2 (.A1(n_0_27), .A2(n_0_468_2), .ZN(n_0_468_1));
   INV_X1 i_0_468_3 (.A(in_data[0]), .ZN(n_0_468_2));
   INV_X1 i_0_469_0 (.A(n_0_469_0), .ZN(n_0_486));
   OAI21_X1 i_0_469_1 (.A(n_0_469_1), .B1(n_1130), .B2(n_0_64), .ZN(n_0_469_0));
   NAND2_X1 i_0_469_2 (.A1(n_0_64), .A2(n_0_469_2), .ZN(n_0_469_1));
   INV_X1 i_0_469_3 (.A(in_data[0]), .ZN(n_0_469_2));
   INV_X1 i_0_470_0 (.A(n_0_470_0), .ZN(n_0_489));
   OAI21_X1 i_0_470_1 (.A(n_0_470_1), .B1(n_1131), .B2(n_0_26), .ZN(n_0_470_0));
   NAND2_X1 i_0_470_2 (.A1(n_0_26), .A2(n_0_470_2), .ZN(n_0_470_1));
   INV_X1 i_0_470_3 (.A(in_data[0]), .ZN(n_0_470_2));
   INV_X1 i_0_471_0 (.A(n_0_95), .ZN(n_0_471_0));
   AOI22_X1 i_0_471_1 (.A1(n_0_471_0), .A2(n_1132), .B1(in_data[0]), .B2(n_0_95), 
      .ZN(n_0_471_1));
   INV_X1 i_0_471_2 (.A(n_0_471_1), .ZN(n_0_492));
   INV_X1 i_0_472_0 (.A(n_0_25), .ZN(n_0_472_0));
   AOI22_X1 i_0_472_1 (.A1(n_0_472_0), .A2(n_1133), .B1(in_data[0]), .B2(n_0_25), 
      .ZN(n_0_472_1));
   INV_X1 i_0_472_2 (.A(n_0_472_1), .ZN(n_0_495));
   INV_X1 i_0_473_0 (.A(n_0_63), .ZN(n_0_473_0));
   AOI22_X1 i_0_473_1 (.A1(n_0_473_0), .A2(n_1134), .B1(in_data[0]), .B2(n_0_63), 
      .ZN(n_0_473_1));
   INV_X1 i_0_473_2 (.A(n_0_473_1), .ZN(n_0_498));
   INV_X1 i_0_474_0 (.A(n_0_24), .ZN(n_0_474_0));
   AOI22_X1 i_0_474_1 (.A1(n_0_474_0), .A2(n_1135), .B1(in_data[0]), .B2(n_0_24), 
      .ZN(n_0_474_1));
   INV_X1 i_0_474_2 (.A(n_0_474_1), .ZN(n_0_501));
   INV_X1 i_0_475_0 (.A(n_0_475_0), .ZN(n_0_504));
   OAI21_X1 i_0_475_1 (.A(n_0_475_1), .B1(n_1136), .B2(n_0_23), .ZN(n_0_475_0));
   NAND2_X1 i_0_475_2 (.A1(n_0_23), .A2(n_0_475_2), .ZN(n_0_475_1));
   INV_X1 i_0_475_3 (.A(in_data[0]), .ZN(n_0_475_2));
   INV_X1 i_0_476_0 (.A(n_0_62), .ZN(n_0_476_0));
   AOI22_X1 i_0_476_1 (.A1(n_0_476_0), .A2(n_1137), .B1(in_data[0]), .B2(n_0_62), 
      .ZN(n_0_476_1));
   INV_X1 i_0_476_2 (.A(n_0_476_1), .ZN(n_0_507));
   INV_X1 i_0_477_0 (.A(n_0_22), .ZN(n_0_477_0));
   AOI22_X1 i_0_477_1 (.A1(n_0_477_0), .A2(n_1138), .B1(in_data[0]), .B2(n_0_22), 
      .ZN(n_0_477_1));
   INV_X1 i_0_477_2 (.A(n_0_477_1), .ZN(n_0_510));
   INV_X1 i_0_478_0 (.A(n_0_478_0), .ZN(n_0_513));
   OAI21_X1 i_0_478_1 (.A(n_0_478_1), .B1(n_1139), .B2(n_0_117), .ZN(n_0_478_0));
   NAND2_X1 i_0_478_2 (.A1(n_0_117), .A2(n_0_478_2), .ZN(n_0_478_1));
   INV_X1 i_0_478_3 (.A(in_data[0]), .ZN(n_0_478_2));
   INV_X1 i_0_479_0 (.A(n_0_21), .ZN(n_0_479_0));
   AOI22_X1 i_0_479_1 (.A1(n_0_479_0), .A2(n_1140), .B1(in_data[0]), .B2(n_0_21), 
      .ZN(n_0_479_1));
   INV_X1 i_0_479_2 (.A(n_0_479_1), .ZN(n_0_516));
   INV_X1 i_0_480_0 (.A(n_0_61), .ZN(n_0_480_0));
   AOI22_X1 i_0_480_1 (.A1(n_0_480_0), .A2(n_1141), .B1(in_data[0]), .B2(n_0_61), 
      .ZN(n_0_480_1));
   INV_X1 i_0_480_2 (.A(n_0_480_1), .ZN(n_0_519));
   INV_X1 i_0_481_0 (.A(n_0_20), .ZN(n_0_481_0));
   AOI22_X1 i_0_481_1 (.A1(n_0_481_0), .A2(n_1142), .B1(in_data[0]), .B2(n_0_20), 
      .ZN(n_0_481_1));
   INV_X1 i_0_481_2 (.A(n_0_481_1), .ZN(n_0_522));
   INV_X1 i_0_482_0 (.A(n_0_482_0), .ZN(n_0_525));
   OAI21_X1 i_0_482_1 (.A(n_0_482_1), .B1(n_1143), .B2(n_0_82), .ZN(n_0_482_0));
   NAND2_X1 i_0_482_2 (.A1(n_0_82), .A2(n_0_482_2), .ZN(n_0_482_1));
   INV_X1 i_0_482_3 (.A(in_data[0]), .ZN(n_0_482_2));
   INV_X1 i_0_483_0 (.A(n_0_19), .ZN(n_0_483_0));
   AOI22_X1 i_0_483_1 (.A1(n_0_483_0), .A2(n_1144), .B1(in_data[0]), .B2(n_0_19), 
      .ZN(n_0_483_1));
   INV_X1 i_0_483_2 (.A(n_0_483_1), .ZN(n_0_528));
   INV_X1 i_0_484_0 (.A(n_0_60), .ZN(n_0_484_0));
   AOI22_X1 i_0_484_1 (.A1(n_0_484_0), .A2(n_1145), .B1(in_data[0]), .B2(n_0_60), 
      .ZN(n_0_484_1));
   INV_X1 i_0_484_2 (.A(n_0_484_1), .ZN(n_0_531));
   INV_X1 i_0_485_0 (.A(n_0_485_0), .ZN(n_0_534));
   OAI21_X1 i_0_485_1 (.A(n_0_485_1), .B1(n_1146), .B2(n_0_18), .ZN(n_0_485_0));
   NAND2_X1 i_0_485_2 (.A1(n_0_18), .A2(n_0_485_2), .ZN(n_0_485_1));
   INV_X1 i_0_485_3 (.A(in_data[0]), .ZN(n_0_485_2));
   INV_X1 i_0_486_0 (.A(n_0_94), .ZN(n_0_486_0));
   AOI22_X1 i_0_486_1 (.A1(n_0_486_0), .A2(n_1147), .B1(in_data[0]), .B2(n_0_94), 
      .ZN(n_0_486_1));
   INV_X1 i_0_486_2 (.A(n_0_486_1), .ZN(n_0_537));
   INV_X1 i_0_487_0 (.A(n_0_487_0), .ZN(n_0_540));
   OAI21_X1 i_0_487_1 (.A(n_0_487_1), .B1(n_1148), .B2(n_0_17), .ZN(n_0_487_0));
   NAND2_X1 i_0_487_2 (.A1(n_0_17), .A2(n_0_487_2), .ZN(n_0_487_1));
   INV_X1 i_0_487_3 (.A(in_data[0]), .ZN(n_0_487_2));
   INV_X1 i_0_488_0 (.A(n_0_81), .ZN(n_0_488_0));
   AOI22_X1 i_0_488_1 (.A1(n_0_488_0), .A2(n_1149), .B1(in_data[0]), .B2(n_0_81), 
      .ZN(n_0_488_1));
   INV_X1 i_0_488_2 (.A(n_0_488_1), .ZN(n_0_543));
   INV_X1 i_0_489_0 (.A(n_0_58), .ZN(n_0_489_0));
   AOI22_X1 i_0_489_1 (.A1(n_0_489_0), .A2(n_1150), .B1(in_data[0]), .B2(n_0_58), 
      .ZN(n_0_489_1));
   INV_X1 i_0_489_2 (.A(n_0_489_1), .ZN(n_0_547));
   INV_X1 i_0_490_0 (.A(n_0_490_0), .ZN(n_0_548));
   OAI21_X1 i_0_490_1 (.A(n_0_490_1), .B1(n_1151), .B2(n_0_13), .ZN(n_0_490_0));
   NAND2_X1 i_0_490_2 (.A1(n_0_13), .A2(n_0_490_2), .ZN(n_0_490_1));
   INV_X1 i_0_490_3 (.A(in_data[0]), .ZN(n_0_490_2));
   INV_X1 i_0_491_0 (.A(n_0_12), .ZN(n_0_491_0));
   AOI22_X1 i_0_491_1 (.A1(n_0_491_0), .A2(n_1152), .B1(in_data[0]), .B2(n_0_12), 
      .ZN(n_0_491_1));
   INV_X1 i_0_491_2 (.A(n_0_491_1), .ZN(n_0_549));
   INV_X1 i_0_492_0 (.A(n_0_492_0), .ZN(n_0_552));
   OAI21_X1 i_0_492_1 (.A(n_0_492_1), .B1(n_1153), .B2(n_0_11), .ZN(n_0_492_0));
   NAND2_X1 i_0_492_2 (.A1(n_0_11), .A2(n_0_492_2), .ZN(n_0_492_1));
   INV_X1 i_0_492_3 (.A(in_data[0]), .ZN(n_0_492_2));
   INV_X1 i_0_493_0 (.A(n_0_493_0), .ZN(n_0_555));
   OAI21_X1 i_0_493_1 (.A(n_0_493_1), .B1(n_1154), .B2(n_0_111), .ZN(n_0_493_0));
   NAND2_X1 i_0_493_2 (.A1(n_0_111), .A2(n_0_493_2), .ZN(n_0_493_1));
   INV_X1 i_0_493_3 (.A(in_data[0]), .ZN(n_0_493_2));
   INV_X1 i_0_494_0 (.A(n_0_494_0), .ZN(n_0_558));
   OAI21_X1 i_0_494_1 (.A(n_0_494_1), .B1(n_1155), .B2(n_0_106), .ZN(n_0_494_0));
   NAND2_X1 i_0_494_2 (.A1(n_0_106), .A2(n_0_494_2), .ZN(n_0_494_1));
   INV_X1 i_0_494_3 (.A(in_data[0]), .ZN(n_0_494_2));
   INV_X1 i_0_495_0 (.A(n_0_10), .ZN(n_0_495_0));
   AOI22_X1 i_0_495_1 (.A1(n_0_495_0), .A2(n_1156), .B1(in_data[0]), .B2(n_0_10), 
      .ZN(n_0_495_1));
   INV_X1 i_0_495_2 (.A(n_0_495_1), .ZN(n_0_561));
   INV_X1 i_0_496_0 (.A(n_0_496_0), .ZN(n_0_564));
   OAI21_X1 i_0_496_1 (.A(n_0_496_1), .B1(n_1157), .B2(n_0_110), .ZN(n_0_496_0));
   NAND2_X1 i_0_496_2 (.A1(n_0_110), .A2(n_0_496_2), .ZN(n_0_496_1));
   INV_X1 i_0_496_3 (.A(in_data[0]), .ZN(n_0_496_2));
   INV_X1 i_0_497_0 (.A(n_0_497_0), .ZN(n_0_567));
   OAI21_X1 i_0_497_1 (.A(n_0_497_1), .B1(n_1158), .B2(n_0_114), .ZN(n_0_497_0));
   NAND2_X1 i_0_497_2 (.A1(n_0_114), .A2(n_0_497_2), .ZN(n_0_497_1));
   INV_X1 i_0_497_3 (.A(in_data[0]), .ZN(n_0_497_2));
   INV_X1 i_0_498_0 (.A(n_0_498_0), .ZN(n_0_570));
   OAI21_X1 i_0_498_1 (.A(n_0_498_1), .B1(n_1159), .B2(n_0_116), .ZN(n_0_498_0));
   NAND2_X1 i_0_498_2 (.A1(n_0_116), .A2(n_0_498_2), .ZN(n_0_498_1));
   INV_X1 i_0_498_3 (.A(in_data[0]), .ZN(n_0_498_2));
   INV_X1 i_0_499_0 (.A(n_0_499_0), .ZN(n_0_573));
   OAI21_X1 i_0_499_1 (.A(n_0_499_1), .B1(n_1160), .B2(n_0_6), .ZN(n_0_499_0));
   NAND2_X1 i_0_499_2 (.A1(n_0_6), .A2(n_0_499_2), .ZN(n_0_499_1));
   INV_X1 i_0_499_3 (.A(in_data[0]), .ZN(n_0_499_2));
   INV_X1 i_0_500_0 (.A(n_0_500_0), .ZN(n_0_576));
   OAI21_X1 i_0_500_1 (.A(n_0_500_1), .B1(n_1161), .B2(n_0_109), .ZN(n_0_500_0));
   NAND2_X1 i_0_500_2 (.A1(n_0_109), .A2(n_0_500_2), .ZN(n_0_500_1));
   INV_X1 i_0_500_3 (.A(in_data[0]), .ZN(n_0_500_2));
   INV_X1 i_0_501_0 (.A(n_0_501_0), .ZN(n_0_579));
   OAI21_X1 i_0_501_1 (.A(n_0_501_1), .B1(n_1162), .B2(n_0_105), .ZN(n_0_501_0));
   NAND2_X1 i_0_501_2 (.A1(n_0_105), .A2(n_0_501_2), .ZN(n_0_501_1));
   INV_X1 i_0_501_3 (.A(in_data[0]), .ZN(n_0_501_2));
   INV_X1 i_0_502_0 (.A(n_0_502_0), .ZN(n_0_582));
   OAI21_X1 i_0_502_1 (.A(n_0_502_1), .B1(n_1163), .B2(n_0_113), .ZN(n_0_502_0));
   NAND2_X1 i_0_502_2 (.A1(n_0_113), .A2(n_0_502_2), .ZN(n_0_502_1));
   INV_X1 i_0_502_3 (.A(in_data[0]), .ZN(n_0_502_2));
   INV_X1 i_0_503_0 (.A(n_0_503_0), .ZN(n_0_585));
   OAI21_X1 i_0_503_1 (.A(n_0_503_1), .B1(n_1164), .B2(n_0_104), .ZN(n_0_503_0));
   NAND2_X1 i_0_503_2 (.A1(n_0_104), .A2(n_0_503_2), .ZN(n_0_503_1));
   INV_X1 i_0_503_3 (.A(in_data[0]), .ZN(n_0_503_2));
   INV_X1 i_0_504_0 (.A(n_0_504_0), .ZN(n_0_588));
   OAI21_X1 i_0_504_1 (.A(n_0_504_1), .B1(n_1165), .B2(n_0_108), .ZN(n_0_504_0));
   NAND2_X1 i_0_504_2 (.A1(n_0_108), .A2(n_0_504_2), .ZN(n_0_504_1));
   INV_X1 i_0_504_3 (.A(in_data[0]), .ZN(n_0_504_2));
   INV_X1 i_0_505_0 (.A(n_0_115), .ZN(n_0_505_0));
   AOI22_X1 i_0_505_1 (.A1(n_0_505_0), .A2(n_1166), .B1(in_data[0]), .B2(n_0_115), 
      .ZN(n_0_505_1));
   INV_X1 i_0_505_2 (.A(n_0_505_1), .ZN(n_0_591));
   INV_X1 i_0_506_0 (.A(n_0_103), .ZN(n_0_506_0));
   AOI22_X1 i_0_506_1 (.A1(n_0_506_0), .A2(n_1167), .B1(in_data[0]), .B2(n_0_103), 
      .ZN(n_0_506_1));
   INV_X1 i_0_506_2 (.A(n_0_506_1), .ZN(n_0_594));
   INV_X1 i_0_507_0 (.A(n_0_112), .ZN(n_0_507_0));
   AOI22_X1 i_0_507_1 (.A1(n_0_507_0), .A2(n_1168), .B1(in_data[0]), .B2(n_0_112), 
      .ZN(n_0_507_1));
   INV_X1 i_0_507_2 (.A(n_0_507_1), .ZN(n_0_595));
   INV_X1 i_0_508_0 (.A(n_0_508_0), .ZN(n_0_596));
   OAI21_X1 i_0_508_1 (.A(n_0_508_1), .B1(n_1169), .B2(n_0_102), .ZN(n_0_508_0));
   NAND2_X1 i_0_508_2 (.A1(n_0_102), .A2(n_0_508_2), .ZN(n_0_508_1));
   INV_X1 i_0_508_3 (.A(in_data[0]), .ZN(n_0_508_2));
   INV_X1 i_0_509_0 (.A(n_0_509_0), .ZN(n_0_599));
   OAI21_X1 i_0_509_1 (.A(n_0_509_1), .B1(n_1170), .B2(n_0_107), .ZN(n_0_509_0));
   NAND2_X1 i_0_509_2 (.A1(n_0_107), .A2(n_0_509_2), .ZN(n_0_509_1));
   INV_X1 i_0_509_3 (.A(in_data[0]), .ZN(n_0_509_2));
   OAI21_X1 i_0_511_0 (.A(n_0_511_0), .B1(n_0_511_1), .B2(n_0_3), .ZN(n_0_602));
   NAND2_X1 i_0_511_1 (.A1(n_0_3), .A2(in_data[0]), .ZN(n_0_511_0));
   INV_X1 i_0_511_2 (.A(n_0_901), .ZN(n_0_511_1));
   INV_X1 i_0_512_0 (.A(n_0_512_0), .ZN(n_0_605));
   OAI21_X1 i_0_512_1 (.A(n_0_512_1), .B1(n_0_900), .B2(n_0_55), .ZN(n_0_512_0));
   NAND2_X1 i_0_512_2 (.A1(n_0_55), .A2(n_0_512_2), .ZN(n_0_512_1));
   INV_X1 i_0_512_3 (.A(in_data[0]), .ZN(n_0_512_2));
   INV_X1 i_0_513_0 (.A(n_0_513_0), .ZN(n_0_608));
   OAI21_X1 i_0_513_1 (.A(n_0_513_1), .B1(n_1087), .B2(n_0_4), .ZN(n_0_513_0));
   NAND2_X1 i_0_513_2 (.A1(n_0_4), .A2(n_0_513_2), .ZN(n_0_513_1));
   INV_X1 i_0_513_3 (.A(in_data[0]), .ZN(n_0_513_2));
   INV_X1 i_0_514_0 (.A(n_0_514_0), .ZN(n_0_611));
   OAI21_X1 i_0_514_1 (.A(n_0_514_1), .B1(n_1086), .B2(n_0_7), .ZN(n_0_514_0));
   NAND2_X1 i_0_514_2 (.A1(n_0_7), .A2(n_0_514_2), .ZN(n_0_514_1));
   INV_X1 i_0_514_3 (.A(in_data[0]), .ZN(n_0_514_2));
   INV_X1 i_0_515_0 (.A(n_0_515_0), .ZN(n_0_614));
   OAI21_X1 i_0_515_1 (.A(n_0_515_1), .B1(n_1085), .B2(n_0_56), .ZN(n_0_515_0));
   NAND2_X1 i_0_515_2 (.A1(n_0_56), .A2(n_0_515_2), .ZN(n_0_515_1));
   INV_X1 i_0_515_3 (.A(in_data[0]), .ZN(n_0_515_2));
   INV_X1 i_0_516_0 (.A(n_0_516_0), .ZN(n_0_617));
   OAI21_X1 i_0_516_1 (.A(n_0_516_1), .B1(n_0_899), .B2(n_0_8), .ZN(n_0_516_0));
   NAND2_X1 i_0_516_2 (.A1(n_0_8), .A2(n_0_516_2), .ZN(n_0_516_1));
   INV_X1 i_0_516_3 (.A(in_data[0]), .ZN(n_0_516_2));
   INV_X1 i_0_517_0 (.A(n_0_517_0), .ZN(n_0_620));
   OAI21_X1 i_0_517_1 (.A(n_0_517_1), .B1(n_1084), .B2(n_0_9), .ZN(n_0_517_0));
   NAND2_X1 i_0_517_2 (.A1(n_0_9), .A2(n_0_517_2), .ZN(n_0_517_1));
   INV_X1 i_0_517_3 (.A(in_data[0]), .ZN(n_0_517_2));
   INV_X1 i_0_518_0 (.A(n_0_518_0), .ZN(n_0_623));
   OAI21_X1 i_0_518_1 (.A(n_0_518_1), .B1(n_1171), .B2(n_0_93), .ZN(n_0_518_0));
   NAND2_X1 i_0_518_2 (.A1(n_0_93), .A2(n_0_518_2), .ZN(n_0_518_1));
   INV_X1 i_0_518_3 (.A(in_data[0]), .ZN(n_0_518_2));
   INV_X1 i_0_519_0 (.A(n_0_80), .ZN(n_0_519_0));
   AOI22_X1 i_0_519_1 (.A1(n_0_519_0), .A2(n_1172), .B1(in_data[0]), .B2(n_0_80), 
      .ZN(n_0_519_1));
   INV_X1 i_0_519_2 (.A(n_0_519_1), .ZN(n_0_626));
   INV_X1 i_0_520_0 (.A(n_0_57), .ZN(n_0_520_0));
   AOI22_X1 i_0_520_1 (.A1(n_0_520_0), .A2(n_1173), .B1(in_data[0]), .B2(n_0_57), 
      .ZN(n_0_520_1));
   INV_X1 i_0_520_2 (.A(n_0_520_1), .ZN(n_0_629));
   INV_X1 i_0_521_0 (.A(n_0_99), .ZN(n_0_521_0));
   AOI22_X1 i_0_521_1 (.A1(n_0_521_0), .A2(n_1174), .B1(in_data[0]), .B2(n_0_99), 
      .ZN(n_0_521_1));
   INV_X1 i_0_521_2 (.A(n_0_521_1), .ZN(n_0_632));
   INV_X1 i_0_522_0 (.A(n_0_522_0), .ZN(n_0_635));
   OAI21_X1 i_0_522_1 (.A(n_0_522_1), .B1(n_0_121), .B2(n_0_14), .ZN(n_0_522_0));
   NAND2_X1 i_0_522_2 (.A1(n_0_14), .A2(n_0_522_2), .ZN(n_0_522_1));
   INV_X1 i_0_522_3 (.A(in_data[0]), .ZN(n_0_522_2));
   INV_X1 i_0_523_0 (.A(n_0_15), .ZN(n_0_523_0));
   AOI22_X1 i_0_523_1 (.A1(n_0_523_0), .A2(n_1175), .B1(in_data[0]), .B2(n_0_15), 
      .ZN(n_0_523_1));
   INV_X1 i_0_523_2 (.A(n_0_523_1), .ZN(n_0_638));
   INV_X1 i_0_524_0 (.A(n_0_524_0), .ZN(n_0_641));
   OAI21_X1 i_0_524_1 (.A(n_0_524_1), .B1(n_0_898), .B2(n_0_16), .ZN(n_0_524_0));
   NAND2_X1 i_0_524_2 (.A1(n_0_16), .A2(n_0_524_2), .ZN(n_0_524_1));
   INV_X1 i_0_524_3 (.A(in_data[0]), .ZN(n_0_524_2));
   INV_X1 i_0_525_0 (.A(n_0_59), .ZN(n_0_525_0));
   AOI22_X1 i_0_525_1 (.A1(n_0_525_0), .A2(n_1176), .B1(in_data[0]), .B2(n_0_59), 
      .ZN(n_0_525_1));
   INV_X1 i_0_525_2 (.A(n_0_525_1), .ZN(n_0_644));
   INV_X1 i_0_526_0 (.A(n_0_83), .ZN(n_0_526_0));
   AOI22_X1 i_0_526_1 (.A1(n_0_526_0), .A2(n_1177), .B1(in_data[0]), .B2(n_0_83), 
      .ZN(n_0_526_1));
   INV_X1 i_0_526_2 (.A(n_0_526_1), .ZN(n_0_647));
   INV_X1 i_0_527_0 (.A(n_0_527_0), .ZN(n_0_650));
   OAI21_X1 i_0_527_1 (.A(n_0_527_1), .B1(n_1178), .B2(n_0_84), .ZN(n_0_527_0));
   NAND2_X1 i_0_527_2 (.A1(n_0_84), .A2(n_0_527_2), .ZN(n_0_527_1));
   INV_X1 i_0_527_3 (.A(in_data[0]), .ZN(n_0_527_2));
   INV_X1 i_0_528_0 (.A(n_0_30), .ZN(n_0_528_0));
   AOI22_X1 i_0_528_1 (.A1(n_0_528_0), .A2(n_1179), .B1(in_data[0]), .B2(n_0_30), 
      .ZN(n_0_528_1));
   INV_X1 i_0_528_2 (.A(n_0_528_1), .ZN(n_0_653));
   OAI21_X1 i_0_529_0 (.A(n_0_529_0), .B1(n_0_529_1), .B2(n_0_98), .ZN(n_0_656));
   NAND2_X1 i_0_529_1 (.A1(n_0_98), .A2(in_data[0]), .ZN(n_0_529_0));
   INV_X1 i_0_529_2 (.A(n_0_897), .ZN(n_0_529_1));
   INV_X1 i_0_530_0 (.A(n_0_38), .ZN(n_0_530_0));
   AOI22_X1 i_0_530_1 (.A1(n_0_530_0), .A2(n_1180), .B1(in_data[0]), .B2(n_0_38), 
      .ZN(n_0_530_1));
   INV_X1 i_0_530_2 (.A(n_0_530_1), .ZN(n_0_659));
   INV_X1 i_0_531_0 (.A(n_0_69), .ZN(n_0_531_0));
   AOI22_X1 i_0_531_1 (.A1(n_0_531_0), .A2(n_1181), .B1(in_data[0]), .B2(n_0_69), 
      .ZN(n_0_531_1));
   INV_X1 i_0_531_2 (.A(n_0_531_1), .ZN(n_0_660));
   INV_X1 i_0_532_0 (.A(n_0_39), .ZN(n_0_532_0));
   AOI22_X1 i_0_532_1 (.A1(n_0_532_0), .A2(n_1182), .B1(in_data[0]), .B2(n_0_39), 
      .ZN(n_0_532_1));
   INV_X1 i_0_532_2 (.A(n_0_532_1), .ZN(n_0_661));
   INV_X1 i_0_533_0 (.A(n_0_87), .ZN(n_0_533_0));
   AOI22_X1 i_0_533_1 (.A1(n_0_533_0), .A2(n_1183), .B1(in_data[0]), .B2(n_0_87), 
      .ZN(n_0_533_1));
   INV_X1 i_0_533_2 (.A(n_0_533_1), .ZN(n_0_662));
   INV_X1 i_0_534_0 (.A(n_0_97), .ZN(n_0_534_0));
   AOI22_X1 i_0_534_1 (.A1(n_0_534_0), .A2(n_1184), .B1(in_data[0]), .B2(n_0_97), 
      .ZN(n_0_534_1));
   INV_X1 i_0_534_2 (.A(n_0_534_1), .ZN(n_0_663));
   INV_X1 i_0_535_0 (.A(n_0_43), .ZN(n_0_535_0));
   AOI22_X1 i_0_535_1 (.A1(n_0_535_0), .A2(n_1185), .B1(in_data[0]), .B2(n_0_43), 
      .ZN(n_0_535_1));
   INV_X1 i_0_535_2 (.A(n_0_535_1), .ZN(n_0_666));
   INV_X1 i_0_536_0 (.A(n_0_47), .ZN(n_0_536_0));
   AOI22_X1 i_0_536_1 (.A1(n_0_536_0), .A2(n_1186), .B1(in_data[0]), .B2(n_0_47), 
      .ZN(n_0_536_1));
   INV_X1 i_0_536_2 (.A(n_0_536_1), .ZN(n_0_669));
   INV_X1 i_0_537_0 (.A(n_0_537_0), .ZN(n_0_670));
   OAI21_X1 i_0_537_1 (.A(n_0_537_1), .B1(n_0_896), .B2(n_0_89), .ZN(n_0_537_0));
   NAND2_X1 i_0_537_2 (.A1(n_0_89), .A2(n_0_537_2), .ZN(n_0_537_1));
   INV_X1 i_0_537_3 (.A(in_data[0]), .ZN(n_0_537_2));
   INV_X1 i_0_538_0 (.A(n_0_538_0), .ZN(n_0_671));
   OAI21_X1 i_0_538_1 (.A(n_0_538_1), .B1(n_1187), .B2(n_0_73), .ZN(n_0_538_0));
   NAND2_X1 i_0_538_2 (.A1(n_0_73), .A2(n_0_538_2), .ZN(n_0_538_1));
   INV_X1 i_0_538_3 (.A(in_data[0]), .ZN(n_0_538_2));
   INV_X1 i_0_539_0 (.A(n_0_53), .ZN(n_0_539_0));
   AOI22_X1 i_0_539_1 (.A1(n_0_539_0), .A2(n_1189), .B1(in_data[0]), .B2(n_0_53), 
      .ZN(n_0_539_1));
   INV_X1 i_0_539_2 (.A(n_0_539_1), .ZN(n_0_674));
   INV_X1 i_0_540_0 (.A(n_0_540_0), .ZN(n_0_675));
   OAI21_X1 i_0_540_1 (.A(n_0_540_1), .B1(n_0_895), .B2(n_0_76), .ZN(n_0_540_0));
   NAND2_X1 i_0_540_2 (.A1(n_0_76), .A2(n_0_540_2), .ZN(n_0_540_1));
   INV_X1 i_0_540_3 (.A(in_data[0]), .ZN(n_0_540_2));
   INV_X1 i_0_541_0 (.A(n_0_130), .ZN(n_0_541_0));
   AOI22_X1 i_0_541_1 (.A1(n_0_541_0), .A2(n_0_119), .B1(in_data[0]), .B2(
      n_0_130), .ZN(n_0_541_1));
   INV_X1 i_0_541_2 (.A(n_0_541_1), .ZN(n_0_676));
   OR2_X1 i_0_542_0 (.A1(n_1012), .A2(n_0_393), .ZN(n_0_679));
   NAND2_X1 i_0_543_0 (.A1(n_0_543_0), .A2(n_0_543_1), .ZN(n_0_682));
   INV_X1 i_0_543_1 (.A(n_0_395), .ZN(n_0_543_0));
   INV_X1 i_0_543_2 (.A(n_1013), .ZN(n_0_543_1));
   OR2_X1 i_0_544_0 (.A1(n_1014), .A2(n_0_398), .ZN(n_0_685));
   OR2_X1 i_0_545_0 (.A1(n_1266), .A2(n_0_401), .ZN(n_0_686));
   NAND2_X1 i_0_546_0 (.A1(n_0_546_0), .A2(n_0_546_1), .ZN(n_0_687));
   INV_X1 i_0_546_1 (.A(n_0_406), .ZN(n_0_546_0));
   INV_X1 i_0_546_2 (.A(n_1015), .ZN(n_0_546_1));
   NAND2_X1 i_0_547_0 (.A1(n_0_547_0), .A2(n_0_547_1), .ZN(n_0_690));
   INV_X1 i_0_547_1 (.A(n_0_409), .ZN(n_0_547_0));
   INV_X1 i_0_547_2 (.A(n_1017), .ZN(n_0_547_1));
   OR2_X1 i_0_548_0 (.A1(n_1261), .A2(n_0_412), .ZN(n_0_691));
   OR2_X1 i_0_549_0 (.A1(n_1018), .A2(n_0_415), .ZN(n_0_692));
   OR2_X1 i_0_550_0 (.A1(n_1258), .A2(n_0_418), .ZN(n_0_693));
   OR2_X1 i_0_551_0 (.A1(n_1257), .A2(n_0_421), .ZN(n_0_694));
   OR2_X1 i_0_552_0 (.A1(n_1256), .A2(n_0_424), .ZN(n_0_695));
   OR2_X1 i_0_553_0 (.A1(n_1019), .A2(n_0_427), .ZN(n_0_696));
   OR2_X1 i_0_554_0 (.A1(n_1255), .A2(n_0_430), .ZN(n_0_697));
   OR2_X1 i_0_555_0 (.A1(n_1254), .A2(n_0_433), .ZN(n_0_698));
   OR2_X1 i_0_556_0 (.A1(n_1253), .A2(n_0_435), .ZN(n_0_699));
   OR2_X1 i_0_557_0 (.A1(n_1020), .A2(n_0_438), .ZN(n_0_700));
   OR2_X1 i_0_558_0 (.A1(n_1021), .A2(n_0_441), .ZN(n_0_703));
   OR2_X1 i_0_559_0 (.A1(n_1022), .A2(n_0_444), .ZN(n_0_704));
   NAND2_X1 i_0_560_0 (.A1(n_0_560_0), .A2(n_0_560_1), .ZN(n_0_705));
   INV_X1 i_0_560_1 (.A(n_0_447), .ZN(n_0_560_0));
   INV_X1 i_0_560_2 (.A(n_1252), .ZN(n_0_560_1));
   OR2_X1 i_0_561_0 (.A1(n_1023), .A2(n_0_450), .ZN(n_0_706));
   OR2_X1 i_0_562_0 (.A1(n_1250), .A2(n_0_453), .ZN(n_0_707));
   OR2_X1 i_0_563_0 (.A1(n_1024), .A2(n_708), .ZN(n_0_710));
   NAND2_X1 i_0_564_0 (.A1(n_0_564_0), .A2(n_0_564_1), .ZN(n_0_713));
   INV_X1 i_0_564_1 (.A(n_0_458), .ZN(n_0_564_0));
   INV_X1 i_0_564_2 (.A(n_1025), .ZN(n_0_564_1));
   NAND2_X1 i_0_565_0 (.A1(n_0_565_0), .A2(n_0_565_1), .ZN(n_0_714));
   INV_X1 i_0_565_1 (.A(n_0_461), .ZN(n_0_565_0));
   INV_X1 i_0_565_2 (.A(n_1026), .ZN(n_0_565_1));
   NAND2_X1 i_0_566_0 (.A1(n_0_566_0), .A2(n_0_566_1), .ZN(n_0_715));
   INV_X1 i_0_566_1 (.A(n_0_464), .ZN(n_0_566_0));
   INV_X1 i_0_566_2 (.A(n_1027), .ZN(n_0_566_1));
   NAND2_X1 i_0_567_0 (.A1(n_0_567_0), .A2(n_0_567_1), .ZN(n_0_716));
   INV_X1 i_0_567_1 (.A(n_0_467), .ZN(n_0_567_0));
   INV_X1 i_0_567_2 (.A(n_1028), .ZN(n_0_567_1));
   OR2_X1 i_0_568_0 (.A1(n_1249), .A2(n_0_470), .ZN(n_0_717));
   OR2_X1 i_0_569_0 (.A1(n_1248), .A2(n_0_473), .ZN(n_0_718));
   NAND2_X1 i_0_570_0 (.A1(n_0_570_0), .A2(n_0_570_1), .ZN(n_0_719));
   INV_X1 i_0_570_1 (.A(n_0_476), .ZN(n_0_570_0));
   INV_X1 i_0_570_2 (.A(n_1247), .ZN(n_0_570_1));
   OR2_X1 i_0_571_0 (.A1(n_1029), .A2(n_0_479), .ZN(n_0_720));
   OR2_X1 i_0_572_0 (.A1(n_1030), .A2(n_0_482), .ZN(n_0_721));
   OR2_X1 i_0_573_0 (.A1(n_1031), .A2(n_0_485), .ZN(n_0_722));
   OR2_X1 i_0_574_0 (.A1(n_1032), .A2(n_0_488), .ZN(n_0_723));
   OR2_X1 i_0_575_0 (.A1(n_1246), .A2(n_0_491), .ZN(n_0_724));
   OR2_X1 i_0_576_0 (.A1(n_1033), .A2(n_0_494), .ZN(n_0_725));
   OR2_X1 i_0_577_0 (.A1(n_1034), .A2(n_0_497), .ZN(n_0_726));
   OR2_X1 i_0_578_0 (.A1(n_1035), .A2(n_0_500), .ZN(n_0_727));
   NAND2_X1 i_0_579_0 (.A1(n_0_579_0), .A2(n_0_579_1), .ZN(n_0_728));
   INV_X1 i_0_579_1 (.A(n_0_503), .ZN(n_0_579_0));
   INV_X1 i_0_579_2 (.A(n_1036), .ZN(n_0_579_1));
   OR2_X1 i_0_580_0 (.A1(n_1037), .A2(n_0_506), .ZN(n_0_729));
   OR2_X1 i_0_581_0 (.A1(n_1038), .A2(n_0_509), .ZN(n_0_730));
   OR2_X1 i_0_582_0 (.A1(n_1245), .A2(n_0_512), .ZN(n_0_731));
   OR2_X1 i_0_583_0 (.A1(n_1039), .A2(n_0_515), .ZN(n_0_732));
   OR2_X1 i_0_584_0 (.A1(n_1040), .A2(n_0_518), .ZN(n_0_733));
   OR2_X1 i_0_585_0 (.A1(n_1244), .A2(n_0_521), .ZN(n_0_734));
   OR2_X1 i_0_586_0 (.A1(n_1041), .A2(n_0_524), .ZN(n_0_735));
   OR2_X1 i_0_587_0 (.A1(n_1042), .A2(n_0_527), .ZN(n_0_736));
   OR2_X1 i_0_588_0 (.A1(n_1243), .A2(n_0_530), .ZN(n_0_737));
   OR2_X1 i_0_589_0 (.A1(n_1043), .A2(n_0_533), .ZN(n_0_738));
   OR2_X1 i_0_590_0 (.A1(n_1242), .A2(n_0_536), .ZN(n_0_739));
   NAND2_X1 i_0_591_0 (.A1(n_0_591_0), .A2(n_0_591_1), .ZN(n_0_740));
   INV_X1 i_0_591_1 (.A(n_0_539), .ZN(n_0_591_0));
   INV_X1 i_0_591_2 (.A(n_1044), .ZN(n_0_591_1));
   OR2_X1 i_0_592_0 (.A1(n_1241), .A2(n_0_542), .ZN(n_0_741));
   OR2_X1 i_0_593_0 (.A1(n_1239), .A2(n_0_546), .ZN(n_0_742));
   OR2_X1 i_0_594_0 (.A1(n_1238), .A2(n_837), .ZN(n_0_743));
   OR2_X1 i_0_595_0 (.A1(n_1237), .A2(n_0_551), .ZN(n_0_744));
   OR2_X1 i_0_596_0 (.A1(n_1045), .A2(n_0_554), .ZN(n_0_745));
   OR2_X1 i_0_597_0 (.A1(n_1046), .A2(n_0_557), .ZN(n_0_746));
   OR2_X1 i_0_598_0 (.A1(n_1047), .A2(n_0_560), .ZN(n_0_747));
   OR2_X1 i_0_599_0 (.A1(n_1048), .A2(n_0_563), .ZN(n_0_748));
   OR2_X1 i_0_600_0 (.A1(n_1049), .A2(n_0_566), .ZN(n_0_749));
   OR2_X1 i_0_601_0 (.A1(n_1050), .A2(n_0_569), .ZN(n_0_750));
   OR2_X1 i_0_602_0 (.A1(n_1051), .A2(n_0_572), .ZN(n_0_751));
   OR2_X1 i_0_603_0 (.A1(n_1052), .A2(n_0_575), .ZN(n_0_752));
   OR2_X1 i_0_604_0 (.A1(n_1053), .A2(n_0_578), .ZN(n_0_753));
   OR2_X1 i_0_605_0 (.A1(n_1054), .A2(n_0_581), .ZN(n_0_754));
   OR2_X1 i_0_606_0 (.A1(n_1055), .A2(n_0_584), .ZN(n_0_755));
   OR2_X1 i_0_607_0 (.A1(n_1056), .A2(n_0_587), .ZN(n_0_756));
   OR2_X1 i_0_608_0 (.A1(n_1236), .A2(n_0_590), .ZN(n_0_757));
   OR2_X1 i_0_609_0 (.A1(n_1235), .A2(n_0_593), .ZN(n_0_758));
   OR2_X1 i_0_610_0 (.A1(n_1057), .A2(n_677), .ZN(n_0_759));
   OR2_X1 i_0_611_0 (.A1(n_1234), .A2(n_0_598), .ZN(n_0_760));
   OR2_X1 i_0_612_0 (.A1(n_1058), .A2(n_0_601), .ZN(n_0_761));
   OR2_X1 i_0_613_0 (.A1(n_1233), .A2(n_0_604), .ZN(n_0_762));
   OR2_X1 i_0_614_0 (.A1(n_1232), .A2(n_0_607), .ZN(n_0_763));
   OR2_X1 i_0_615_0 (.A1(n_1231), .A2(n_0_610), .ZN(n_0_764));
   OR2_X1 i_0_616_0 (.A1(n_1059), .A2(n_0_613), .ZN(n_0_765));
   OR2_X1 i_0_617_0 (.A1(n_1060), .A2(n_0_616), .ZN(n_0_766));
   OR2_X1 i_0_618_0 (.A1(n_1061), .A2(n_0_619), .ZN(n_0_767));
   OR2_X1 i_0_619_0 (.A1(n_1062), .A2(n_0_622), .ZN(n_0_768));
   OR2_X1 i_0_620_0 (.A1(n_1063), .A2(n_0_625), .ZN(n_0_769));
   NAND2_X1 i_0_621_0 (.A1(n_0_621_0), .A2(n_0_621_1), .ZN(n_0_770));
   INV_X1 i_0_621_1 (.A(n_0_628), .ZN(n_0_621_0));
   INV_X1 i_0_621_2 (.A(n_1064), .ZN(n_0_621_1));
   OR2_X1 i_0_622_0 (.A1(n_1230), .A2(n_0_631), .ZN(n_0_771));
   OR2_X1 i_0_623_0 (.A1(n_1065), .A2(n_0_634), .ZN(n_0_772));
   OR2_X1 i_0_624_0 (.A1(n_1066), .A2(n_0_637), .ZN(n_0_773));
   OR2_X1 i_0_625_0 (.A1(n_1229), .A2(n_0_640), .ZN(n_0_774));
   OR2_X1 i_0_626_0 (.A1(n_1228), .A2(n_0_643), .ZN(n_0_775));
   OR2_X1 i_0_627_0 (.A1(n_1067), .A2(n_0_646), .ZN(n_0_776));
   OR2_X1 i_0_628_0 (.A1(n_1068), .A2(n_0_649), .ZN(n_0_777));
   OR2_X1 i_0_629_0 (.A1(n_1227), .A2(n_0_652), .ZN(n_0_778));
   OR2_X1 i_0_630_0 (.A1(n_1069), .A2(n_0_655), .ZN(n_0_779));
   OR2_X1 i_0_631_0 (.A1(n_1070), .A2(n_0_658), .ZN(n_0_780));
   OR2_X1 i_0_632_0 (.A1(n_836), .A2(n_1071), .ZN(n_0_781));
   OR2_X1 i_0_633_0 (.A1(n_1226), .A2(n_676), .ZN(n_0_782));
   OR2_X1 i_0_634_0 (.A1(n_1225), .A2(n_0_665), .ZN(n_0_783));
   OR2_X1 i_0_635_0 (.A1(n_1224), .A2(n_0_668), .ZN(n_0_784));
   OR2_X1 i_0_636_0 (.A1(n_1223), .A2(n_675), .ZN(n_0_785));
   OR2_X1 i_0_637_0 (.A1(n_1072), .A2(n_0_673), .ZN(n_0_786));
   OR2_X1 i_0_638_0 (.A1(n_1222), .A2(n_674), .ZN(n_0_787));
   OR2_X1 i_0_639_0 (.A1(n_1073), .A2(n_0_678), .ZN(n_0_788));
   OR2_X1 i_0_640_0 (.A1(n_1074), .A2(n_0_681), .ZN(n_0_789));
   OR2_X1 i_0_641_0 (.A1(n_1075), .A2(n_0_684), .ZN(n_0_790));
   OR2_X1 i_0_642_0 (.A1(n_1221), .A2(n_673), .ZN(n_0_791));
   OR2_X1 i_0_643_0 (.A1(n_1220), .A2(n_0_689), .ZN(n_0_792));
   OR2_X1 i_0_644_0 (.A1(n_1219), .A2(n_672), .ZN(n_0_793));
   OR2_X1 i_0_645_0 (.A1(n_1076), .A2(n_671), .ZN(n_0_794));
   OR2_X1 i_0_646_0 (.A1(n_1218), .A2(n_670), .ZN(n_0_795));
   OR2_X1 i_0_647_0 (.A1(n_1077), .A2(n_835), .ZN(n_0_796));
   OR2_X1 i_0_648_0 (.A1(n_1078), .A2(n_669), .ZN(n_0_797));
   OR2_X1 i_0_649_0 (.A1(n_1079), .A2(n_0_702), .ZN(n_0_798));
   OR2_X1 i_0_650_0 (.A1(n_1217), .A2(n_668), .ZN(n_0_799));
   OR2_X1 i_0_651_0 (.A1(n_1080), .A2(n_667), .ZN(n_0_800));
   OR2_X1 i_0_652_0 (.A1(n_1081), .A2(n_0_709), .ZN(n_0_801));
   OR2_X1 i_0_653_0 (.A1(n_1082), .A2(n_0_712), .ZN(n_0_802));
   OR2_X1 i_0_654_0 (.A1(n_1216), .A2(n_666), .ZN(n_0_803));
   OR2_X1 i_0_655_0 (.A1(n_1083), .A2(n_665), .ZN(n_0_804));
   OR2_X1 i_0_656_0 (.A1(n_1215), .A2(n_664), .ZN(n_0_805));
   OAI21_X1 i_0_658_0 (.A(n_0_658_0), .B1(n_0_658_3), .B2(n_0_658_1), .ZN(
      n_0_901));
   NAND2_X1 i_0_658_1 (.A1(n_1198), .A2(n_0_658_1), .ZN(n_0_658_0));
   OAI22_X1 i_0_658_2 (.A1(n_952), .A2(n_1211), .B1(n_0_658_2), .B2(n_1210), 
      .ZN(n_0_658_1));
   INV_X1 i_0_658_3 (.A(n_952), .ZN(n_0_658_2));
   INV_X1 i_0_658_4 (.A(in_data[4]), .ZN(n_0_658_3));
   DFF_X1 \buf_reg[127]  (.D(n_0_816), .CK(clk), .Q(n_857), .QN());
   DFF_X1 \buf_reg[126]  (.D(n_0_817), .CK(clk), .Q(n_858), .QN());
   DFF_X1 \buf_reg[125]  (.D(n_0_818), .CK(clk), .Q(n_859), .QN());
   DFF_X1 \buf_reg[124]  (.D(n_0_819), .CK(clk), .Q(n_860), .QN());
   DFF_X1 \buf_reg[121]  (.D(n_0_822), .CK(clk), .Q(n_861), .QN());
   DFF_X1 \buf_reg[120]  (.D(n_0_823), .CK(clk), .Q(n_862), .QN());
   DFF_X1 \buf_reg[119]  (.D(n_0_824), .CK(clk), .Q(n_863), .QN());
   DFF_X1 \buf_reg[117]  (.D(n_0_826), .CK(clk), .Q(n_864), .QN());
   DFF_X1 \buf_reg[116]  (.D(n_0_827), .CK(clk), .Q(n_865), .QN());
   DFF_X1 \buf_reg[114]  (.D(n_0_829), .CK(clk), .Q(n_866), .QN());
   DFF_X1 \buf_reg[113]  (.D(n_0_830), .CK(clk), .Q(n_867), .QN());
   DFF_X1 \buf_reg[112]  (.D(n_0_831), .CK(clk), .Q(n_868), .QN());
   DFF_X1 \buf_reg[111]  (.D(n_0_832), .CK(clk), .Q(n_869), .QN());
   DFF_X1 \buf_reg[110]  (.D(n_0_833), .CK(clk), .Q(n_870), .QN());
   DFF_X1 \buf_reg[108]  (.D(n_0_835), .CK(clk), .Q(n_871), .QN());
   DFF_X1 \buf_reg[107]  (.D(n_0_836), .CK(clk), .Q(n_872), .QN());
   DFF_X1 \buf_reg[106]  (.D(n_0_837), .CK(clk), .Q(n_873), .QN());
   DFF_X1 \buf_reg[105]  (.D(n_0_838), .CK(clk), .Q(n_874), .QN());
   DFF_X1 \buf_reg[104]  (.D(n_0_839), .CK(clk), .Q(n_875), .QN());
   DFF_X1 \buf_reg[103]  (.D(n_0_840), .CK(clk), .Q(n_876), .QN());
   DFF_X2 \buf_reg[101]  (.D(n_0_842), .CK(clk), .Q(n_877), .QN());
   DFF_X1 \buf_reg[100]  (.D(n_0_843), .CK(clk), .Q(n_878), .QN());
   DFF_X1 \buf_reg[99]  (.D(n_0_844), .CK(clk), .Q(n_879), .QN());
   DFF_X1 \buf_reg[98]  (.D(n_0_845), .CK(clk), .Q(n_880), .QN());
   DFF_X1 \buf_reg[97]  (.D(n_0_846), .CK(clk), .Q(n_881), .QN());
   DFF_X1 \buf_reg[94]  (.D(n_0_849), .CK(clk), .Q(n_882), .QN());
   DFF_X1 \buf_reg[93]  (.D(n_0_850), .CK(clk), .Q(n_883), .QN());
   DFF_X1 \buf_reg[92]  (.D(n_0_851), .CK(clk), .Q(n_884), .QN());
   DFF_X1 \buf_reg[90]  (.D(n_0_853), .CK(clk), .Q(n_885), .QN());
   DFF_X1 \buf_reg[89]  (.D(n_0_854), .CK(clk), .Q(n_886), .QN());
   DFF_X1 \buf_reg[87]  (.D(n_0_856), .CK(clk), .Q(n_887), .QN());
   DFF_X1 \buf_reg[85]  (.D(n_0_858), .CK(clk), .Q(n_888), .QN());
   DFF_X1 \buf_reg[84]  (.D(n_0_859), .CK(clk), .Q(n_889), .QN());
   DFF_X1 \buf_reg[83]  (.D(n_0_860), .CK(clk), .Q(n_890), .QN());
   DFF_X1 \buf_reg[81]  (.D(n_0_862), .CK(clk), .Q(n_891), .QN());
   DFF_X1 \buf_reg[80]  (.D(n_0_863), .CK(clk), .Q(n_892), .QN());
   DFF_X1 \buf_reg[79]  (.D(n_0_864), .CK(clk), .Q(n_893), .QN());
   DFF_X1 \buf_reg[78]  (.D(n_0_865), .CK(clk), .Q(n_894), .QN());
   DFF_X2 \buf_reg[77]  (.D(n_0_866), .CK(clk), .Q(n_895), .QN());
   DFF_X1 \buf_reg[76]  (.D(n_0_867), .CK(clk), .Q(n_896), .QN());
   DFF_X2 \buf_reg[71]  (.D(n_0_872), .CK(clk), .Q(n_897), .QN());
   DFF_X2 \buf_reg[70]  (.D(n_0_873), .CK(clk), .Q(n_898), .QN());
   DFF_X2 \buf_reg[69]  (.D(n_0_874), .CK(clk), .Q(n_899), .QN());
   DFF_X1 \buf_reg[68]  (.D(n_0_875), .CK(clk), .Q(n_900), .QN());
   DFF_X2 \buf_reg[67]  (.D(n_0_876), .CK(clk), .Q(n_901), .QN());
   DFF_X2 \buf_reg[66]  (.D(n_0_877), .CK(clk), .Q(n_902), .QN());
   DFF_X2 \buf_reg[65]  (.D(n_0_878), .CK(clk), .Q(n_903), .QN());
   DFF_X1 \buf_reg[63]  (.D(n_0_880), .CK(clk), .Q(n_904), .QN());
   DFF_X1 \buf_reg[62]  (.D(n_0_881), .CK(clk), .Q(n_905), .QN());
   DFF_X1 \buf_reg[61]  (.D(n_0_882), .CK(clk), .Q(n_906), .QN());
   DFF_X2 \buf_reg[60]  (.D(n_0_883), .CK(clk), .Q(n_907), .QN());
   DFF_X1 \buf_reg[59]  (.D(n_0_884), .CK(clk), .Q(n_908), .QN());
   DFF_X1 \buf_reg[57]  (.D(n_0_886), .CK(clk), .Q(n_909), .QN());
   DFF_X1 \buf_reg[54]  (.D(n_0_889), .CK(clk), .Q(n_910), .QN());
   DFF_X1 \buf_reg[51]  (.D(n_0_892), .CK(clk), .Q(n_911), .QN());
   DFF_X1 \buf_reg[50]  (.D(n_0_893), .CK(clk), .Q(n_912), .QN());
   DFF_X1 \buf_reg[49]  (.D(n_0_894), .CK(clk), .Q(n_913), .QN());
   DFF_X2 \buf_reg[48]  (.D(n_0_902), .CK(clk), .Q(n_914), .QN());
   DFF_X1 \buf_reg[44]  (.D(n_0_906), .CK(clk), .Q(n_915), .QN());
   DFF_X1 \buf_reg[38]  (.D(n_0_912), .CK(clk), .Q(n_916), .QN());
   DFF_X1 \buf_reg[37]  (.D(n_0_913), .CK(clk), .Q(n_917), .QN());
   DFF_X2 \buf_reg[36]  (.D(n_0_914), .CK(clk), .Q(n_918), .QN());
   DFF_X2 \buf_reg[35]  (.D(n_0_915), .CK(clk), .Q(n_919), .QN());
   DFF_X1 \buf_reg[34]  (.D(n_0_916), .CK(clk), .Q(n_920), .QN());
   DFF_X1 \buf_reg[33]  (.D(n_0_917), .CK(clk), .Q(n_921), .QN());
   DFF_X1 \buf_reg[32]  (.D(n_0_918), .CK(clk), .Q(n_922), .QN());
   DFF_X1 \buf_reg[31]  (.D(n_0_919), .CK(clk), .Q(n_923), .QN());
   DFF_X1 \buf_reg[30]  (.D(n_0_920), .CK(clk), .Q(n_924), .QN());
   DFF_X1 \buf_reg[29]  (.D(n_0_921), .CK(clk), .Q(n_925), .QN());
   DFF_X1 \buf_reg[27]  (.D(n_0_923), .CK(clk), .Q(n_926), .QN());
   DFF_X1 \buf_reg[26]  (.D(n_0_924), .CK(clk), .Q(n_927), .QN());
   DFF_X1 \buf_reg[25]  (.D(n_0_925), .CK(clk), .Q(n_928), .QN());
   DFF_X1 \buf_reg[24]  (.D(n_0_926), .CK(clk), .Q(n_929), .QN());
   DFF_X1 \buf_reg[23]  (.D(n_0_927), .CK(clk), .Q(n_930), .QN());
   DFF_X1 \buf_reg[22]  (.D(n_0_928), .CK(clk), .Q(n_931), .QN());
   DFF_X1 \buf_reg[21]  (.D(n_0_929), .CK(clk), .Q(n_932), .QN());
   DFF_X1 \buf_reg[20]  (.D(n_0_930), .CK(clk), .Q(n_933), .QN());
   DFF_X1 \buf_reg[19]  (.D(n_0_931), .CK(clk), .Q(n_934), .QN());
   DFF_X1 \buf_reg[18]  (.D(n_0_932), .CK(clk), .Q(n_935), .QN());
   DFF_X1 \buf_reg[17]  (.D(n_0_933), .CK(clk), .Q(n_936), .QN());
   DFF_X1 \buf_reg[16]  (.D(n_0_934), .CK(clk), .Q(n_937), .QN());
   DFF_X1 \buf_reg[13]  (.D(n_0_937), .CK(clk), .Q(n_938), .QN());
   DFF_X1 \buf_reg[12]  (.D(n_0_938), .CK(clk), .Q(n_939), .QN());
   DFF_X1 \buf_reg[11]  (.D(n_0_939), .CK(clk), .Q(n_940), .QN());
   DFF_X1 \buf_reg[10]  (.D(n_0_940), .CK(clk), .Q(n_941), .QN());
   DFF_X1 \buf_reg[9]  (.D(n_0_941), .CK(clk), .Q(n_942), .QN());
   DFF_X1 \buf_reg[8]  (.D(n_0_942), .CK(clk), .Q(n_943), .QN());
   DFF_X1 \buf_reg[7]  (.D(n_0_943), .CK(clk), .Q(n_944), .QN());
   DFF_X1 \buf_reg[6]  (.D(n_0_944), .CK(clk), .Q(n_945), .QN());
   DFF_X1 \buf_reg[5]  (.D(n_0_945), .CK(clk), .Q(n_946), .QN());
   DFF_X1 \buf_reg[4]  (.D(n_0_946), .CK(clk), .Q(n_947), .QN());
   DFF_X1 \buf_reg[2]  (.D(n_0_948), .CK(clk), .Q(n_948), .QN());
   DFF_X1 \buf_reg[1]  (.D(n_0_949), .CK(clk), .Q(n_949), .QN());
   DFF_X1 \buf_reg[0]  (.D(n_0_950), .CK(clk), .Q(n_950), .QN());
   DFF_X1 \buf_reg[15]  (.D(n_0_935), .CK(clk), .Q(n_951), .QN());
   range_extractor ranges_7_range_extr_i (.in_a(\out_bs[6] ), .in_size({
      in_data[3], in_data[2], in_data[1]}), .out_a(\out_as[7] ), .out_b(
      \out_bs[7] ));
   datapath__1_7663 i_0_660 (.\out_as[6] (\out_as[6] ), .\out_bs[6] (\out_bs[6] ), 
      .p_0(n_952));
   datapath__1_12443 i_0_510 (.\out_as[7] (\out_as[7] ), .\out_bs[7] (
      \out_bs[7] ), .p_0(n_0_806));
   datapath__1_14009 i_0_662 (.to_int6126({uc_149, \out_bs[7] [6], 
      \out_bs[7] [5], \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], 
      \out_bs[7] [1], \out_bs[7] [0]}), .p_0(n_953));
   datapath__1_13993 i_0_663 (.to_int6126({uc_150, \out_bs[7] [6], 
      \out_bs[7] [5], \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], 
      \out_bs[7] [1], \out_bs[7] [0]}), .p_0(n_954));
   datapath__1_13977 i_0_664 (.to_int6126({uc_151, \out_bs[7] [6], 
      \out_bs[7] [5], \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], 
      \out_bs[7] [1], \out_bs[7] [0]}), .p_0(n_955));
   datapath__1_13969 i_0_665 (.to_int6126({uc_152, \out_bs[7] [6], 
      \out_bs[7] [5], \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], 
      \out_bs[7] [1], \out_bs[7] [0]}), .p_0(n_956));
   datapath__1_13921 i_0_666 (.to_int6126({uc_153, \out_bs[7] [6], 
      \out_bs[7] [5], \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], 
      \out_bs[7] [1], \out_bs[7] [0]}), .p_0(n_957));
   datapath__1_14013 i_0_667 (.to_int6126({uc_154, \out_bs[7] [6], 
      \out_bs[7] [5], \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], 
      \out_bs[7] [1], uc_155}), .p_0(n_958));
   datapath__1_13981 i_0_668 (.to_int6126({uc_156, \out_bs[7] [6], 
      \out_bs[7] [5], \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], 
      \out_bs[7] [1], uc_157}), .p_0(n_959));
   datapath__1_13965 i_0_669 (.to_int6126({uc_158, \out_bs[7] [6], 
      \out_bs[7] [5], \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], 
      \out_bs[7] [1], uc_159}), .p_0(n_960));
   datapath__1_13933 i_0_670 (.to_int6126({uc_160, \out_bs[7] [6], 
      \out_bs[7] [5], \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], 
      \out_bs[7] [1], uc_161}), .p_0(n_961));
   datapath__1_13917 i_0_671 (.to_int6126({uc_162, \out_bs[7] [6], 
      \out_bs[7] [5], \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], 
      \out_bs[7] [1], uc_163}), .p_0(n_962));
   datapath__1_14005 i_0_672 (.to_int6126({uc_164, \out_bs[7] [6], 
      \out_bs[7] [5], \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], uc_165, 
      uc_166}), .p_0(n_963));
   datapath__1_13973 i_0_673 (.to_int6126({uc_167, \out_bs[7] [6], 
      \out_bs[7] [5], \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], uc_168, 
      uc_169}), .p_0(n_964));
   datapath__1_13941 i_0_674 (.to_int6126({uc_170, \out_bs[7] [6], 
      \out_bs[7] [5], \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], uc_171, 
      uc_172}), .p_0(n_965));
   datapath__1_13989 i_0_675 (.to_int6126({uc_173, \out_bs[7] [6], 
      \out_bs[7] [5], \out_bs[7] [4], \out_bs[7] [3], uc_174, uc_175, uc_176}), 
      .p_0(n_966));
   datapath__1_13957 i_0_676 (.to_int6126({uc_177, \out_bs[7] [6], 
      \out_bs[7] [5], \out_bs[7] [4], uc_178, uc_179, uc_180, uc_181}), .p_0(
      n_967));
   datapath__1_13829 i_0_677 (.to_int6126({uc_182, \out_bs[7] [6], 
      \out_bs[7] [5], \out_bs[7] [4], uc_183, uc_184, uc_185, uc_186}), .p_0(
      n_968));
   datapath__1_13638 i_0_678 (.to_int6126({uc_187, \out_bs[7] [6], 
      \out_bs[7] [5], uc_188, uc_189, uc_190, uc_191, uc_192}), .p_0(n_969));
   datapath__1_13765 i_0_679 (.to_int6128({1'b0, \out_as[7] [6], \out_as[7] [5], 
      \out_as[7] [4], \out_as[7] [3], \out_as[7] [2], \out_as[7] [1], 
      \out_as[7] [0]}), .p_0(n_970));
   OAI21_X1 i_0_680_0 (.A(n_0_680_0), .B1(n_0_680_3), .B2(n_0_680_1), .ZN(
      n_0_100));
   NAND2_X1 i_0_680_1 (.A1(n_99), .A2(n_0_680_1), .ZN(n_0_680_0));
   OAI22_X1 i_0_680_2 (.A1(n_952), .A2(n_508), .B1(n_0_680_2), .B2(n_507), 
      .ZN(n_0_680_1));
   INV_X1 i_0_680_3 (.A(n_952), .ZN(n_0_680_2));
   INV_X1 i_0_680_4 (.A(in_data[4]), .ZN(n_0_680_3));
   OAI21_X1 i_0_681_0 (.A(n_0_681_0), .B1(n_0_681_3), .B2(n_0_681_1), .ZN(
      n_0_101));
   NAND2_X1 i_0_681_1 (.A1(n_95), .A2(n_0_681_1), .ZN(n_0_681_0));
   OAI22_X1 i_0_681_2 (.A1(n_952), .A2(n_461), .B1(n_0_681_2), .B2(n_460), 
      .ZN(n_0_681_1));
   INV_X1 i_0_681_3 (.A(n_952), .ZN(n_0_681_2));
   INV_X1 i_0_681_4 (.A(in_data[4]), .ZN(n_0_681_3));
   AND2_X1 i_0_682_0 (.A1(n_772), .A2(n_953), .ZN(n_0_102));
   AND2_X1 i_0_683_0 (.A1(n_954), .A2(n_776), .ZN(n_0_103));
   AND2_X1 i_0_684_0 (.A1(n_839), .A2(n_955), .ZN(n_0_104));
   AND2_X1 i_0_685_0 (.A1(n_781), .A2(n_956), .ZN(n_0_105));
   AND2_X1 i_0_686_0 (.A1(n_793), .A2(n_957), .ZN(n_0_106));
   AND2_X1 i_0_687_0 (.A1(n_771), .A2(n_958), .ZN(n_0_107));
   AND2_X1 i_0_688_0 (.A1(n_779), .A2(n_959), .ZN(n_0_108));
   AND2_X1 i_0_689_0 (.A1(n_782), .A2(n_960), .ZN(n_0_109));
   AND2_X1 i_0_690_0 (.A1(n_790), .A2(n_961), .ZN(n_0_110));
   AND2_X1 i_0_691_0 (.A1(n_840), .A2(n_962), .ZN(n_0_111));
   AND2_X1 i_0_692_0 (.A1(n_773), .A2(n_963), .ZN(n_0_112));
   AND2_X1 i_0_693_0 (.A1(n_780), .A2(n_964), .ZN(n_0_113));
   AND2_X1 i_0_694_0 (.A1(n_788), .A2(n_965), .ZN(n_0_114));
   AND2_X1 i_0_695_0 (.A1(n_966), .A2(n_777), .ZN(n_0_115));
   AND2_X1 i_0_696_0 (.A1(n_784), .A2(n_967), .ZN(n_0_116));
   INV_X1 i_0_697_0 (.A(n_0_697_0), .ZN(n_0_117));
   NAND2_X1 i_0_697_1 (.A1(n_968), .A2(n_815), .ZN(n_0_697_0));
   AND2_X1 i_0_698_0 (.A1(n_709), .A2(n_969), .ZN(n_0_118));
   OAI21_X1 i_0_699_0 (.A(n_0_699_0), .B1(n_0_699_1), .B2(n_1310), .ZN(n_0_807));
   NAND2_X1 i_0_699_1 (.A1(n_1310), .A2(in_data[0]), .ZN(n_0_699_0));
   INV_X1 i_0_699_2 (.A(n_977), .ZN(n_0_699_1));
   INV_X1 i_0_700_0 (.A(n_0_700_0), .ZN(n_0_808));
   OAI21_X1 i_0_700_1 (.A(n_0_700_1), .B1(n_1125), .B2(n_0_126), .ZN(n_0_700_0));
   NAND2_X1 i_0_700_2 (.A1(n_0_126), .A2(n_0_700_2), .ZN(n_0_700_1));
   INV_X1 i_0_700_3 (.A(in_data[0]), .ZN(n_0_700_2));
   OAI21_X1 i_0_701_0 (.A(n_0_701_0), .B1(n_0_701_1), .B2(n_1287), .ZN(n_0_809));
   NAND2_X1 i_0_701_1 (.A1(n_1287), .A2(in_data[0]), .ZN(n_0_701_0));
   INV_X1 i_0_701_2 (.A(n_976), .ZN(n_0_701_1));
   OAI21_X1 i_0_702_0 (.A(n_0_702_0), .B1(n_0_702_1), .B2(n_1289), .ZN(n_0_810));
   NAND2_X1 i_0_702_1 (.A1(n_1289), .A2(in_data[0]), .ZN(n_0_702_0));
   INV_X1 i_0_702_2 (.A(n_975), .ZN(n_0_702_1));
   OAI21_X1 i_0_703_0 (.A(n_0_703_0), .B1(n_0_703_1), .B2(n_1281), .ZN(n_0_811));
   NAND2_X1 i_0_703_1 (.A1(n_1281), .A2(in_data[0]), .ZN(n_0_703_0));
   INV_X1 i_0_703_2 (.A(n_973), .ZN(n_0_703_1));
   OAI21_X1 i_0_704_0 (.A(n_0_704_0), .B1(n_0_704_1), .B2(n_1278), .ZN(n_0_812));
   NAND2_X1 i_0_704_1 (.A1(n_1278), .A2(in_data[0]), .ZN(n_0_704_0));
   INV_X1 i_0_704_2 (.A(n_972), .ZN(n_0_704_1));
   INV_X1 i_0_705_0 (.A(n_0_705_0), .ZN(n_0_813));
   OAI21_X1 i_0_705_1 (.A(n_0_705_1), .B1(n_1095), .B2(n_0_127), .ZN(n_0_705_0));
   NAND2_X1 i_0_705_2 (.A1(n_0_127), .A2(n_0_705_2), .ZN(n_0_705_1));
   INV_X1 i_0_705_3 (.A(in_data[0]), .ZN(n_0_705_2));
   INV_X1 i_0_706_0 (.A(n_0_706_0), .ZN(n_0_814));
   OAI21_X1 i_0_706_1 (.A(n_0_706_1), .B1(n_1094), .B2(n_0_125), .ZN(n_0_706_0));
   NAND2_X1 i_0_706_2 (.A1(n_0_125), .A2(n_0_706_2), .ZN(n_0_706_1));
   INV_X1 i_0_706_3 (.A(in_data[0]), .ZN(n_0_706_2));
   OAI21_X1 i_0_707_0 (.A(n_0_707_0), .B1(n_0_707_1), .B2(n_1275), .ZN(n_0_815));
   NAND2_X1 i_0_707_1 (.A1(n_1275), .A2(in_data[0]), .ZN(n_0_707_0));
   INV_X1 i_0_707_2 (.A(n_971), .ZN(n_0_707_1));
   OAI21_X1 i_0_708_0 (.A(n_0_708_0), .B1(n_0_708_3), .B2(n_0_708_1), .ZN(
      n_0_119));
   NAND2_X1 i_0_708_1 (.A1(n_126), .A2(n_0_708_1), .ZN(n_0_708_0));
   OAI22_X1 i_0_708_2 (.A1(n_952), .A2(n_1200), .B1(n_0_708_2), .B2(n_1199), 
      .ZN(n_0_708_1));
   INV_X1 i_0_708_3 (.A(n_952), .ZN(n_0_708_2));
   INV_X1 i_0_708_4 (.A(in_data[4]), .ZN(n_0_708_3));
   OAI21_X1 i_0_709_0 (.A(n_0_709_0), .B1(n_0_709_3), .B2(n_0_709_1), .ZN(n_971));
   NAND2_X1 i_0_709_1 (.A1(n_124), .A2(n_0_709_1), .ZN(n_0_709_0));
   OAI22_X1 i_0_709_2 (.A1(n_952), .A2(n_1308), .B1(n_0_709_2), .B2(n_1307), 
      .ZN(n_0_709_1));
   INV_X1 i_0_709_3 (.A(n_952), .ZN(n_0_709_2));
   INV_X1 i_0_709_4 (.A(in_data[4]), .ZN(n_0_709_3));
   OAI21_X1 i_0_710_0 (.A(n_0_710_0), .B1(n_0_710_3), .B2(n_0_710_1), .ZN(n_972));
   NAND2_X1 i_0_710_1 (.A1(n_120), .A2(n_0_710_1), .ZN(n_0_710_0));
   OAI22_X1 i_0_710_2 (.A1(n_952), .A2(n_1304), .B1(n_0_710_2), .B2(n_1303), 
      .ZN(n_0_710_1));
   INV_X1 i_0_710_3 (.A(n_952), .ZN(n_0_710_2));
   INV_X1 i_0_710_4 (.A(in_data[4]), .ZN(n_0_710_3));
   OAI21_X1 i_0_711_0 (.A(n_0_711_0), .B1(n_0_711_3), .B2(n_0_711_1), .ZN(n_973));
   NAND2_X1 i_0_711_1 (.A1(n_118), .A2(n_0_711_1), .ZN(n_0_711_0));
   OAI22_X1 i_0_711_2 (.A1(n_952), .A2(n_1302), .B1(n_0_711_2), .B2(n_1301), 
      .ZN(n_0_711_1));
   INV_X1 i_0_711_3 (.A(n_952), .ZN(n_0_711_2));
   INV_X1 i_0_711_4 (.A(in_data[4]), .ZN(n_0_711_3));
   OAI21_X1 i_0_712_0 (.A(n_0_712_0), .B1(n_0_712_3), .B2(n_0_712_1), .ZN(n_974));
   NAND2_X1 i_0_712_1 (.A1(n_117), .A2(n_0_712_1), .ZN(n_0_712_0));
   OAI22_X1 i_0_712_2 (.A1(n_952), .A2(n_1202), .B1(n_0_712_2), .B2(n_1201), 
      .ZN(n_0_712_1));
   INV_X1 i_0_712_3 (.A(n_952), .ZN(n_0_712_2));
   INV_X1 i_0_712_4 (.A(in_data[4]), .ZN(n_0_712_3));
   OAI21_X1 i_0_713_0 (.A(n_0_713_0), .B1(n_0_713_3), .B2(n_0_713_1), .ZN(n_975));
   NAND2_X1 i_0_713_1 (.A1(n_115), .A2(n_0_713_1), .ZN(n_0_713_0));
   OAI22_X1 i_0_713_2 (.A1(n_952), .A2(n_1298), .B1(n_0_713_2), .B2(n_1297), 
      .ZN(n_0_713_1));
   INV_X1 i_0_713_3 (.A(n_952), .ZN(n_0_713_2));
   INV_X1 i_0_713_4 (.A(in_data[4]), .ZN(n_0_713_3));
   OAI21_X1 i_0_714_0 (.A(n_0_714_0), .B1(n_0_714_3), .B2(n_0_714_1), .ZN(n_976));
   NAND2_X1 i_0_714_1 (.A1(n_107), .A2(n_0_714_1), .ZN(n_0_714_0));
   OAI22_X1 i_0_714_2 (.A1(n_952), .A2(n_1292), .B1(n_0_714_2), .B2(n_1291), 
      .ZN(n_0_714_1));
   INV_X1 i_0_714_3 (.A(n_952), .ZN(n_0_714_2));
   INV_X1 i_0_714_4 (.A(in_data[4]), .ZN(n_0_714_3));
   OAI21_X1 i_0_715_0 (.A(n_0_715_0), .B1(n_0_715_3), .B2(n_0_715_1), .ZN(
      n_0_900));
   NAND2_X1 i_0_715_1 (.A1(n_1197), .A2(n_0_715_1), .ZN(n_0_715_0));
   OAI22_X1 i_0_715_2 (.A1(n_952), .A2(n_1209), .B1(n_0_715_2), .B2(n_1208), 
      .ZN(n_0_715_1));
   INV_X1 i_0_715_3 (.A(n_952), .ZN(n_0_715_2));
   INV_X1 i_0_715_4 (.A(in_data[4]), .ZN(n_0_715_3));
   OAI21_X1 i_0_716_0 (.A(n_0_716_0), .B1(n_0_716_3), .B2(n_0_716_1), .ZN(
      n_0_899));
   NAND2_X1 i_0_716_1 (.A1(n_1090), .A2(n_0_716_1), .ZN(n_0_716_0));
   OAI22_X1 i_0_716_2 (.A1(n_952), .A2(n_1207), .B1(n_0_716_2), .B2(n_1206), 
      .ZN(n_0_716_1));
   INV_X1 i_0_716_3 (.A(n_952), .ZN(n_0_716_2));
   INV_X1 i_0_716_4 (.A(in_data[4]), .ZN(n_0_716_3));
   OAI21_X1 i_0_717_0 (.A(n_0_717_0), .B1(n_0_717_3), .B2(n_0_717_1), .ZN(
      n_0_898));
   NAND2_X1 i_0_717_1 (.A1(n_1195), .A2(n_0_717_1), .ZN(n_0_717_0));
   OAI22_X1 i_0_717_2 (.A1(n_952), .A2(n_1205), .B1(n_0_717_2), .B2(n_1204), 
      .ZN(n_0_717_1));
   INV_X1 i_0_717_3 (.A(n_952), .ZN(n_0_717_2));
   INV_X1 i_0_717_4 (.A(in_data[4]), .ZN(n_0_717_3));
   OAI21_X1 i_0_718_0 (.A(n_0_718_0), .B1(n_0_718_3), .B2(n_0_718_1), .ZN(
      n_0_897));
   NAND2_X1 i_0_718_1 (.A1(n_1193), .A2(n_0_718_1), .ZN(n_0_718_0));
   OAI22_X1 i_0_718_2 (.A1(n_952), .A2(n_465), .B1(n_0_718_2), .B2(n_1203), 
      .ZN(n_0_718_1));
   INV_X1 i_0_718_3 (.A(n_952), .ZN(n_0_718_2));
   INV_X1 i_0_718_4 (.A(in_data[4]), .ZN(n_0_718_3));
   OAI21_X1 i_0_719_0 (.A(n_0_719_0), .B1(n_0_719_3), .B2(n_0_719_1), .ZN(
      n_0_896));
   NAND2_X1 i_0_719_1 (.A1(n_1192), .A2(n_0_719_1), .ZN(n_0_719_0));
   OAI22_X1 i_0_719_2 (.A1(n_952), .A2(n_1294), .B1(n_0_719_2), .B2(n_1293), 
      .ZN(n_0_719_1));
   INV_X1 i_0_719_3 (.A(n_952), .ZN(n_0_719_2));
   INV_X1 i_0_719_4 (.A(in_data[4]), .ZN(n_0_719_3));
   OAI21_X1 i_0_720_0 (.A(n_0_720_0), .B1(n_0_720_3), .B2(n_0_720_1), .ZN(n_977));
   NAND2_X1 i_0_720_1 (.A1(n_1191), .A2(n_0_720_1), .ZN(n_0_720_0));
   OAI22_X1 i_0_720_2 (.A1(n_952), .A2(n_1296), .B1(n_0_720_2), .B2(n_1295), 
      .ZN(n_0_720_1));
   INV_X1 i_0_720_3 (.A(n_952), .ZN(n_0_720_2));
   INV_X1 i_0_720_4 (.A(in_data[4]), .ZN(n_0_720_3));
   OAI21_X1 i_0_721_0 (.A(n_0_721_0), .B1(n_0_721_3), .B2(n_0_721_1), .ZN(
      n_0_895));
   NAND2_X1 i_0_721_1 (.A1(n_1190), .A2(n_0_721_1), .ZN(n_0_721_0));
   OAI22_X1 i_0_721_2 (.A1(n_952), .A2(n_1300), .B1(n_0_721_2), .B2(n_1299), 
      .ZN(n_0_721_1));
   INV_X1 i_0_721_3 (.A(n_952), .ZN(n_0_721_2));
   INV_X1 i_0_721_4 (.A(in_data[4]), .ZN(n_0_721_3));
   OAI21_X1 i_0_722_0 (.A(n_0_722_0), .B1(n_0_722_3), .B2(n_0_722_1), .ZN(
      n_0_120));
   NAND2_X1 i_0_722_1 (.A1(n_1194), .A2(n_0_722_1), .ZN(n_0_722_0));
   OAI22_X1 i_0_722_2 (.A1(n_952), .A2(n_387), .B1(n_0_722_2), .B2(n_386), 
      .ZN(n_0_722_1));
   INV_X1 i_0_722_3 (.A(n_952), .ZN(n_0_722_2));
   INV_X1 i_0_722_4 (.A(in_data[4]), .ZN(n_0_722_3));
   OAI21_X1 i_0_723_0 (.A(n_0_723_0), .B1(n_0_723_3), .B2(n_0_723_1), .ZN(
      n_0_121));
   NAND2_X1 i_0_723_1 (.A1(n_1196), .A2(n_0_723_1), .ZN(n_0_723_0));
   OAI22_X1 i_0_723_2 (.A1(n_952), .A2(n_262), .B1(n_0_723_2), .B2(n_261), 
      .ZN(n_0_723_1));
   INV_X1 i_0_723_3 (.A(n_952), .ZN(n_0_723_2));
   INV_X1 i_0_723_4 (.A(in_data[4]), .ZN(n_0_723_3));
   OAI21_X1 i_0_724_0 (.A(n_0_724_0), .B1(n_0_724_3), .B2(n_0_724_1), .ZN(
      n_0_122));
   NAND2_X1 i_0_724_1 (.A1(n_84), .A2(n_0_724_1), .ZN(n_0_724_0));
   OAI22_X1 i_0_724_2 (.A1(n_952), .A2(n_407), .B1(n_0_724_2), .B2(n_406), 
      .ZN(n_0_724_1));
   INV_X1 i_0_724_3 (.A(n_952), .ZN(n_0_724_2));
   INV_X1 i_0_724_4 (.A(in_data[4]), .ZN(n_0_724_3));
   OAI21_X1 i_0_725_0 (.A(n_0_725_0), .B1(n_0_725_3), .B2(n_0_725_1), .ZN(
      n_0_123));
   NAND2_X1 i_0_725_1 (.A1(n_101), .A2(n_0_725_1), .ZN(n_0_725_0));
   OAI22_X1 i_0_725_2 (.A1(n_952), .A2(n_523), .B1(n_0_725_2), .B2(n_522), 
      .ZN(n_0_725_1));
   INV_X1 i_0_725_3 (.A(n_952), .ZN(n_0_725_2));
   INV_X1 i_0_725_4 (.A(in_data[4]), .ZN(n_0_725_3));
   OAI21_X1 i_0_726_0 (.A(n_0_726_0), .B1(n_0_726_3), .B2(n_0_726_1), .ZN(
      n_0_124));
   NAND2_X1 i_0_726_1 (.A1(n_102), .A2(n_0_726_1), .ZN(n_0_726_0));
   OAI22_X1 i_0_726_2 (.A1(n_952), .A2(n_528), .B1(n_0_726_2), .B2(n_527), 
      .ZN(n_0_726_1));
   INV_X1 i_0_726_3 (.A(n_952), .ZN(n_0_726_2));
   INV_X1 i_0_726_4 (.A(in_data[4]), .ZN(n_0_726_3));
   AND2_X1 i_0_727_0 (.A1(n_735), .A2(n_0_403), .ZN(n_0_125));
   AND2_X1 i_0_728_0 (.A1(n_678), .A2(n_0_544), .ZN(n_0_126));
   AND2_X1 i_0_729_0 (.A1(n_731), .A2(n_0_404), .ZN(n_0_127));
   DFF_X1 \buf_reg[14]  (.D(n_0_936), .CK(clk), .Q(n_978), .QN());
   DFF_X1 \buf_reg[28]  (.D(n_0_922), .CK(clk), .Q(n_979), .QN());
   DFF_X1 \buf_reg[39]  (.D(n_0_911), .CK(clk), .Q(n_980), .QN());
   DFF_X1 \buf_reg[64]  (.D(n_0_879), .CK(clk), .Q(n_981), .QN());
   DFF_X1 \buf_reg[91]  (.D(n_0_852), .CK(clk), .Q(n_982), .QN());
   DFF_X1 \buf_reg[95]  (.D(n_0_848), .CK(clk), .Q(n_983), .QN());
   DFF_X1 \buf_reg[109]  (.D(n_0_834), .CK(clk), .Q(n_984), .QN());
   DFF_X1 \buf_reg[122]  (.D(n_0_821), .CK(clk), .Q(n_985), .QN());
   DFF_X1 \buf_reg[123]  (.D(n_0_820), .CK(clk), .Q(n_986), .QN());
   INV_X1 i_0_657_0 (.A(n_0_657_1), .ZN(n_0_657_0));
   NAND2_X1 i_0_657_1 (.A1(n_0_253), .A2(n_0_657_964), .ZN(n_0_657_1));
   INV_X1 i_0_657_2 (.A(n_0_657_3), .ZN(n_0_657_2));
   NAND2_X1 i_0_657_3 (.A1(n_0_232), .A2(n_0_657_964), .ZN(n_0_657_3));
   OAI21_X1 i_0_657_4 (.A(n_0_657_4), .B1(n_0_806), .B2(n_0_657_7), .ZN(n_0_848));
   OAI221_X1 i_0_657_5 (.A(n_0_806), .B1(n_983), .B2(n_0_657_5), .C1(n_0_635), 
      .C2(n_0_657_6), .ZN(n_0_657_4));
   INV_X1 i_0_657_6 (.A(n_0_657_6), .ZN(n_0_657_5));
   NAND2_X1 i_0_657_7 (.A1(n_0_226), .A2(n_0_657_964), .ZN(n_0_657_6));
   AOI22_X1 i_0_657_8 (.A1(n_983), .A2(n_0_657_9), .B1(n_0_349), .B2(n_0_657_8), 
      .ZN(n_0_657_7));
   INV_X1 i_0_657_9 (.A(n_0_657_9), .ZN(n_0_657_8));
   NAND2_X1 i_0_657_10 (.A1(n_0_774), .A2(n_0_657_964), .ZN(n_0_657_9));
   INV_X1 i_0_657_11 (.A(n_0_657_11), .ZN(n_0_657_10));
   NAND2_X1 i_0_657_12 (.A1(n_0_208), .A2(n_0_657_964), .ZN(n_0_657_11));
   INV_X1 i_0_657_13 (.A(n_0_657_13), .ZN(n_0_657_12));
   NAND2_X1 i_0_657_14 (.A1(n_0_202), .A2(n_0_657_964), .ZN(n_0_657_13));
   INV_X1 i_0_657_15 (.A(n_0_657_15), .ZN(n_0_657_14));
   NAND2_X1 i_0_657_16 (.A1(n_0_201), .A2(n_0_657_964), .ZN(n_0_657_15));
   INV_X1 i_0_657_17 (.A(n_0_657_17), .ZN(n_0_657_16));
   NAND2_X1 i_0_657_18 (.A1(n_0_200), .A2(n_0_657_964), .ZN(n_0_657_17));
   INV_X1 i_0_657_19 (.A(n_0_657_19), .ZN(n_0_657_18));
   NAND2_X1 i_0_657_20 (.A1(n_0_198), .A2(n_0_657_964), .ZN(n_0_657_19));
   INV_X1 i_0_657_21 (.A(n_0_657_21), .ZN(n_0_657_20));
   NAND2_X1 i_0_657_22 (.A1(n_0_196), .A2(n_0_657_964), .ZN(n_0_657_21));
   OAI21_X1 i_0_657_23 (.A(n_0_657_22), .B1(n_0_806), .B2(n_0_657_25), .ZN(
      n_0_879));
   OAI221_X1 i_0_657_24 (.A(n_0_806), .B1(n_981), .B2(n_0_657_23), .C1(n_0_262), 
      .C2(n_0_657_24), .ZN(n_0_657_22));
   INV_X1 i_0_657_25 (.A(n_0_657_24), .ZN(n_0_657_23));
   NAND2_X1 i_0_657_26 (.A1(n_0_195), .A2(n_0_657_964), .ZN(n_0_657_24));
   AOI22_X1 i_0_657_27 (.A1(n_981), .A2(n_0_657_27), .B1(n_0_318), .B2(
      n_0_657_26), .ZN(n_0_657_25));
   INV_X1 i_0_657_28 (.A(n_0_657_27), .ZN(n_0_657_26));
   NAND2_X1 i_0_657_29 (.A1(n_0_743), .A2(n_0_657_964), .ZN(n_0_657_27));
   OAI21_X1 i_0_657_30 (.A(n_0_657_28), .B1(n_0_806), .B2(n_0_657_31), .ZN(
      n_0_911));
   OAI221_X1 i_0_657_31 (.A(n_0_806), .B1(n_980), .B2(n_0_657_29), .C1(n_0_428), 
      .C2(n_0_657_30), .ZN(n_0_657_28));
   INV_X1 i_0_657_32 (.A(n_0_657_30), .ZN(n_0_657_29));
   NAND2_X1 i_0_657_33 (.A1(n_0_170), .A2(n_0_657_964), .ZN(n_0_657_30));
   AOI22_X1 i_0_657_34 (.A1(n_980), .A2(n_0_657_33), .B1(n_0_293), .B2(
      n_0_657_32), .ZN(n_0_657_31));
   INV_X1 i_0_657_35 (.A(n_0_657_33), .ZN(n_0_657_32));
   NAND2_X1 i_0_657_36 (.A1(n_0_719), .A2(n_0_657_964), .ZN(n_0_657_33));
   OAI21_X1 i_0_657_37 (.A(n_0_657_34), .B1(n_0_806), .B2(n_0_657_37), .ZN(
      n_0_920));
   OAI221_X1 i_0_657_38 (.A(n_0_806), .B1(n_924), .B2(n_0_657_35), .C1(n_0_809), 
      .C2(n_0_657_36), .ZN(n_0_657_34));
   INV_X1 i_0_657_39 (.A(n_0_657_36), .ZN(n_0_657_35));
   NAND2_X1 i_0_657_40 (.A1(n_0_161), .A2(n_0_657_964), .ZN(n_0_657_36));
   AOI22_X1 i_0_657_41 (.A1(n_924), .A2(n_0_657_39), .B1(n_1286), .B2(n_0_657_38), 
      .ZN(n_0_657_37));
   INV_X1 i_0_657_42 (.A(n_0_657_39), .ZN(n_0_657_38));
   NAND2_X1 i_0_657_43 (.A1(n_1285), .A2(n_0_657_964), .ZN(n_0_657_39));
   OAI21_X1 i_0_657_44 (.A(n_0_657_40), .B1(n_0_806), .B2(n_0_657_43), .ZN(
      n_0_922));
   OAI221_X1 i_0_657_45 (.A(n_0_806), .B1(n_979), .B2(n_0_657_41), .C1(n_0_670), 
      .C2(n_0_657_42), .ZN(n_0_657_40));
   INV_X1 i_0_657_46 (.A(n_0_657_42), .ZN(n_0_657_41));
   NAND2_X1 i_0_657_47 (.A1(n_0_159), .A2(n_0_657_964), .ZN(n_0_657_42));
   AOI22_X1 i_0_657_48 (.A1(n_979), .A2(n_0_657_45), .B1(n_0_283), .B2(
      n_0_657_44), .ZN(n_0_657_43));
   INV_X1 i_0_657_49 (.A(n_0_657_45), .ZN(n_0_657_44));
   NAND2_X1 i_0_657_50 (.A1(n_0_705), .A2(n_0_657_964), .ZN(n_0_657_45));
   OAI21_X1 i_0_657_51 (.A(n_0_657_46), .B1(n_0_806), .B2(n_0_657_49), .ZN(
      n_0_934));
   OAI221_X1 i_0_657_52 (.A(n_0_806), .B1(n_937), .B2(n_0_657_47), .C1(n_0_807), 
      .C2(n_0_657_48), .ZN(n_0_657_46));
   INV_X1 i_0_657_53 (.A(n_0_657_48), .ZN(n_0_657_47));
   NAND2_X1 i_0_657_54 (.A1(n_0_147), .A2(n_0_657_964), .ZN(n_0_657_48));
   AOI22_X1 i_0_657_55 (.A1(n_937), .A2(n_0_657_51), .B1(n_1284), .B2(n_0_657_50), 
      .ZN(n_0_657_49));
   INV_X1 i_0_657_56 (.A(n_0_657_51), .ZN(n_0_657_50));
   NAND2_X1 i_0_657_57 (.A1(n_1283), .A2(n_0_657_964), .ZN(n_0_657_51));
   INV_X1 i_0_657_58 (.A(n_0_657_53), .ZN(n_0_657_52));
   NAND2_X1 i_0_657_59 (.A1(n_0_146), .A2(n_0_657_964), .ZN(n_0_657_53));
   INV_X1 i_0_657_60 (.A(n_0_657_55), .ZN(n_0_657_54));
   NAND2_X1 i_0_657_61 (.A1(n_0_143), .A2(n_0_657_964), .ZN(n_0_657_55));
   OAI21_X1 i_0_657_62 (.A(n_0_657_56), .B1(n_0_806), .B2(n_0_657_59), .ZN(
      n_0_939));
   OAI221_X1 i_0_657_63 (.A(n_0_806), .B1(n_940), .B2(n_0_657_57), .C1(n_0_811), 
      .C2(n_0_657_58), .ZN(n_0_657_56));
   INV_X1 i_0_657_64 (.A(n_0_657_58), .ZN(n_0_657_57));
   NAND2_X1 i_0_657_65 (.A1(n_0_142), .A2(n_0_657_964), .ZN(n_0_657_58));
   AOI22_X1 i_0_657_66 (.A1(n_940), .A2(n_0_657_61), .B1(n_1280), .B2(n_0_657_60), 
      .ZN(n_0_657_59));
   INV_X1 i_0_657_67 (.A(n_0_657_61), .ZN(n_0_657_60));
   NAND2_X1 i_0_657_68 (.A1(n_1279), .A2(n_0_657_964), .ZN(n_0_657_61));
   OAI21_X1 i_0_657_69 (.A(n_0_657_62), .B1(n_0_806), .B2(n_0_657_65), .ZN(
      n_0_941));
   OAI221_X1 i_0_657_70 (.A(n_0_806), .B1(n_942), .B2(n_0_657_63), .C1(n_0_812), 
      .C2(n_0_657_64), .ZN(n_0_657_62));
   INV_X1 i_0_657_71 (.A(n_0_657_64), .ZN(n_0_657_63));
   NAND2_X1 i_0_657_72 (.A1(n_0_140), .A2(n_0_657_964), .ZN(n_0_657_64));
   AOI22_X1 i_0_657_73 (.A1(n_942), .A2(n_0_657_67), .B1(n_1277), .B2(n_0_657_66), 
      .ZN(n_0_657_65));
   INV_X1 i_0_657_74 (.A(n_0_657_67), .ZN(n_0_657_66));
   NAND2_X1 i_0_657_75 (.A1(n_1276), .A2(n_0_657_964), .ZN(n_0_657_67));
   OAI21_X1 i_0_657_76 (.A(n_0_657_68), .B1(n_0_806), .B2(n_0_657_71), .ZN(
      n_0_945));
   OAI221_X1 i_0_657_77 (.A(n_0_806), .B1(n_946), .B2(n_0_657_69), .C1(n_0_815), 
      .C2(n_0_657_70), .ZN(n_0_657_68));
   INV_X1 i_0_657_78 (.A(n_0_657_70), .ZN(n_0_657_69));
   NAND2_X1 i_0_657_79 (.A1(n_0_136), .A2(n_0_657_964), .ZN(n_0_657_70));
   AOI22_X1 i_0_657_80 (.A1(n_946), .A2(n_0_657_73), .B1(n_1274), .B2(n_0_657_72), 
      .ZN(n_0_657_71));
   INV_X1 i_0_657_81 (.A(n_0_657_73), .ZN(n_0_657_72));
   NAND2_X1 i_0_657_82 (.A1(n_1273), .A2(n_0_657_964), .ZN(n_0_657_73));
   INV_X1 i_0_657_83 (.A(n_0_657_75), .ZN(n_0_657_74));
   NAND2_X1 i_0_657_84 (.A1(n_0_682), .A2(n_0_657_964), .ZN(n_0_657_75));
   OAI33_X1 i_0_657_85 (.A1(n_0_806), .A2(n_0_657_813), .A3(n_0_657_80), 
      .B1(n_0_657_87), .B2(n_0_657_76), .B3(n_0_657_77), .ZN(n_0_950));
   AOI21_X1 i_0_657_86 (.A(n_950), .B1(n_0_131), .B2(n_0_657_964), .ZN(
      n_0_657_76));
   NOR3_X1 i_0_657_87 (.A1(n_0_657_79), .A2(n_0_657_813), .A3(n_1268), .ZN(
      n_0_657_77));
   INV_X1 i_0_657_88 (.A(enbl_in), .ZN(n_0_657_78));
   INV_X1 i_0_657_89 (.A(n_0_131), .ZN(n_0_657_79));
   INV_X1 i_0_657_90 (.A(in_data[0]), .ZN(n_0_657_80));
   OAI21_X1 i_0_657_91 (.A(n_0_657_81), .B1(n_0_657_82), .B2(n_0_657_87), 
      .ZN(n_0_816));
   NAND2_X1 i_0_657_92 (.A1(n_0_657_87), .A2(in_data[0]), .ZN(n_0_657_81));
   AOI21_X1 i_0_657_93 (.A(n_0_657_83), .B1(n_0_261), .B2(n_0_657_85), .ZN(
      n_0_657_82));
   AOI21_X1 i_0_657_94 (.A(n_0_657_84), .B1(n_0_258), .B2(n_0_657_964), .ZN(
      n_0_657_83));
   INV_X1 i_0_657_95 (.A(n_857), .ZN(n_0_657_84));
   INV_X1 i_0_657_96 (.A(n_0_657_86), .ZN(n_0_657_85));
   NAND2_X1 i_0_657_97 (.A1(n_0_258), .A2(n_0_657_964), .ZN(n_0_657_86));
   NOR2_X1 i_0_657_98 (.A1(n_0_806), .A2(n_0_657_813), .ZN(n_0_657_87));
   NAND2_X1 i_0_657_99 (.A1(n_0_657_91), .A2(n_0_657_88), .ZN(n_0_817));
   OAI21_X1 i_0_657_100 (.A(n_0_657_89), .B1(n_0_380), .B2(n_0_657_90), .ZN(
      n_0_657_88));
   AOI21_X1 i_0_657_101 (.A(n_0_806), .B1(n_0_657_90), .B2(n_0_657_93), .ZN(
      n_0_657_89));
   NAND2_X1 i_0_657_102 (.A1(n_0_805), .A2(n_0_657_964), .ZN(n_0_657_90));
   OAI21_X1 i_0_657_103 (.A(n_0_657_92), .B1(n_0_599), .B2(n_0_657_94), .ZN(
      n_0_657_91));
   AOI21_X1 i_0_657_104 (.A(n_0_657_959), .B1(n_0_657_94), .B2(n_0_657_93), 
      .ZN(n_0_657_92));
   INV_X1 i_0_657_105 (.A(n_858), .ZN(n_0_657_93));
   NAND2_X1 i_0_657_106 (.A1(n_0_257), .A2(n_0_657_964), .ZN(n_0_657_94));
   NAND2_X1 i_0_657_107 (.A1(n_0_657_95), .A2(n_0_657_98), .ZN(n_0_818));
   OAI21_X1 i_0_657_108 (.A(n_0_657_96), .B1(n_0_379), .B2(n_0_657_97), .ZN(
      n_0_657_95));
   AOI21_X1 i_0_657_109 (.A(n_0_806), .B1(n_0_657_97), .B2(n_0_657_100), 
      .ZN(n_0_657_96));
   NAND2_X1 i_0_657_110 (.A1(n_0_804), .A2(n_0_657_964), .ZN(n_0_657_97));
   OAI21_X1 i_0_657_111 (.A(n_0_657_99), .B1(n_0_596), .B2(n_0_657_101), 
      .ZN(n_0_657_98));
   AOI21_X1 i_0_657_112 (.A(n_0_657_959), .B1(n_0_657_101), .B2(n_0_657_100), 
      .ZN(n_0_657_99));
   INV_X1 i_0_657_113 (.A(n_859), .ZN(n_0_657_100));
   NAND2_X1 i_0_657_114 (.A1(n_0_256), .A2(n_0_657_964), .ZN(n_0_657_101));
   NAND2_X1 i_0_657_115 (.A1(n_0_657_102), .A2(n_0_657_105), .ZN(n_0_819));
   OAI21_X1 i_0_657_116 (.A(n_0_657_103), .B1(n_0_378), .B2(n_0_657_104), 
      .ZN(n_0_657_102));
   AOI21_X1 i_0_657_117 (.A(n_0_806), .B1(n_0_657_104), .B2(n_0_657_107), 
      .ZN(n_0_657_103));
   NAND2_X1 i_0_657_118 (.A1(n_0_803), .A2(n_0_657_964), .ZN(n_0_657_104));
   OAI21_X1 i_0_657_119 (.A(n_0_657_106), .B1(n_0_595), .B2(n_0_657_108), 
      .ZN(n_0_657_105));
   AOI21_X1 i_0_657_120 (.A(n_0_657_959), .B1(n_0_657_108), .B2(n_0_657_107), 
      .ZN(n_0_657_106));
   INV_X1 i_0_657_121 (.A(n_860), .ZN(n_0_657_107));
   NAND2_X1 i_0_657_122 (.A1(n_0_255), .A2(n_0_657_964), .ZN(n_0_657_108));
   NAND2_X1 i_0_657_123 (.A1(n_0_657_109), .A2(n_0_657_112), .ZN(n_0_820));
   OAI21_X1 i_0_657_124 (.A(n_0_657_110), .B1(n_0_377), .B2(n_0_657_111), 
      .ZN(n_0_657_109));
   AOI21_X1 i_0_657_125 (.A(n_0_806), .B1(n_0_657_111), .B2(n_0_657_114), 
      .ZN(n_0_657_110));
   NAND2_X1 i_0_657_126 (.A1(n_0_802), .A2(n_0_657_964), .ZN(n_0_657_111));
   OAI211_X1 i_0_657_127 (.A(n_0_657_113), .B(n_0_806), .C1(n_0_602), .C2(
      n_0_657_115), .ZN(n_0_657_112));
   NAND2_X1 i_0_657_128 (.A1(n_0_657_115), .A2(n_0_657_114), .ZN(n_0_657_113));
   INV_X1 i_0_657_129 (.A(n_986), .ZN(n_0_657_114));
   NAND2_X1 i_0_657_130 (.A1(n_0_254), .A2(n_0_657_964), .ZN(n_0_657_115));
   OAI21_X1 i_0_657_131 (.A(n_0_657_118), .B1(n_0_657_117), .B2(n_0_657_116), 
      .ZN(n_0_821));
   OAI21_X1 i_0_657_132 (.A(n_0_806), .B1(n_0_657_0), .B2(n_985), .ZN(
      n_0_657_116));
   NOR2_X1 i_0_657_133 (.A1(n_0_605), .A2(n_0_657_1), .ZN(n_0_657_117));
   OAI21_X1 i_0_657_134 (.A(n_0_657_119), .B1(n_0_376), .B2(n_0_657_121), 
      .ZN(n_0_657_118));
   AOI21_X1 i_0_657_135 (.A(n_0_806), .B1(n_0_657_121), .B2(n_0_657_120), 
      .ZN(n_0_657_119));
   INV_X1 i_0_657_136 (.A(n_985), .ZN(n_0_657_120));
   NAND2_X1 i_0_657_137 (.A1(n_0_801), .A2(n_0_657_964), .ZN(n_0_657_121));
   NAND2_X1 i_0_657_138 (.A1(n_0_657_122), .A2(n_0_657_125), .ZN(n_0_822));
   OAI21_X1 i_0_657_139 (.A(n_0_657_123), .B1(n_0_375), .B2(n_0_657_124), 
      .ZN(n_0_657_122));
   AOI21_X1 i_0_657_140 (.A(n_0_806), .B1(n_0_657_124), .B2(n_0_657_127), 
      .ZN(n_0_657_123));
   NAND2_X1 i_0_657_141 (.A1(n_0_800), .A2(n_0_657_964), .ZN(n_0_657_124));
   OAI21_X1 i_0_657_142 (.A(n_0_657_126), .B1(n_0_594), .B2(n_0_657_128), 
      .ZN(n_0_657_125));
   AOI21_X1 i_0_657_143 (.A(n_0_657_959), .B1(n_0_657_128), .B2(n_0_657_127), 
      .ZN(n_0_657_126));
   INV_X1 i_0_657_144 (.A(n_861), .ZN(n_0_657_127));
   NAND2_X1 i_0_657_145 (.A1(n_0_252), .A2(n_0_657_964), .ZN(n_0_657_128));
   NAND2_X1 i_0_657_146 (.A1(n_0_657_129), .A2(n_0_657_132), .ZN(n_0_823));
   OAI21_X1 i_0_657_147 (.A(n_0_657_130), .B1(n_0_374), .B2(n_0_657_131), 
      .ZN(n_0_657_129));
   AOI21_X1 i_0_657_148 (.A(n_0_806), .B1(n_0_657_131), .B2(n_0_657_134), 
      .ZN(n_0_657_130));
   NAND2_X1 i_0_657_149 (.A1(n_0_799), .A2(n_0_657_964), .ZN(n_0_657_131));
   OAI21_X1 i_0_657_150 (.A(n_0_657_133), .B1(n_0_591), .B2(n_0_657_135), 
      .ZN(n_0_657_132));
   AOI21_X1 i_0_657_151 (.A(n_0_657_959), .B1(n_0_657_135), .B2(n_0_657_134), 
      .ZN(n_0_657_133));
   INV_X1 i_0_657_152 (.A(n_862), .ZN(n_0_657_134));
   NAND2_X1 i_0_657_153 (.A1(n_0_251), .A2(n_0_657_964), .ZN(n_0_657_135));
   NAND2_X1 i_0_657_154 (.A1(n_0_657_136), .A2(n_0_657_139), .ZN(n_0_824));
   OAI21_X1 i_0_657_155 (.A(n_0_657_137), .B1(n_0_373), .B2(n_0_657_138), 
      .ZN(n_0_657_136));
   AOI21_X1 i_0_657_156 (.A(n_0_806), .B1(n_0_657_138), .B2(n_0_657_141), 
      .ZN(n_0_657_137));
   NAND2_X1 i_0_657_157 (.A1(n_0_798), .A2(n_0_657_964), .ZN(n_0_657_138));
   OAI21_X1 i_0_657_158 (.A(n_0_657_140), .B1(n_0_608), .B2(n_0_657_142), 
      .ZN(n_0_657_139));
   AOI21_X1 i_0_657_159 (.A(n_0_657_959), .B1(n_0_657_141), .B2(n_0_657_142), 
      .ZN(n_0_657_140));
   INV_X1 i_0_657_160 (.A(n_863), .ZN(n_0_657_141));
   NAND2_X1 i_0_657_161 (.A1(n_0_250), .A2(n_0_657_964), .ZN(n_0_657_142));
   OAI21_X1 i_0_657_162 (.A(n_0_657_147), .B1(n_0_657_143), .B2(n_0_657_145), 
      .ZN(n_0_825));
   OAI21_X1 i_0_657_163 (.A(n_0_657_959), .B1(n_0_657_144), .B2(n_987), .ZN(
      n_0_657_143));
   INV_X1 i_0_657_164 (.A(n_0_657_146), .ZN(n_0_657_144));
   NOR2_X1 i_0_657_165 (.A1(n_0_372), .A2(n_0_657_146), .ZN(n_0_657_145));
   NAND2_X1 i_0_657_166 (.A1(n_0_797), .A2(n_0_657_964), .ZN(n_0_657_146));
   OAI21_X1 i_0_657_167 (.A(n_0_657_148), .B1(n_0_588), .B2(n_0_657_150), 
      .ZN(n_0_657_147));
   AOI21_X1 i_0_657_168 (.A(n_0_657_959), .B1(n_0_657_150), .B2(n_0_657_149), 
      .ZN(n_0_657_148));
   INV_X1 i_0_657_169 (.A(n_987), .ZN(n_0_657_149));
   NAND2_X1 i_0_657_170 (.A1(n_0_249), .A2(n_0_657_964), .ZN(n_0_657_150));
   NAND2_X1 i_0_657_171 (.A1(n_0_657_151), .A2(n_0_657_154), .ZN(n_0_826));
   OAI21_X1 i_0_657_172 (.A(n_0_657_152), .B1(n_0_371), .B2(n_0_657_153), 
      .ZN(n_0_657_151));
   AOI21_X1 i_0_657_173 (.A(n_0_806), .B1(n_0_657_153), .B2(n_0_657_156), 
      .ZN(n_0_657_152));
   NAND2_X1 i_0_657_174 (.A1(n_0_796), .A2(n_0_657_964), .ZN(n_0_657_153));
   OAI211_X1 i_0_657_175 (.A(n_0_657_155), .B(n_0_806), .C1(n_0_585), .C2(
      n_0_657_157), .ZN(n_0_657_154));
   NAND2_X1 i_0_657_176 (.A1(n_0_657_157), .A2(n_0_657_156), .ZN(n_0_657_155));
   INV_X1 i_0_657_177 (.A(n_864), .ZN(n_0_657_156));
   NAND2_X1 i_0_657_178 (.A1(n_0_248), .A2(n_0_657_964), .ZN(n_0_657_157));
   NAND2_X1 i_0_657_179 (.A1(n_0_657_158), .A2(n_0_657_161), .ZN(n_0_827));
   OAI21_X1 i_0_657_180 (.A(n_0_657_159), .B1(n_0_370), .B2(n_0_657_160), 
      .ZN(n_0_657_158));
   AOI21_X1 i_0_657_181 (.A(n_0_806), .B1(n_0_657_160), .B2(n_0_657_163), 
      .ZN(n_0_657_159));
   NAND2_X1 i_0_657_182 (.A1(n_0_795), .A2(n_0_657_964), .ZN(n_0_657_160));
   OAI21_X1 i_0_657_183 (.A(n_0_657_162), .B1(n_0_582), .B2(n_0_657_164), 
      .ZN(n_0_657_161));
   AOI21_X1 i_0_657_184 (.A(n_0_657_959), .B1(n_0_657_164), .B2(n_0_657_163), 
      .ZN(n_0_657_162));
   INV_X1 i_0_657_185 (.A(n_865), .ZN(n_0_657_163));
   NAND2_X1 i_0_657_186 (.A1(n_0_247), .A2(n_0_657_964), .ZN(n_0_657_164));
   OAI21_X1 i_0_657_187 (.A(n_0_657_169), .B1(n_0_657_165), .B2(n_0_657_167), 
      .ZN(n_0_828));
   OAI21_X1 i_0_657_188 (.A(n_0_657_959), .B1(n_0_657_166), .B2(n_988), .ZN(
      n_0_657_165));
   INV_X1 i_0_657_189 (.A(n_0_657_168), .ZN(n_0_657_166));
   NOR2_X1 i_0_657_190 (.A1(n_0_369), .A2(n_0_657_168), .ZN(n_0_657_167));
   NAND2_X1 i_0_657_191 (.A1(n_0_794), .A2(n_0_657_964), .ZN(n_0_657_168));
   OAI21_X1 i_0_657_192 (.A(n_0_657_170), .B1(n_0_579), .B2(n_0_657_172), 
      .ZN(n_0_657_169));
   AOI21_X1 i_0_657_193 (.A(n_0_657_959), .B1(n_0_657_172), .B2(n_0_657_171), 
      .ZN(n_0_657_170));
   INV_X1 i_0_657_194 (.A(n_988), .ZN(n_0_657_171));
   NAND2_X1 i_0_657_195 (.A1(n_0_246), .A2(n_0_657_964), .ZN(n_0_657_172));
   NAND2_X1 i_0_657_196 (.A1(n_0_657_173), .A2(n_0_657_176), .ZN(n_0_829));
   OAI21_X1 i_0_657_197 (.A(n_0_657_174), .B1(n_0_368), .B2(n_0_657_175), 
      .ZN(n_0_657_173));
   AOI21_X1 i_0_657_198 (.A(n_0_806), .B1(n_0_657_175), .B2(n_0_657_178), 
      .ZN(n_0_657_174));
   NAND2_X1 i_0_657_199 (.A1(n_0_793), .A2(n_0_657_964), .ZN(n_0_657_175));
   OAI21_X1 i_0_657_200 (.A(n_0_657_177), .B1(n_0_576), .B2(n_0_657_179), 
      .ZN(n_0_657_176));
   AOI21_X1 i_0_657_201 (.A(n_0_657_959), .B1(n_0_657_179), .B2(n_0_657_178), 
      .ZN(n_0_657_177));
   INV_X1 i_0_657_202 (.A(n_866), .ZN(n_0_657_178));
   NAND2_X1 i_0_657_203 (.A1(n_0_245), .A2(n_0_657_964), .ZN(n_0_657_179));
   NAND2_X1 i_0_657_204 (.A1(n_0_657_180), .A2(n_0_657_183), .ZN(n_0_830));
   OAI21_X1 i_0_657_205 (.A(n_0_657_181), .B1(n_0_367), .B2(n_0_657_182), 
      .ZN(n_0_657_180));
   AOI21_X1 i_0_657_206 (.A(n_0_806), .B1(n_0_657_182), .B2(n_0_657_185), 
      .ZN(n_0_657_181));
   NAND2_X1 i_0_657_207 (.A1(n_0_792), .A2(n_0_657_964), .ZN(n_0_657_182));
   OAI21_X1 i_0_657_208 (.A(n_0_657_184), .B1(n_0_573), .B2(n_0_657_186), 
      .ZN(n_0_657_183));
   AOI21_X1 i_0_657_209 (.A(n_0_657_959), .B1(n_0_657_185), .B2(n_0_657_186), 
      .ZN(n_0_657_184));
   INV_X1 i_0_657_210 (.A(n_867), .ZN(n_0_657_185));
   NAND2_X1 i_0_657_211 (.A1(n_0_244), .A2(n_0_657_964), .ZN(n_0_657_186));
   NAND2_X1 i_0_657_212 (.A1(n_0_657_187), .A2(n_0_657_190), .ZN(n_0_831));
   OAI21_X1 i_0_657_213 (.A(n_0_657_188), .B1(n_0_366), .B2(n_0_657_189), 
      .ZN(n_0_657_187));
   AOI21_X1 i_0_657_214 (.A(n_0_806), .B1(n_0_657_189), .B2(n_0_657_192), 
      .ZN(n_0_657_188));
   NAND2_X1 i_0_657_215 (.A1(n_0_791), .A2(n_0_657_964), .ZN(n_0_657_189));
   OAI21_X1 i_0_657_216 (.A(n_0_657_191), .B1(n_0_570), .B2(n_0_657_193), 
      .ZN(n_0_657_190));
   AOI21_X1 i_0_657_217 (.A(n_0_657_959), .B1(n_0_657_192), .B2(n_0_657_193), 
      .ZN(n_0_657_191));
   INV_X1 i_0_657_218 (.A(n_868), .ZN(n_0_657_192));
   NAND2_X1 i_0_657_219 (.A1(n_0_243), .A2(n_0_657_964), .ZN(n_0_657_193));
   NAND2_X1 i_0_657_220 (.A1(n_0_657_194), .A2(n_0_657_197), .ZN(n_0_832));
   OAI21_X1 i_0_657_221 (.A(n_0_657_195), .B1(n_0_365), .B2(n_0_657_196), 
      .ZN(n_0_657_194));
   AOI21_X1 i_0_657_222 (.A(n_0_806), .B1(n_0_657_196), .B2(n_0_657_199), 
      .ZN(n_0_657_195));
   NAND2_X1 i_0_657_223 (.A1(n_0_790), .A2(n_0_657_964), .ZN(n_0_657_196));
   OAI21_X1 i_0_657_224 (.A(n_0_657_198), .B1(n_0_611), .B2(n_0_657_200), 
      .ZN(n_0_657_197));
   AOI21_X1 i_0_657_225 (.A(n_0_657_959), .B1(n_0_657_200), .B2(n_0_657_199), 
      .ZN(n_0_657_198));
   INV_X1 i_0_657_226 (.A(n_869), .ZN(n_0_657_199));
   NAND2_X1 i_0_657_227 (.A1(n_0_242), .A2(n_0_657_964), .ZN(n_0_657_200));
   NAND2_X1 i_0_657_228 (.A1(n_0_657_201), .A2(n_0_657_204), .ZN(n_0_833));
   OAI21_X1 i_0_657_229 (.A(n_0_657_202), .B1(n_0_364), .B2(n_0_657_203), 
      .ZN(n_0_657_201));
   AOI21_X1 i_0_657_230 (.A(n_0_806), .B1(n_0_657_203), .B2(n_0_657_206), 
      .ZN(n_0_657_202));
   NAND2_X1 i_0_657_231 (.A1(n_0_789), .A2(n_0_657_964), .ZN(n_0_657_203));
   OAI21_X1 i_0_657_232 (.A(n_0_657_205), .B1(n_0_614), .B2(n_0_657_207), 
      .ZN(n_0_657_204));
   AOI21_X1 i_0_657_233 (.A(n_0_657_959), .B1(n_0_657_207), .B2(n_0_657_206), 
      .ZN(n_0_657_205));
   INV_X1 i_0_657_234 (.A(n_870), .ZN(n_0_657_206));
   NAND2_X1 i_0_657_235 (.A1(n_0_241), .A2(n_0_657_964), .ZN(n_0_657_207));
   NAND2_X1 i_0_657_236 (.A1(n_0_657_208), .A2(n_0_657_211), .ZN(n_0_834));
   OAI21_X1 i_0_657_237 (.A(n_0_657_209), .B1(n_0_363), .B2(n_0_657_210), 
      .ZN(n_0_657_208));
   AOI21_X1 i_0_657_238 (.A(n_0_806), .B1(n_0_657_210), .B2(n_0_657_213), 
      .ZN(n_0_657_209));
   NAND2_X1 i_0_657_239 (.A1(n_0_788), .A2(n_0_657_964), .ZN(n_0_657_210));
   OAI21_X1 i_0_657_240 (.A(n_0_657_212), .B1(n_0_617), .B2(n_0_657_214), 
      .ZN(n_0_657_211));
   AOI21_X1 i_0_657_241 (.A(n_0_657_959), .B1(n_0_657_213), .B2(n_0_657_214), 
      .ZN(n_0_657_212));
   INV_X1 i_0_657_242 (.A(n_984), .ZN(n_0_657_213));
   NAND2_X1 i_0_657_243 (.A1(n_0_240), .A2(n_0_657_964), .ZN(n_0_657_214));
   NAND2_X1 i_0_657_244 (.A1(n_0_657_215), .A2(n_0_657_218), .ZN(n_0_835));
   OAI21_X1 i_0_657_245 (.A(n_0_657_216), .B1(n_0_362), .B2(n_0_657_217), 
      .ZN(n_0_657_215));
   AOI21_X1 i_0_657_246 (.A(n_0_806), .B1(n_0_657_217), .B2(n_0_657_220), 
      .ZN(n_0_657_216));
   NAND2_X1 i_0_657_247 (.A1(n_0_787), .A2(n_0_657_964), .ZN(n_0_657_217));
   OAI21_X1 i_0_657_248 (.A(n_0_657_219), .B1(n_0_567), .B2(n_0_657_221), 
      .ZN(n_0_657_218));
   AOI21_X1 i_0_657_249 (.A(n_0_657_959), .B1(n_0_657_220), .B2(n_0_657_221), 
      .ZN(n_0_657_219));
   INV_X1 i_0_657_250 (.A(n_871), .ZN(n_0_657_220));
   NAND2_X1 i_0_657_251 (.A1(n_0_239), .A2(n_0_657_964), .ZN(n_0_657_221));
   NAND2_X1 i_0_657_252 (.A1(n_0_657_222), .A2(n_0_657_225), .ZN(n_0_836));
   OAI21_X1 i_0_657_253 (.A(n_0_657_223), .B1(n_0_361), .B2(n_0_657_224), 
      .ZN(n_0_657_222));
   AOI21_X1 i_0_657_254 (.A(n_0_806), .B1(n_0_657_224), .B2(n_0_657_227), 
      .ZN(n_0_657_223));
   NAND2_X1 i_0_657_255 (.A1(n_0_786), .A2(n_0_657_964), .ZN(n_0_657_224));
   OAI21_X1 i_0_657_256 (.A(n_0_657_226), .B1(n_0_620), .B2(n_0_657_228), 
      .ZN(n_0_657_225));
   AOI21_X1 i_0_657_257 (.A(n_0_657_959), .B1(n_0_657_228), .B2(n_0_657_227), 
      .ZN(n_0_657_226));
   INV_X1 i_0_657_258 (.A(n_872), .ZN(n_0_657_227));
   NAND2_X1 i_0_657_259 (.A1(n_0_238), .A2(n_0_657_964), .ZN(n_0_657_228));
   NAND2_X1 i_0_657_260 (.A1(n_0_657_232), .A2(n_0_657_229), .ZN(n_0_837));
   OAI21_X1 i_0_657_261 (.A(n_0_657_230), .B1(n_0_360), .B2(n_0_657_231), 
      .ZN(n_0_657_229));
   AOI21_X1 i_0_657_262 (.A(n_0_806), .B1(n_0_657_231), .B2(n_0_657_234), 
      .ZN(n_0_657_230));
   NAND2_X1 i_0_657_263 (.A1(n_0_785), .A2(n_0_657_964), .ZN(n_0_657_231));
   OAI21_X1 i_0_657_264 (.A(n_0_657_233), .B1(n_0_564), .B2(n_0_657_235), 
      .ZN(n_0_657_232));
   AOI21_X1 i_0_657_265 (.A(n_0_657_959), .B1(n_0_657_235), .B2(n_0_657_234), 
      .ZN(n_0_657_233));
   INV_X1 i_0_657_266 (.A(n_873), .ZN(n_0_657_234));
   NAND2_X1 i_0_657_267 (.A1(n_0_237), .A2(n_0_657_964), .ZN(n_0_657_235));
   NAND2_X1 i_0_657_268 (.A1(n_0_657_236), .A2(n_0_657_239), .ZN(n_0_838));
   OAI21_X1 i_0_657_269 (.A(n_0_657_237), .B1(n_0_359), .B2(n_0_657_238), 
      .ZN(n_0_657_236));
   AOI21_X1 i_0_657_270 (.A(n_0_806), .B1(n_0_657_238), .B2(n_0_657_241), 
      .ZN(n_0_657_237));
   NAND2_X1 i_0_657_271 (.A1(n_0_784), .A2(n_0_657_964), .ZN(n_0_657_238));
   OAI21_X1 i_0_657_272 (.A(n_0_657_240), .B1(n_0_561), .B2(n_0_657_242), 
      .ZN(n_0_657_239));
   AOI21_X1 i_0_657_273 (.A(n_0_657_959), .B1(n_0_657_242), .B2(n_0_657_241), 
      .ZN(n_0_657_240));
   INV_X1 i_0_657_274 (.A(n_874), .ZN(n_0_657_241));
   NAND2_X1 i_0_657_275 (.A1(n_0_236), .A2(n_0_657_964), .ZN(n_0_657_242));
   NAND2_X1 i_0_657_276 (.A1(n_0_657_243), .A2(n_0_657_246), .ZN(n_0_839));
   OAI21_X1 i_0_657_277 (.A(n_0_657_244), .B1(n_0_358), .B2(n_0_657_245), 
      .ZN(n_0_657_243));
   AOI21_X1 i_0_657_278 (.A(n_0_806), .B1(n_0_657_245), .B2(n_0_657_248), 
      .ZN(n_0_657_244));
   NAND2_X1 i_0_657_279 (.A1(n_0_783), .A2(n_0_657_964), .ZN(n_0_657_245));
   OAI21_X1 i_0_657_280 (.A(n_0_657_247), .B1(n_0_623), .B2(n_0_657_249), 
      .ZN(n_0_657_246));
   AOI21_X1 i_0_657_281 (.A(n_0_657_959), .B1(n_0_657_249), .B2(n_0_657_248), 
      .ZN(n_0_657_247));
   INV_X1 i_0_657_282 (.A(n_875), .ZN(n_0_657_248));
   NAND2_X1 i_0_657_283 (.A1(n_0_235), .A2(n_0_657_964), .ZN(n_0_657_249));
   NAND2_X1 i_0_657_284 (.A1(n_0_657_250), .A2(n_0_657_253), .ZN(n_0_840));
   OAI21_X1 i_0_657_285 (.A(n_0_657_251), .B1(n_0_357), .B2(n_0_657_252), 
      .ZN(n_0_657_250));
   AOI21_X1 i_0_657_286 (.A(n_0_806), .B1(n_0_657_252), .B2(n_0_657_255), 
      .ZN(n_0_657_251));
   NAND2_X1 i_0_657_287 (.A1(n_0_782), .A2(n_0_657_964), .ZN(n_0_657_252));
   OAI21_X1 i_0_657_288 (.A(n_0_657_254), .B1(n_0_558), .B2(n_0_657_256), 
      .ZN(n_0_657_253));
   AOI21_X1 i_0_657_289 (.A(n_0_657_959), .B1(n_0_657_256), .B2(n_0_657_255), 
      .ZN(n_0_657_254));
   INV_X1 i_0_657_290 (.A(n_876), .ZN(n_0_657_255));
   NAND2_X1 i_0_657_291 (.A1(n_0_234), .A2(n_0_657_964), .ZN(n_0_657_256));
   OAI21_X1 i_0_657_292 (.A(n_0_657_261), .B1(n_0_657_259), .B2(n_0_657_257), 
      .ZN(n_0_841));
   OAI21_X1 i_0_657_293 (.A(n_0_657_959), .B1(n_0_657_258), .B2(n_989), .ZN(
      n_0_657_257));
   INV_X1 i_0_657_294 (.A(n_0_657_260), .ZN(n_0_657_258));
   NOR2_X1 i_0_657_295 (.A1(n_0_356), .A2(n_0_657_260), .ZN(n_0_657_259));
   NAND2_X1 i_0_657_296 (.A1(n_0_781), .A2(n_0_657_964), .ZN(n_0_657_260));
   OAI21_X1 i_0_657_297 (.A(n_0_657_262), .B1(n_0_555), .B2(n_0_657_264), 
      .ZN(n_0_657_261));
   AOI21_X1 i_0_657_298 (.A(n_0_657_959), .B1(n_0_657_263), .B2(n_0_657_264), 
      .ZN(n_0_657_262));
   INV_X1 i_0_657_299 (.A(n_989), .ZN(n_0_657_263));
   NAND2_X1 i_0_657_300 (.A1(n_0_233), .A2(n_0_657_964), .ZN(n_0_657_264));
   OAI22_X1 i_0_657_301 (.A1(n_0_657_269), .A2(n_0_657_267), .B1(n_0_657_266), 
      .B2(n_0_657_265), .ZN(n_0_842));
   OAI21_X1 i_0_657_302 (.A(n_0_806), .B1(n_0_657_2), .B2(n_877), .ZN(
      n_0_657_265));
   NOR2_X1 i_0_657_303 (.A1(n_0_552), .A2(n_0_657_3), .ZN(n_0_657_266));
   OAI21_X1 i_0_657_304 (.A(n_0_657_959), .B1(n_0_657_268), .B2(n_877), .ZN(
      n_0_657_267));
   INV_X1 i_0_657_305 (.A(n_0_657_270), .ZN(n_0_657_268));
   NOR2_X1 i_0_657_306 (.A1(n_0_355), .A2(n_0_657_270), .ZN(n_0_657_269));
   NAND2_X1 i_0_657_307 (.A1(n_0_780), .A2(n_0_657_964), .ZN(n_0_657_270));
   NAND2_X1 i_0_657_308 (.A1(n_0_657_271), .A2(n_0_657_274), .ZN(n_0_843));
   OAI21_X1 i_0_657_309 (.A(n_0_657_272), .B1(n_0_354), .B2(n_0_657_273), 
      .ZN(n_0_657_271));
   AOI21_X1 i_0_657_310 (.A(n_0_806), .B1(n_0_657_273), .B2(n_0_657_276), 
      .ZN(n_0_657_272));
   NAND2_X1 i_0_657_311 (.A1(n_0_779), .A2(n_0_657_964), .ZN(n_0_657_273));
   OAI21_X1 i_0_657_312 (.A(n_0_657_275), .B1(n_0_626), .B2(n_0_657_277), 
      .ZN(n_0_657_274));
   AOI21_X1 i_0_657_313 (.A(n_0_657_959), .B1(n_0_657_277), .B2(n_0_657_276), 
      .ZN(n_0_657_275));
   INV_X1 i_0_657_314 (.A(n_878), .ZN(n_0_657_276));
   NAND2_X1 i_0_657_315 (.A1(n_0_231), .A2(n_0_657_964), .ZN(n_0_657_277));
   NAND2_X1 i_0_657_316 (.A1(n_0_657_278), .A2(n_0_657_281), .ZN(n_0_844));
   OAI21_X1 i_0_657_317 (.A(n_0_657_279), .B1(n_0_353), .B2(n_0_657_280), 
      .ZN(n_0_657_278));
   AOI21_X1 i_0_657_318 (.A(n_0_806), .B1(n_0_657_280), .B2(n_0_657_283), 
      .ZN(n_0_657_279));
   NAND2_X1 i_0_657_319 (.A1(n_0_778), .A2(n_0_657_964), .ZN(n_0_657_280));
   OAI21_X1 i_0_657_320 (.A(n_0_657_282), .B1(n_0_549), .B2(n_0_657_284), 
      .ZN(n_0_657_281));
   AOI21_X1 i_0_657_321 (.A(n_0_657_959), .B1(n_0_657_284), .B2(n_0_657_283), 
      .ZN(n_0_657_282));
   INV_X1 i_0_657_322 (.A(n_879), .ZN(n_0_657_283));
   NAND2_X1 i_0_657_323 (.A1(n_0_230), .A2(n_0_657_964), .ZN(n_0_657_284));
   OAI21_X1 i_0_657_324 (.A(n_0_657_285), .B1(n_0_657_291), .B2(n_0_657_289), 
      .ZN(n_0_845));
   OAI21_X1 i_0_657_325 (.A(n_0_657_286), .B1(n_0_352), .B2(n_0_657_288), 
      .ZN(n_0_657_285));
   AOI21_X1 i_0_657_326 (.A(n_0_806), .B1(n_0_657_288), .B2(n_0_657_287), 
      .ZN(n_0_657_286));
   INV_X1 i_0_657_327 (.A(n_880), .ZN(n_0_657_287));
   NAND2_X1 i_0_657_328 (.A1(n_0_777), .A2(n_0_657_964), .ZN(n_0_657_288));
   OAI21_X1 i_0_657_329 (.A(n_0_806), .B1(n_0_657_290), .B2(n_880), .ZN(
      n_0_657_289));
   INV_X1 i_0_657_330 (.A(n_0_657_292), .ZN(n_0_657_290));
   NOR2_X1 i_0_657_331 (.A1(n_0_629), .A2(n_0_657_292), .ZN(n_0_657_291));
   NAND2_X1 i_0_657_332 (.A1(n_0_229), .A2(n_0_657_964), .ZN(n_0_657_292));
   NAND2_X1 i_0_657_333 (.A1(n_0_657_293), .A2(n_0_657_296), .ZN(n_0_846));
   OAI21_X1 i_0_657_334 (.A(n_0_657_294), .B1(n_0_351), .B2(n_0_657_295), 
      .ZN(n_0_657_293));
   AOI21_X1 i_0_657_335 (.A(n_0_806), .B1(n_0_657_295), .B2(n_0_657_298), 
      .ZN(n_0_657_294));
   NAND2_X1 i_0_657_336 (.A1(n_0_776), .A2(n_0_657_964), .ZN(n_0_657_295));
   OAI21_X1 i_0_657_337 (.A(n_0_657_297), .B1(n_0_548), .B2(n_0_657_299), 
      .ZN(n_0_657_296));
   AOI21_X1 i_0_657_338 (.A(n_0_657_959), .B1(n_0_657_298), .B2(n_0_657_299), 
      .ZN(n_0_657_297));
   INV_X1 i_0_657_339 (.A(n_881), .ZN(n_0_657_298));
   NAND2_X1 i_0_657_340 (.A1(n_0_228), .A2(n_0_657_964), .ZN(n_0_657_299));
   OAI21_X1 i_0_657_341 (.A(n_0_657_304), .B1(n_0_657_302), .B2(n_0_657_300), 
      .ZN(n_0_847));
   OAI21_X1 i_0_657_342 (.A(n_0_657_959), .B1(n_0_657_301), .B2(n_990), .ZN(
      n_0_657_300));
   INV_X1 i_0_657_343 (.A(n_0_657_303), .ZN(n_0_657_301));
   NOR2_X1 i_0_657_344 (.A1(n_0_350), .A2(n_0_657_303), .ZN(n_0_657_302));
   NAND2_X1 i_0_657_345 (.A1(n_0_775), .A2(n_0_657_964), .ZN(n_0_657_303));
   OAI21_X1 i_0_657_346 (.A(n_0_657_305), .B1(n_0_632), .B2(n_0_657_307), 
      .ZN(n_0_657_304));
   AOI21_X1 i_0_657_347 (.A(n_0_657_959), .B1(n_0_657_307), .B2(n_0_657_306), 
      .ZN(n_0_657_305));
   INV_X1 i_0_657_348 (.A(n_990), .ZN(n_0_657_306));
   NAND2_X1 i_0_657_349 (.A1(n_0_227), .A2(n_0_657_964), .ZN(n_0_657_307));
   NAND2_X1 i_0_657_350 (.A1(n_0_657_308), .A2(n_0_657_311), .ZN(n_0_849));
   OAI21_X1 i_0_657_351 (.A(n_0_657_309), .B1(n_0_348), .B2(n_0_657_310), 
      .ZN(n_0_657_308));
   AOI21_X1 i_0_657_352 (.A(n_0_806), .B1(n_0_657_310), .B2(n_0_657_313), 
      .ZN(n_0_657_309));
   NAND2_X1 i_0_657_353 (.A1(n_0_773), .A2(n_0_657_964), .ZN(n_0_657_310));
   OAI21_X1 i_0_657_354 (.A(n_0_657_312), .B1(n_0_547), .B2(n_0_657_314), 
      .ZN(n_0_657_311));
   AOI21_X1 i_0_657_355 (.A(n_0_657_959), .B1(n_0_657_314), .B2(n_0_657_313), 
      .ZN(n_0_657_312));
   INV_X1 i_0_657_356 (.A(n_882), .ZN(n_0_657_313));
   NAND2_X1 i_0_657_357 (.A1(n_0_225), .A2(n_0_657_964), .ZN(n_0_657_314));
   NAND2_X1 i_0_657_358 (.A1(n_0_657_315), .A2(n_0_657_318), .ZN(n_0_850));
   OAI21_X1 i_0_657_359 (.A(n_0_657_316), .B1(n_0_347), .B2(n_0_657_317), 
      .ZN(n_0_657_315));
   AOI21_X1 i_0_657_360 (.A(n_0_806), .B1(n_0_657_317), .B2(n_0_657_320), 
      .ZN(n_0_657_316));
   NAND2_X1 i_0_657_361 (.A1(n_0_772), .A2(n_0_657_964), .ZN(n_0_657_317));
   OAI21_X1 i_0_657_362 (.A(n_0_657_319), .B1(n_0_638), .B2(n_0_657_321), 
      .ZN(n_0_657_318));
   AOI21_X1 i_0_657_363 (.A(n_0_657_959), .B1(n_0_657_321), .B2(n_0_657_320), 
      .ZN(n_0_657_319));
   INV_X1 i_0_657_364 (.A(n_883), .ZN(n_0_657_320));
   NAND2_X1 i_0_657_365 (.A1(n_0_224), .A2(n_0_657_964), .ZN(n_0_657_321));
   NAND2_X1 i_0_657_366 (.A1(n_0_657_322), .A2(n_0_657_325), .ZN(n_0_851));
   OAI21_X1 i_0_657_367 (.A(n_0_657_323), .B1(n_0_346), .B2(n_0_657_324), 
      .ZN(n_0_657_322));
   AOI21_X1 i_0_657_368 (.A(n_0_806), .B1(n_0_657_324), .B2(n_0_657_327), 
      .ZN(n_0_657_323));
   NAND2_X1 i_0_657_369 (.A1(n_0_771), .A2(n_0_657_964), .ZN(n_0_657_324));
   OAI21_X1 i_0_657_370 (.A(n_0_657_326), .B1(n_0_543), .B2(n_0_657_328), 
      .ZN(n_0_657_325));
   AOI21_X1 i_0_657_371 (.A(n_0_657_959), .B1(n_0_657_328), .B2(n_0_657_327), 
      .ZN(n_0_657_326));
   INV_X1 i_0_657_372 (.A(n_884), .ZN(n_0_657_327));
   NAND2_X1 i_0_657_373 (.A1(n_0_223), .A2(n_0_657_964), .ZN(n_0_657_328));
   NAND2_X1 i_0_657_374 (.A1(n_0_657_329), .A2(n_0_657_332), .ZN(n_0_852));
   OAI21_X1 i_0_657_375 (.A(n_0_657_330), .B1(n_0_345), .B2(n_0_657_331), 
      .ZN(n_0_657_329));
   AOI21_X1 i_0_657_376 (.A(n_0_806), .B1(n_0_657_331), .B2(n_0_657_334), 
      .ZN(n_0_657_330));
   NAND2_X1 i_0_657_377 (.A1(n_0_770), .A2(n_0_657_964), .ZN(n_0_657_331));
   OAI211_X1 i_0_657_378 (.A(n_0_657_333), .B(n_0_806), .C1(n_0_641), .C2(
      n_0_657_335), .ZN(n_0_657_332));
   NAND2_X1 i_0_657_379 (.A1(n_0_657_335), .A2(n_0_657_334), .ZN(n_0_657_333));
   INV_X1 i_0_657_380 (.A(n_982), .ZN(n_0_657_334));
   NAND2_X1 i_0_657_381 (.A1(n_0_222), .A2(n_0_657_964), .ZN(n_0_657_335));
   NAND2_X1 i_0_657_382 (.A1(n_0_657_336), .A2(n_0_657_339), .ZN(n_0_853));
   OAI21_X1 i_0_657_383 (.A(n_0_657_337), .B1(n_0_344), .B2(n_0_657_338), 
      .ZN(n_0_657_336));
   AOI21_X1 i_0_657_384 (.A(n_0_806), .B1(n_0_657_338), .B2(n_0_657_341), 
      .ZN(n_0_657_337));
   NAND2_X1 i_0_657_385 (.A1(n_0_769), .A2(n_0_657_964), .ZN(n_0_657_338));
   OAI21_X1 i_0_657_386 (.A(n_0_657_340), .B1(n_0_644), .B2(n_0_657_342), 
      .ZN(n_0_657_339));
   AOI21_X1 i_0_657_387 (.A(n_0_657_959), .B1(n_0_657_342), .B2(n_0_657_341), 
      .ZN(n_0_657_340));
   INV_X1 i_0_657_388 (.A(n_885), .ZN(n_0_657_341));
   NAND2_X1 i_0_657_389 (.A1(n_0_221), .A2(n_0_657_964), .ZN(n_0_657_342));
   OAI21_X1 i_0_657_390 (.A(n_0_657_347), .B1(n_0_657_345), .B2(n_0_657_343), 
      .ZN(n_0_854));
   OAI21_X1 i_0_657_391 (.A(n_0_657_959), .B1(n_0_657_344), .B2(n_886), .ZN(
      n_0_657_343));
   INV_X1 i_0_657_392 (.A(n_0_657_346), .ZN(n_0_657_344));
   NOR2_X1 i_0_657_393 (.A1(n_0_343), .A2(n_0_657_346), .ZN(n_0_657_345));
   NAND2_X1 i_0_657_394 (.A1(n_0_768), .A2(n_0_657_964), .ZN(n_0_657_346));
   OAI211_X1 i_0_657_395 (.A(n_0_657_348), .B(n_0_806), .C1(n_886), .C2(
      n_0_657_350), .ZN(n_0_657_347));
   NAND2_X1 i_0_657_396 (.A1(n_0_657_349), .A2(n_0_657_350), .ZN(n_0_657_348));
   INV_X1 i_0_657_397 (.A(n_0_540), .ZN(n_0_657_349));
   INV_X1 i_0_657_398 (.A(n_0_657_351), .ZN(n_0_657_350));
   NAND2_X1 i_0_657_399 (.A1(n_0_220), .A2(n_0_657_964), .ZN(n_0_657_351));
   OAI21_X1 i_0_657_400 (.A(n_0_657_356), .B1(n_0_657_354), .B2(n_0_657_352), 
      .ZN(n_0_855));
   OAI21_X1 i_0_657_401 (.A(n_0_657_959), .B1(n_0_657_353), .B2(n_991), .ZN(
      n_0_657_352));
   INV_X1 i_0_657_402 (.A(n_0_657_355), .ZN(n_0_657_353));
   NOR2_X1 i_0_657_403 (.A1(n_0_342), .A2(n_0_657_355), .ZN(n_0_657_354));
   NAND2_X1 i_0_657_404 (.A1(n_0_767), .A2(n_0_657_964), .ZN(n_0_657_355));
   OAI21_X1 i_0_657_405 (.A(n_0_657_357), .B1(n_0_537), .B2(n_0_657_359), 
      .ZN(n_0_657_356));
   AOI21_X1 i_0_657_406 (.A(n_0_657_959), .B1(n_0_657_358), .B2(n_0_657_359), 
      .ZN(n_0_657_357));
   INV_X1 i_0_657_407 (.A(n_991), .ZN(n_0_657_358));
   NAND2_X1 i_0_657_408 (.A1(n_0_219), .A2(n_0_657_964), .ZN(n_0_657_359));
   OAI21_X1 i_0_657_409 (.A(n_0_657_364), .B1(n_0_657_362), .B2(n_0_657_360), 
      .ZN(n_0_856));
   OAI21_X1 i_0_657_410 (.A(n_0_657_959), .B1(n_0_657_361), .B2(n_887), .ZN(
      n_0_657_360));
   INV_X1 i_0_657_411 (.A(n_0_657_363), .ZN(n_0_657_361));
   NOR2_X1 i_0_657_412 (.A1(n_0_341), .A2(n_0_657_363), .ZN(n_0_657_362));
   NAND2_X1 i_0_657_413 (.A1(n_0_766), .A2(n_0_657_964), .ZN(n_0_657_363));
   OAI211_X1 i_0_657_414 (.A(n_0_657_365), .B(n_0_806), .C1(n_887), .C2(
      n_0_657_367), .ZN(n_0_657_364));
   NAND2_X1 i_0_657_415 (.A1(n_0_657_366), .A2(n_0_657_367), .ZN(n_0_657_365));
   INV_X1 i_0_657_416 (.A(n_0_534), .ZN(n_0_657_366));
   INV_X1 i_0_657_417 (.A(n_0_657_368), .ZN(n_0_657_367));
   NAND2_X1 i_0_657_418 (.A1(n_0_218), .A2(n_0_657_964), .ZN(n_0_657_368));
   OAI21_X1 i_0_657_419 (.A(n_0_657_373), .B1(n_0_657_371), .B2(n_0_657_369), 
      .ZN(n_0_857));
   OAI21_X1 i_0_657_420 (.A(n_0_657_959), .B1(n_0_657_370), .B2(n_992), .ZN(
      n_0_657_369));
   INV_X1 i_0_657_421 (.A(n_0_657_372), .ZN(n_0_657_370));
   NOR2_X1 i_0_657_422 (.A1(n_0_340), .A2(n_0_657_372), .ZN(n_0_657_371));
   NAND2_X1 i_0_657_423 (.A1(n_0_765), .A2(n_0_657_964), .ZN(n_0_657_372));
   OAI21_X1 i_0_657_424 (.A(n_0_657_374), .B1(n_0_531), .B2(n_0_657_376), 
      .ZN(n_0_657_373));
   AOI21_X1 i_0_657_425 (.A(n_0_657_959), .B1(n_0_657_375), .B2(n_0_657_376), 
      .ZN(n_0_657_374));
   INV_X1 i_0_657_426 (.A(n_992), .ZN(n_0_657_375));
   NAND2_X1 i_0_657_427 (.A1(n_0_217), .A2(n_0_657_964), .ZN(n_0_657_376));
   NAND2_X1 i_0_657_428 (.A1(n_0_657_377), .A2(n_0_657_380), .ZN(n_0_858));
   OAI21_X1 i_0_657_429 (.A(n_0_657_378), .B1(n_0_339), .B2(n_0_657_379), 
      .ZN(n_0_657_377));
   AOI21_X1 i_0_657_430 (.A(n_0_806), .B1(n_0_657_379), .B2(n_0_657_382), 
      .ZN(n_0_657_378));
   NAND2_X1 i_0_657_431 (.A1(n_0_764), .A2(n_0_657_964), .ZN(n_0_657_379));
   OAI21_X1 i_0_657_432 (.A(n_0_657_381), .B1(n_0_528), .B2(n_0_657_383), 
      .ZN(n_0_657_380));
   AOI21_X1 i_0_657_433 (.A(n_0_657_959), .B1(n_0_657_383), .B2(n_0_657_382), 
      .ZN(n_0_657_381));
   INV_X1 i_0_657_434 (.A(n_888), .ZN(n_0_657_382));
   NAND2_X1 i_0_657_435 (.A1(n_0_216), .A2(n_0_657_964), .ZN(n_0_657_383));
   NAND2_X1 i_0_657_436 (.A1(n_0_657_384), .A2(n_0_657_387), .ZN(n_0_859));
   OAI21_X1 i_0_657_437 (.A(n_0_657_385), .B1(n_0_338), .B2(n_0_657_386), 
      .ZN(n_0_657_384));
   AOI21_X1 i_0_657_438 (.A(n_0_806), .B1(n_0_657_386), .B2(n_0_657_389), 
      .ZN(n_0_657_385));
   NAND2_X1 i_0_657_439 (.A1(n_0_763), .A2(n_0_657_964), .ZN(n_0_657_386));
   OAI211_X1 i_0_657_440 (.A(n_0_657_388), .B(n_0_806), .C1(n_0_525), .C2(
      n_0_657_390), .ZN(n_0_657_387));
   NAND2_X1 i_0_657_441 (.A1(n_0_657_390), .A2(n_0_657_389), .ZN(n_0_657_388));
   INV_X1 i_0_657_442 (.A(n_889), .ZN(n_0_657_389));
   NAND2_X1 i_0_657_443 (.A1(n_0_215), .A2(n_0_657_964), .ZN(n_0_657_390));
   NAND2_X1 i_0_657_444 (.A1(n_0_657_391), .A2(n_0_657_394), .ZN(n_0_860));
   OAI21_X1 i_0_657_445 (.A(n_0_657_392), .B1(n_0_337), .B2(n_0_657_393), 
      .ZN(n_0_657_391));
   AOI21_X1 i_0_657_446 (.A(n_0_806), .B1(n_0_657_393), .B2(n_0_657_396), 
      .ZN(n_0_657_392));
   NAND2_X1 i_0_657_447 (.A1(n_0_762), .A2(n_0_657_964), .ZN(n_0_657_393));
   OAI21_X1 i_0_657_448 (.A(n_0_657_395), .B1(n_0_522), .B2(n_0_657_397), 
      .ZN(n_0_657_394));
   AOI21_X1 i_0_657_449 (.A(n_0_657_959), .B1(n_0_657_397), .B2(n_0_657_396), 
      .ZN(n_0_657_395));
   INV_X1 i_0_657_450 (.A(n_890), .ZN(n_0_657_396));
   NAND2_X1 i_0_657_451 (.A1(n_0_214), .A2(n_0_657_964), .ZN(n_0_657_397));
   OAI21_X1 i_0_657_452 (.A(n_0_657_402), .B1(n_0_657_400), .B2(n_0_657_398), 
      .ZN(n_0_861));
   OAI21_X1 i_0_657_453 (.A(n_0_657_959), .B1(n_0_657_399), .B2(n_993), .ZN(
      n_0_657_398));
   INV_X1 i_0_657_454 (.A(n_0_657_401), .ZN(n_0_657_399));
   NOR2_X1 i_0_657_455 (.A1(n_0_336), .A2(n_0_657_401), .ZN(n_0_657_400));
   NAND2_X1 i_0_657_456 (.A1(n_0_761), .A2(n_0_657_964), .ZN(n_0_657_401));
   OAI21_X1 i_0_657_457 (.A(n_0_657_403), .B1(n_0_519), .B2(n_0_657_405), 
      .ZN(n_0_657_402));
   AOI21_X1 i_0_657_458 (.A(n_0_657_959), .B1(n_0_657_404), .B2(n_0_657_405), 
      .ZN(n_0_657_403));
   INV_X1 i_0_657_459 (.A(n_993), .ZN(n_0_657_404));
   NAND2_X1 i_0_657_460 (.A1(n_0_213), .A2(n_0_657_964), .ZN(n_0_657_405));
   NAND2_X1 i_0_657_461 (.A1(n_0_657_406), .A2(n_0_657_409), .ZN(n_0_862));
   OAI21_X1 i_0_657_462 (.A(n_0_657_407), .B1(n_0_335), .B2(n_0_657_408), 
      .ZN(n_0_657_406));
   AOI21_X1 i_0_657_463 (.A(n_0_806), .B1(n_0_657_408), .B2(n_0_657_411), 
      .ZN(n_0_657_407));
   NAND2_X1 i_0_657_464 (.A1(n_0_760), .A2(n_0_657_964), .ZN(n_0_657_408));
   OAI21_X1 i_0_657_465 (.A(n_0_657_410), .B1(n_0_516), .B2(n_0_657_412), 
      .ZN(n_0_657_409));
   AOI21_X1 i_0_657_466 (.A(n_0_657_959), .B1(n_0_657_412), .B2(n_0_657_411), 
      .ZN(n_0_657_410));
   INV_X1 i_0_657_467 (.A(n_891), .ZN(n_0_657_411));
   NAND2_X1 i_0_657_468 (.A1(n_0_212), .A2(n_0_657_964), .ZN(n_0_657_412));
   NAND2_X1 i_0_657_469 (.A1(n_0_657_413), .A2(n_0_657_418), .ZN(n_0_863));
   OAI211_X1 i_0_657_470 (.A(n_0_657_959), .B(n_0_657_414), .C1(n_0_657_416), 
      .C2(n_892), .ZN(n_0_657_413));
   NAND3_X1 i_0_657_471 (.A1(n_0_759), .A2(n_0_657_415), .A3(n_0_657_964), 
      .ZN(n_0_657_414));
   INV_X1 i_0_657_472 (.A(n_0_334), .ZN(n_0_657_415));
   INV_X1 i_0_657_473 (.A(n_0_657_417), .ZN(n_0_657_416));
   NAND2_X1 i_0_657_474 (.A1(n_0_759), .A2(n_0_657_964), .ZN(n_0_657_417));
   OAI211_X1 i_0_657_475 (.A(n_0_657_419), .B(n_0_806), .C1(n_892), .C2(
      n_0_657_421), .ZN(n_0_657_418));
   NAND2_X1 i_0_657_476 (.A1(n_0_657_420), .A2(n_0_657_421), .ZN(n_0_657_419));
   INV_X1 i_0_657_477 (.A(n_0_513), .ZN(n_0_657_420));
   INV_X1 i_0_657_478 (.A(n_0_657_422), .ZN(n_0_657_421));
   NAND2_X1 i_0_657_479 (.A1(n_0_211), .A2(n_0_657_964), .ZN(n_0_657_422));
   NAND2_X1 i_0_657_480 (.A1(n_0_657_423), .A2(n_0_657_426), .ZN(n_0_864));
   OAI21_X1 i_0_657_481 (.A(n_0_657_424), .B1(n_0_333), .B2(n_0_657_425), 
      .ZN(n_0_657_423));
   AOI21_X1 i_0_657_482 (.A(n_0_806), .B1(n_0_657_425), .B2(n_0_657_428), 
      .ZN(n_0_657_424));
   NAND2_X1 i_0_657_483 (.A1(n_0_758), .A2(n_0_657_964), .ZN(n_0_657_425));
   OAI21_X1 i_0_657_484 (.A(n_0_657_427), .B1(n_0_510), .B2(n_0_657_429), 
      .ZN(n_0_657_426));
   AOI21_X1 i_0_657_485 (.A(n_0_657_959), .B1(n_0_657_429), .B2(n_0_657_428), 
      .ZN(n_0_657_427));
   INV_X1 i_0_657_486 (.A(n_893), .ZN(n_0_657_428));
   NAND2_X1 i_0_657_487 (.A1(n_0_210), .A2(n_0_657_964), .ZN(n_0_657_429));
   NAND2_X1 i_0_657_488 (.A1(n_0_657_430), .A2(n_0_657_433), .ZN(n_0_865));
   OAI21_X1 i_0_657_489 (.A(n_0_657_431), .B1(n_0_332), .B2(n_0_657_432), 
      .ZN(n_0_657_430));
   AOI21_X1 i_0_657_490 (.A(n_0_806), .B1(n_0_657_432), .B2(n_0_657_435), 
      .ZN(n_0_657_431));
   NAND2_X1 i_0_657_491 (.A1(n_0_757), .A2(n_0_657_964), .ZN(n_0_657_432));
   OAI21_X1 i_0_657_492 (.A(n_0_657_434), .B1(n_0_507), .B2(n_0_657_436), 
      .ZN(n_0_657_433));
   AOI21_X1 i_0_657_493 (.A(n_0_657_959), .B1(n_0_657_436), .B2(n_0_657_435), 
      .ZN(n_0_657_434));
   INV_X1 i_0_657_494 (.A(n_894), .ZN(n_0_657_435));
   NAND2_X1 i_0_657_495 (.A1(n_0_209), .A2(n_0_657_964), .ZN(n_0_657_436));
   OAI22_X1 i_0_657_496 (.A1(n_0_657_441), .A2(n_0_657_439), .B1(n_0_657_438), 
      .B2(n_0_657_437), .ZN(n_0_866));
   OAI21_X1 i_0_657_497 (.A(n_0_806), .B1(n_0_657_10), .B2(n_895), .ZN(
      n_0_657_437));
   NOR2_X1 i_0_657_498 (.A1(n_0_504), .A2(n_0_657_11), .ZN(n_0_657_438));
   OAI21_X1 i_0_657_499 (.A(n_0_657_959), .B1(n_0_657_440), .B2(n_895), .ZN(
      n_0_657_439));
   INV_X1 i_0_657_500 (.A(n_0_657_442), .ZN(n_0_657_440));
   NOR2_X1 i_0_657_501 (.A1(n_0_331), .A2(n_0_657_442), .ZN(n_0_657_441));
   NAND2_X1 i_0_657_502 (.A1(n_0_756), .A2(n_0_657_964), .ZN(n_0_657_442));
   NAND2_X1 i_0_657_503 (.A1(n_0_657_443), .A2(n_0_657_446), .ZN(n_0_867));
   OAI21_X1 i_0_657_504 (.A(n_0_657_444), .B1(n_0_330), .B2(n_0_657_445), 
      .ZN(n_0_657_443));
   AOI21_X1 i_0_657_505 (.A(n_0_806), .B1(n_0_657_445), .B2(n_0_657_448), 
      .ZN(n_0_657_444));
   NAND2_X1 i_0_657_506 (.A1(n_0_755), .A2(n_0_657_964), .ZN(n_0_657_445));
   OAI21_X1 i_0_657_507 (.A(n_0_657_447), .B1(n_0_647), .B2(n_0_657_449), 
      .ZN(n_0_657_446));
   AOI21_X1 i_0_657_508 (.A(n_0_657_959), .B1(n_0_657_449), .B2(n_0_657_448), 
      .ZN(n_0_657_447));
   INV_X1 i_0_657_509 (.A(n_896), .ZN(n_0_657_448));
   NAND2_X1 i_0_657_510 (.A1(n_0_207), .A2(n_0_657_964), .ZN(n_0_657_449));
   OAI21_X1 i_0_657_511 (.A(n_0_657_454), .B1(n_0_657_452), .B2(n_0_657_450), 
      .ZN(n_0_868));
   OAI21_X1 i_0_657_512 (.A(n_0_657_959), .B1(n_0_657_451), .B2(n_994), .ZN(
      n_0_657_450));
   INV_X1 i_0_657_513 (.A(n_0_657_453), .ZN(n_0_657_451));
   NOR2_X1 i_0_657_514 (.A1(n_0_329), .A2(n_0_657_453), .ZN(n_0_657_452));
   NAND2_X1 i_0_657_515 (.A1(n_0_754), .A2(n_0_657_964), .ZN(n_0_657_453));
   OAI21_X1 i_0_657_516 (.A(n_0_657_455), .B1(n_0_501), .B2(n_0_657_457), 
      .ZN(n_0_657_454));
   AOI21_X1 i_0_657_517 (.A(n_0_657_959), .B1(n_0_657_456), .B2(n_0_657_457), 
      .ZN(n_0_657_455));
   INV_X1 i_0_657_518 (.A(n_994), .ZN(n_0_657_456));
   NAND2_X1 i_0_657_519 (.A1(n_0_206), .A2(n_0_657_964), .ZN(n_0_657_457));
   OAI21_X1 i_0_657_520 (.A(n_0_657_462), .B1(n_0_657_460), .B2(n_0_657_458), 
      .ZN(n_0_869));
   OAI21_X1 i_0_657_521 (.A(n_0_657_959), .B1(n_0_657_459), .B2(n_995), .ZN(
      n_0_657_458));
   INV_X1 i_0_657_522 (.A(n_0_657_461), .ZN(n_0_657_459));
   NOR2_X1 i_0_657_523 (.A1(n_0_328), .A2(n_0_657_461), .ZN(n_0_657_460));
   NAND2_X1 i_0_657_524 (.A1(n_0_753), .A2(n_0_657_964), .ZN(n_0_657_461));
   OAI21_X1 i_0_657_525 (.A(n_0_657_463), .B1(n_0_498), .B2(n_0_657_465), 
      .ZN(n_0_657_462));
   AOI21_X1 i_0_657_526 (.A(n_0_657_959), .B1(n_0_657_464), .B2(n_0_657_465), 
      .ZN(n_0_657_463));
   INV_X1 i_0_657_527 (.A(n_995), .ZN(n_0_657_464));
   NAND2_X1 i_0_657_528 (.A1(n_0_205), .A2(n_0_657_964), .ZN(n_0_657_465));
   OAI21_X1 i_0_657_529 (.A(n_0_657_470), .B1(n_0_657_468), .B2(n_0_657_466), 
      .ZN(n_0_870));
   OAI21_X1 i_0_657_530 (.A(n_0_657_959), .B1(n_0_657_467), .B2(n_996), .ZN(
      n_0_657_466));
   INV_X1 i_0_657_531 (.A(n_0_657_469), .ZN(n_0_657_467));
   NOR2_X1 i_0_657_532 (.A1(n_0_327), .A2(n_0_657_469), .ZN(n_0_657_468));
   NAND2_X1 i_0_657_533 (.A1(n_0_752), .A2(n_0_657_964), .ZN(n_0_657_469));
   OAI21_X1 i_0_657_534 (.A(n_0_657_471), .B1(n_0_495), .B2(n_0_657_473), 
      .ZN(n_0_657_470));
   AOI21_X1 i_0_657_535 (.A(n_0_657_959), .B1(n_0_657_472), .B2(n_0_657_473), 
      .ZN(n_0_657_471));
   INV_X1 i_0_657_536 (.A(n_996), .ZN(n_0_657_472));
   NAND2_X1 i_0_657_537 (.A1(n_0_204), .A2(n_0_657_964), .ZN(n_0_657_473));
   OAI21_X1 i_0_657_538 (.A(n_0_657_478), .B1(n_0_657_476), .B2(n_0_657_474), 
      .ZN(n_0_871));
   OAI21_X1 i_0_657_539 (.A(n_0_657_959), .B1(n_0_657_475), .B2(n_997), .ZN(
      n_0_657_474));
   INV_X1 i_0_657_540 (.A(n_0_657_477), .ZN(n_0_657_475));
   NOR2_X1 i_0_657_541 (.A1(n_0_326), .A2(n_0_657_477), .ZN(n_0_657_476));
   NAND2_X1 i_0_657_542 (.A1(n_0_751), .A2(n_0_657_964), .ZN(n_0_657_477));
   OAI21_X1 i_0_657_543 (.A(n_0_657_479), .B1(n_0_492), .B2(n_0_657_481), 
      .ZN(n_0_657_478));
   AOI21_X1 i_0_657_544 (.A(n_0_657_959), .B1(n_0_657_481), .B2(n_0_657_480), 
      .ZN(n_0_657_479));
   INV_X1 i_0_657_545 (.A(n_997), .ZN(n_0_657_480));
   NAND2_X1 i_0_657_546 (.A1(n_0_203), .A2(n_0_657_964), .ZN(n_0_657_481));
   OAI22_X1 i_0_657_547 (.A1(n_0_657_486), .A2(n_0_657_484), .B1(n_0_657_483), 
      .B2(n_0_657_482), .ZN(n_0_872));
   OAI21_X1 i_0_657_548 (.A(n_0_806), .B1(n_0_657_12), .B2(n_897), .ZN(
      n_0_657_482));
   NOR2_X1 i_0_657_549 (.A1(n_0_489), .A2(n_0_657_13), .ZN(n_0_657_483));
   OAI21_X1 i_0_657_550 (.A(n_0_657_959), .B1(n_0_657_485), .B2(n_897), .ZN(
      n_0_657_484));
   INV_X1 i_0_657_551 (.A(n_0_657_487), .ZN(n_0_657_485));
   NOR2_X1 i_0_657_552 (.A1(n_0_325), .A2(n_0_657_487), .ZN(n_0_657_486));
   NAND2_X1 i_0_657_553 (.A1(n_0_750), .A2(n_0_657_964), .ZN(n_0_657_487));
   OAI22_X1 i_0_657_554 (.A1(n_0_657_492), .A2(n_0_657_490), .B1(n_0_657_489), 
      .B2(n_0_657_488), .ZN(n_0_873));
   OAI21_X1 i_0_657_555 (.A(n_0_806), .B1(n_0_657_14), .B2(n_898), .ZN(
      n_0_657_488));
   NOR2_X1 i_0_657_556 (.A1(n_0_486), .A2(n_0_657_15), .ZN(n_0_657_489));
   OAI21_X1 i_0_657_557 (.A(n_0_657_959), .B1(n_0_657_491), .B2(n_898), .ZN(
      n_0_657_490));
   INV_X1 i_0_657_558 (.A(n_0_657_493), .ZN(n_0_657_491));
   NOR2_X1 i_0_657_559 (.A1(n_0_324), .A2(n_0_657_493), .ZN(n_0_657_492));
   NAND2_X1 i_0_657_560 (.A1(n_0_749), .A2(n_0_657_964), .ZN(n_0_657_493));
   OAI22_X1 i_0_657_561 (.A1(n_0_657_498), .A2(n_0_657_496), .B1(n_0_657_495), 
      .B2(n_0_657_494), .ZN(n_0_874));
   OAI21_X1 i_0_657_562 (.A(n_0_806), .B1(n_0_657_16), .B2(n_899), .ZN(
      n_0_657_494));
   NOR2_X1 i_0_657_563 (.A1(n_0_483), .A2(n_0_657_17), .ZN(n_0_657_495));
   OAI21_X1 i_0_657_564 (.A(n_0_657_959), .B1(n_0_657_497), .B2(n_899), .ZN(
      n_0_657_496));
   INV_X1 i_0_657_565 (.A(n_0_657_499), .ZN(n_0_657_497));
   NOR2_X1 i_0_657_566 (.A1(n_0_323), .A2(n_0_657_499), .ZN(n_0_657_498));
   NAND2_X1 i_0_657_567 (.A1(n_0_748), .A2(n_0_657_964), .ZN(n_0_657_499));
   OAI21_X1 i_0_657_568 (.A(n_0_657_504), .B1(n_0_657_502), .B2(n_0_657_500), 
      .ZN(n_0_875));
   OAI21_X1 i_0_657_569 (.A(n_0_657_959), .B1(n_0_657_501), .B2(n_900), .ZN(
      n_0_657_500));
   INV_X1 i_0_657_570 (.A(n_0_657_503), .ZN(n_0_657_501));
   NOR2_X1 i_0_657_571 (.A1(n_0_322), .A2(n_0_657_503), .ZN(n_0_657_502));
   NAND2_X1 i_0_657_572 (.A1(n_0_747), .A2(n_0_657_964), .ZN(n_0_657_503));
   OAI211_X1 i_0_657_573 (.A(n_0_657_505), .B(n_0_806), .C1(n_900), .C2(
      n_0_657_507), .ZN(n_0_657_504));
   NAND2_X1 i_0_657_574 (.A1(n_0_657_506), .A2(n_0_657_507), .ZN(n_0_657_505));
   INV_X1 i_0_657_575 (.A(n_0_650), .ZN(n_0_657_506));
   INV_X1 i_0_657_576 (.A(n_0_657_508), .ZN(n_0_657_507));
   NAND2_X1 i_0_657_577 (.A1(n_0_199), .A2(n_0_657_964), .ZN(n_0_657_508));
   OAI22_X1 i_0_657_578 (.A1(n_0_657_513), .A2(n_0_657_511), .B1(n_0_657_510), 
      .B2(n_0_657_509), .ZN(n_0_876));
   OAI21_X1 i_0_657_579 (.A(n_0_806), .B1(n_0_657_18), .B2(n_901), .ZN(
      n_0_657_509));
   NOR2_X1 i_0_657_580 (.A1(n_0_480), .A2(n_0_657_19), .ZN(n_0_657_510));
   OAI21_X1 i_0_657_581 (.A(n_0_657_959), .B1(n_0_657_512), .B2(n_901), .ZN(
      n_0_657_511));
   INV_X1 i_0_657_582 (.A(n_0_657_514), .ZN(n_0_657_512));
   NOR2_X1 i_0_657_583 (.A1(n_0_321), .A2(n_0_657_514), .ZN(n_0_657_513));
   NAND2_X1 i_0_657_584 (.A1(n_0_746), .A2(n_0_657_964), .ZN(n_0_657_514));
   NAND2_X1 i_0_657_585 (.A1(n_0_657_515), .A2(n_0_657_518), .ZN(n_0_877));
   OAI21_X1 i_0_657_586 (.A(n_0_657_516), .B1(n_0_320), .B2(n_0_657_517), 
      .ZN(n_0_657_515));
   AOI21_X1 i_0_657_587 (.A(n_0_806), .B1(n_0_657_517), .B2(n_0_657_520), 
      .ZN(n_0_657_516));
   NAND2_X1 i_0_657_588 (.A1(n_0_745), .A2(n_0_657_964), .ZN(n_0_657_517));
   OAI211_X1 i_0_657_589 (.A(n_0_657_519), .B(n_0_806), .C1(n_0_477), .C2(
      n_0_657_521), .ZN(n_0_657_518));
   NAND2_X1 i_0_657_590 (.A1(n_0_657_521), .A2(n_0_657_520), .ZN(n_0_657_519));
   INV_X1 i_0_657_591 (.A(n_902), .ZN(n_0_657_520));
   NAND2_X1 i_0_657_592 (.A1(n_0_197), .A2(n_0_657_964), .ZN(n_0_657_521));
   OAI22_X1 i_0_657_593 (.A1(n_0_657_526), .A2(n_0_657_524), .B1(n_0_657_523), 
      .B2(n_0_657_522), .ZN(n_0_878));
   OAI21_X1 i_0_657_594 (.A(n_0_806), .B1(n_0_657_20), .B2(n_903), .ZN(
      n_0_657_522));
   NOR2_X1 i_0_657_595 (.A1(n_0_474), .A2(n_0_657_21), .ZN(n_0_657_523));
   OAI21_X1 i_0_657_596 (.A(n_0_657_959), .B1(n_0_657_525), .B2(n_903), .ZN(
      n_0_657_524));
   INV_X1 i_0_657_597 (.A(n_0_657_527), .ZN(n_0_657_525));
   NOR2_X1 i_0_657_598 (.A1(n_0_319), .A2(n_0_657_527), .ZN(n_0_657_526));
   NAND2_X1 i_0_657_599 (.A1(n_0_744), .A2(n_0_657_964), .ZN(n_0_657_527));
   NAND2_X1 i_0_657_600 (.A1(n_0_657_528), .A2(n_0_657_531), .ZN(n_0_880));
   OAI21_X1 i_0_657_601 (.A(n_0_657_529), .B1(n_0_317), .B2(n_0_657_530), 
      .ZN(n_0_657_528));
   AOI21_X1 i_0_657_602 (.A(n_0_806), .B1(n_0_657_530), .B2(n_0_657_533), 
      .ZN(n_0_657_529));
   NAND2_X1 i_0_657_603 (.A1(n_0_742), .A2(n_0_657_964), .ZN(n_0_657_530));
   OAI21_X1 i_0_657_604 (.A(n_0_657_532), .B1(n_0_653), .B2(n_0_657_534), 
      .ZN(n_0_657_531));
   AOI21_X1 i_0_657_605 (.A(n_0_657_959), .B1(n_0_657_534), .B2(n_0_657_533), 
      .ZN(n_0_657_532));
   INV_X1 i_0_657_606 (.A(n_904), .ZN(n_0_657_533));
   NAND2_X1 i_0_657_607 (.A1(n_0_194), .A2(n_0_657_964), .ZN(n_0_657_534));
   NAND2_X1 i_0_657_608 (.A1(n_0_657_535), .A2(n_0_657_538), .ZN(n_0_881));
   OAI21_X1 i_0_657_609 (.A(n_0_657_536), .B1(n_0_316), .B2(n_0_657_537), 
      .ZN(n_0_657_535));
   AOI21_X1 i_0_657_610 (.A(n_0_806), .B1(n_0_657_537), .B2(n_0_657_540), 
      .ZN(n_0_657_536));
   NAND2_X1 i_0_657_611 (.A1(n_1290), .A2(n_0_657_964), .ZN(n_0_657_537));
   OAI211_X1 i_0_657_612 (.A(n_0_657_539), .B(n_0_806), .C1(n_0_808), .C2(
      n_0_657_541), .ZN(n_0_657_538));
   NAND2_X1 i_0_657_613 (.A1(n_0_657_541), .A2(n_0_657_540), .ZN(n_0_657_539));
   INV_X1 i_0_657_614 (.A(n_905), .ZN(n_0_657_540));
   NAND2_X1 i_0_657_615 (.A1(n_0_193), .A2(n_0_657_964), .ZN(n_0_657_541));
   NAND2_X1 i_0_657_616 (.A1(n_0_657_542), .A2(n_0_657_545), .ZN(n_0_882));
   OAI21_X1 i_0_657_617 (.A(n_0_657_543), .B1(n_0_315), .B2(n_0_657_544), 
      .ZN(n_0_657_542));
   AOI21_X1 i_0_657_618 (.A(n_0_806), .B1(n_0_657_544), .B2(n_0_657_547), 
      .ZN(n_0_657_543));
   NAND2_X1 i_0_657_619 (.A1(n_0_741), .A2(n_0_657_964), .ZN(n_0_657_544));
   OAI21_X1 i_0_657_620 (.A(n_0_657_546), .B1(n_0_471), .B2(n_0_657_548), 
      .ZN(n_0_657_545));
   AOI21_X1 i_0_657_621 (.A(n_0_657_959), .B1(n_0_657_548), .B2(n_0_657_547), 
      .ZN(n_0_657_546));
   INV_X1 i_0_657_622 (.A(n_906), .ZN(n_0_657_547));
   NAND2_X1 i_0_657_623 (.A1(n_0_192), .A2(n_0_657_964), .ZN(n_0_657_548));
   NAND2_X1 i_0_657_624 (.A1(n_0_657_554), .A2(n_0_657_549), .ZN(n_0_883));
   NAND3_X1 i_0_657_625 (.A1(n_0_657_552), .A2(n_0_657_550), .A3(n_0_657_959), 
      .ZN(n_0_657_549));
   OAI21_X1 i_0_657_626 (.A(n_0_657_559), .B1(n_0_657_551), .B2(n_0_657_813), 
      .ZN(n_0_657_550));
   INV_X1 i_0_657_627 (.A(n_0_740), .ZN(n_0_657_551));
   NAND3_X1 i_0_657_628 (.A1(n_0_657_553), .A2(n_0_740), .A3(n_0_657_964), 
      .ZN(n_0_657_552));
   INV_X1 i_0_657_629 (.A(n_0_314), .ZN(n_0_657_553));
   NAND3_X1 i_0_657_630 (.A1(n_0_657_557), .A2(n_0_806), .A3(n_0_657_555), 
      .ZN(n_0_657_554));
   NAND3_X1 i_0_657_631 (.A1(n_0_191), .A2(n_0_657_556), .A3(n_0_657_964), 
      .ZN(n_0_657_555));
   INV_X1 i_0_657_632 (.A(n_0_468), .ZN(n_0_657_556));
   NAND2_X1 i_0_657_633 (.A1(n_0_657_558), .A2(n_0_657_559), .ZN(n_0_657_557));
   NAND2_X1 i_0_657_634 (.A1(n_0_191), .A2(n_0_657_964), .ZN(n_0_657_558));
   INV_X1 i_0_657_635 (.A(n_907), .ZN(n_0_657_559));
   NAND2_X1 i_0_657_636 (.A1(n_0_657_560), .A2(n_0_657_563), .ZN(n_0_884));
   OAI21_X1 i_0_657_637 (.A(n_0_657_561), .B1(n_0_313), .B2(n_0_657_562), 
      .ZN(n_0_657_560));
   AOI21_X1 i_0_657_638 (.A(n_0_806), .B1(n_0_657_562), .B2(n_0_657_565), 
      .ZN(n_0_657_561));
   NAND2_X1 i_0_657_639 (.A1(n_0_739), .A2(n_0_657_964), .ZN(n_0_657_562));
   OAI21_X1 i_0_657_640 (.A(n_0_657_564), .B1(n_0_465), .B2(n_0_657_566), 
      .ZN(n_0_657_563));
   AOI21_X1 i_0_657_641 (.A(n_0_657_959), .B1(n_0_657_566), .B2(n_0_657_565), 
      .ZN(n_0_657_564));
   INV_X1 i_0_657_642 (.A(n_908), .ZN(n_0_657_565));
   NAND2_X1 i_0_657_643 (.A1(n_0_190), .A2(n_0_657_964), .ZN(n_0_657_566));
   OAI21_X1 i_0_657_644 (.A(n_0_657_571), .B1(n_0_657_569), .B2(n_0_657_567), 
      .ZN(n_0_885));
   OAI21_X1 i_0_657_645 (.A(n_0_657_959), .B1(n_0_657_568), .B2(n_998), .ZN(
      n_0_657_567));
   INV_X1 i_0_657_646 (.A(n_0_657_570), .ZN(n_0_657_568));
   NOR2_X1 i_0_657_647 (.A1(n_0_312), .A2(n_0_657_570), .ZN(n_0_657_569));
   NAND2_X1 i_0_657_648 (.A1(n_0_738), .A2(n_0_657_964), .ZN(n_0_657_570));
   OAI21_X1 i_0_657_649 (.A(n_0_657_572), .B1(n_0_462), .B2(n_0_657_574), 
      .ZN(n_0_657_571));
   AOI21_X1 i_0_657_650 (.A(n_0_657_959), .B1(n_0_657_574), .B2(n_0_657_573), 
      .ZN(n_0_657_572));
   INV_X1 i_0_657_651 (.A(n_998), .ZN(n_0_657_573));
   NAND2_X1 i_0_657_652 (.A1(n_0_189), .A2(n_0_657_964), .ZN(n_0_657_574));
   NAND2_X1 i_0_657_653 (.A1(n_0_657_575), .A2(n_0_657_578), .ZN(n_0_886));
   OAI21_X1 i_0_657_654 (.A(n_0_657_576), .B1(n_0_311), .B2(n_0_657_577), 
      .ZN(n_0_657_575));
   AOI21_X1 i_0_657_655 (.A(n_0_806), .B1(n_0_657_577), .B2(n_0_657_580), 
      .ZN(n_0_657_576));
   NAND2_X1 i_0_657_656 (.A1(n_0_737), .A2(n_0_657_964), .ZN(n_0_657_577));
   OAI21_X1 i_0_657_657 (.A(n_0_657_579), .B1(n_0_459), .B2(n_0_657_581), 
      .ZN(n_0_657_578));
   AOI21_X1 i_0_657_658 (.A(n_0_657_959), .B1(n_0_657_581), .B2(n_0_657_580), 
      .ZN(n_0_657_579));
   INV_X1 i_0_657_659 (.A(n_909), .ZN(n_0_657_580));
   NAND2_X1 i_0_657_660 (.A1(n_0_188), .A2(n_0_657_964), .ZN(n_0_657_581));
   OAI21_X1 i_0_657_661 (.A(n_0_657_586), .B1(n_0_657_584), .B2(n_0_657_582), 
      .ZN(n_0_887));
   OAI21_X1 i_0_657_662 (.A(n_0_657_959), .B1(n_0_657_583), .B2(n_1009), 
      .ZN(n_0_657_582));
   INV_X1 i_0_657_663 (.A(n_0_657_585), .ZN(n_0_657_583));
   NOR2_X1 i_0_657_664 (.A1(n_0_310), .A2(n_0_657_585), .ZN(n_0_657_584));
   NAND2_X1 i_0_657_665 (.A1(n_0_736), .A2(n_0_657_964), .ZN(n_0_657_585));
   OAI21_X1 i_0_657_666 (.A(n_0_657_587), .B1(n_0_456), .B2(n_0_657_589), 
      .ZN(n_0_657_586));
   AOI21_X1 i_0_657_667 (.A(n_0_657_959), .B1(n_0_657_588), .B2(n_0_657_589), 
      .ZN(n_0_657_587));
   INV_X1 i_0_657_668 (.A(n_1009), .ZN(n_0_657_588));
   NAND2_X1 i_0_657_669 (.A1(n_0_187), .A2(n_0_657_964), .ZN(n_0_657_589));
   OAI21_X1 i_0_657_670 (.A(n_0_657_594), .B1(n_0_657_592), .B2(n_0_657_590), 
      .ZN(n_0_888));
   OAI21_X1 i_0_657_671 (.A(n_0_657_959), .B1(n_0_657_591), .B2(n_999), .ZN(
      n_0_657_590));
   INV_X1 i_0_657_672 (.A(n_0_657_593), .ZN(n_0_657_591));
   NOR2_X1 i_0_657_673 (.A1(n_0_309), .A2(n_0_657_593), .ZN(n_0_657_592));
   NAND2_X1 i_0_657_674 (.A1(n_0_735), .A2(n_0_657_964), .ZN(n_0_657_593));
   OAI21_X1 i_0_657_675 (.A(n_0_657_595), .B1(n_0_455), .B2(n_0_657_597), 
      .ZN(n_0_657_594));
   AOI21_X1 i_0_657_676 (.A(n_0_657_959), .B1(n_0_657_596), .B2(n_0_657_597), 
      .ZN(n_0_657_595));
   INV_X1 i_0_657_677 (.A(n_999), .ZN(n_0_657_596));
   NAND2_X1 i_0_657_678 (.A1(n_0_186), .A2(n_0_657_964), .ZN(n_0_657_597));
   NAND2_X1 i_0_657_679 (.A1(n_0_657_598), .A2(n_0_657_601), .ZN(n_0_889));
   OAI21_X1 i_0_657_680 (.A(n_0_657_599), .B1(n_0_308), .B2(n_0_657_600), 
      .ZN(n_0_657_598));
   AOI21_X1 i_0_657_681 (.A(n_0_806), .B1(n_0_657_600), .B2(n_0_657_603), 
      .ZN(n_0_657_599));
   NAND2_X1 i_0_657_682 (.A1(n_0_734), .A2(n_0_657_964), .ZN(n_0_657_600));
   OAI21_X1 i_0_657_683 (.A(n_0_657_602), .B1(n_0_454), .B2(n_0_657_604), 
      .ZN(n_0_657_601));
   AOI21_X1 i_0_657_684 (.A(n_0_657_959), .B1(n_0_657_604), .B2(n_0_657_603), 
      .ZN(n_0_657_602));
   INV_X1 i_0_657_685 (.A(n_910), .ZN(n_0_657_603));
   NAND2_X1 i_0_657_686 (.A1(n_0_185), .A2(n_0_657_964), .ZN(n_0_657_604));
   OAI21_X1 i_0_657_687 (.A(n_0_657_609), .B1(n_0_657_607), .B2(n_0_657_605), 
      .ZN(n_0_890));
   OAI21_X1 i_0_657_688 (.A(n_0_657_959), .B1(n_0_657_606), .B2(n_1000), 
      .ZN(n_0_657_605));
   INV_X1 i_0_657_689 (.A(n_0_657_608), .ZN(n_0_657_606));
   NOR2_X1 i_0_657_690 (.A1(n_0_307), .A2(n_0_657_608), .ZN(n_0_657_607));
   NAND2_X1 i_0_657_691 (.A1(n_0_733), .A2(n_0_657_964), .ZN(n_0_657_608));
   OAI21_X1 i_0_657_692 (.A(n_0_657_610), .B1(n_0_451), .B2(n_0_657_612), 
      .ZN(n_0_657_609));
   AOI21_X1 i_0_657_693 (.A(n_0_657_959), .B1(n_0_657_611), .B2(n_0_657_612), 
      .ZN(n_0_657_610));
   INV_X1 i_0_657_694 (.A(n_1000), .ZN(n_0_657_611));
   NAND2_X1 i_0_657_695 (.A1(n_0_184), .A2(n_0_657_964), .ZN(n_0_657_612));
   OAI21_X1 i_0_657_696 (.A(n_0_657_617), .B1(n_0_657_615), .B2(n_0_657_613), 
      .ZN(n_0_891));
   OAI21_X1 i_0_657_697 (.A(n_0_657_959), .B1(n_0_657_614), .B2(n_1001), 
      .ZN(n_0_657_613));
   INV_X1 i_0_657_698 (.A(n_0_657_616), .ZN(n_0_657_614));
   NOR2_X1 i_0_657_699 (.A1(n_0_306), .A2(n_0_657_616), .ZN(n_0_657_615));
   NAND2_X1 i_0_657_700 (.A1(n_0_732), .A2(n_0_657_964), .ZN(n_0_657_616));
   OAI21_X1 i_0_657_701 (.A(n_0_657_618), .B1(n_0_448), .B2(n_0_657_620), 
      .ZN(n_0_657_617));
   AOI21_X1 i_0_657_702 (.A(n_0_657_959), .B1(n_0_657_619), .B2(n_0_657_620), 
      .ZN(n_0_657_618));
   INV_X1 i_0_657_703 (.A(n_1001), .ZN(n_0_657_619));
   NAND2_X1 i_0_657_704 (.A1(n_0_183), .A2(n_0_657_964), .ZN(n_0_657_620));
   NAND2_X1 i_0_657_705 (.A1(n_0_657_621), .A2(n_0_657_624), .ZN(n_0_892));
   OAI21_X1 i_0_657_706 (.A(n_0_657_622), .B1(n_0_305), .B2(n_0_657_623), 
      .ZN(n_0_657_621));
   AOI21_X1 i_0_657_707 (.A(n_0_806), .B1(n_0_657_623), .B2(n_0_657_626), 
      .ZN(n_0_657_622));
   NAND2_X1 i_0_657_708 (.A1(n_0_731), .A2(n_0_657_964), .ZN(n_0_657_623));
   OAI21_X1 i_0_657_709 (.A(n_0_657_625), .B1(n_0_445), .B2(n_0_657_627), 
      .ZN(n_0_657_624));
   AOI21_X1 i_0_657_710 (.A(n_0_657_959), .B1(n_0_657_627), .B2(n_0_657_626), 
      .ZN(n_0_657_625));
   INV_X1 i_0_657_711 (.A(n_911), .ZN(n_0_657_626));
   NAND2_X1 i_0_657_712 (.A1(n_0_182), .A2(n_0_657_964), .ZN(n_0_657_627));
   NAND2_X1 i_0_657_713 (.A1(n_0_657_628), .A2(n_0_657_631), .ZN(n_0_893));
   OAI21_X1 i_0_657_714 (.A(n_0_657_629), .B1(n_0_304), .B2(n_0_657_630), 
      .ZN(n_0_657_628));
   AOI21_X1 i_0_657_715 (.A(n_0_806), .B1(n_0_657_630), .B2(n_0_657_633), 
      .ZN(n_0_657_629));
   NAND2_X1 i_0_657_716 (.A1(n_0_730), .A2(n_0_657_964), .ZN(n_0_657_630));
   OAI21_X1 i_0_657_717 (.A(n_0_657_632), .B1(n_0_442), .B2(n_0_657_634), 
      .ZN(n_0_657_631));
   AOI21_X1 i_0_657_718 (.A(n_0_657_959), .B1(n_0_657_634), .B2(n_0_657_633), 
      .ZN(n_0_657_632));
   INV_X1 i_0_657_719 (.A(n_912), .ZN(n_0_657_633));
   NAND2_X1 i_0_657_720 (.A1(n_0_181), .A2(n_0_657_964), .ZN(n_0_657_634));
   NAND2_X1 i_0_657_721 (.A1(n_0_657_635), .A2(n_0_657_638), .ZN(n_0_894));
   OAI21_X1 i_0_657_722 (.A(n_0_657_636), .B1(n_0_303), .B2(n_0_657_637), 
      .ZN(n_0_657_635));
   AOI21_X1 i_0_657_723 (.A(n_0_806), .B1(n_0_657_637), .B2(n_0_657_640), 
      .ZN(n_0_657_636));
   NAND2_X1 i_0_657_724 (.A1(n_0_729), .A2(n_0_657_964), .ZN(n_0_657_637));
   OAI21_X1 i_0_657_725 (.A(n_0_657_639), .B1(n_0_439), .B2(n_0_657_641), 
      .ZN(n_0_657_638));
   AOI21_X1 i_0_657_726 (.A(n_0_657_959), .B1(n_0_657_641), .B2(n_0_657_640), 
      .ZN(n_0_657_639));
   INV_X1 i_0_657_727 (.A(n_913), .ZN(n_0_657_640));
   NAND2_X1 i_0_657_728 (.A1(n_0_180), .A2(n_0_657_964), .ZN(n_0_657_641));
   NAND2_X1 i_0_657_729 (.A1(n_0_657_647), .A2(n_0_657_642), .ZN(n_0_902));
   NAND3_X1 i_0_657_730 (.A1(n_0_657_645), .A2(n_0_657_643), .A3(n_0_657_959), 
      .ZN(n_0_657_642));
   OAI21_X1 i_0_657_731 (.A(n_0_657_652), .B1(n_0_657_644), .B2(n_0_657_813), 
      .ZN(n_0_657_643));
   INV_X1 i_0_657_732 (.A(n_0_728), .ZN(n_0_657_644));
   NAND3_X1 i_0_657_733 (.A1(n_0_657_646), .A2(n_0_728), .A3(n_0_657_964), 
      .ZN(n_0_657_645));
   INV_X1 i_0_657_734 (.A(n_0_302), .ZN(n_0_657_646));
   NAND3_X1 i_0_657_735 (.A1(n_0_657_650), .A2(n_0_806), .A3(n_0_657_648), 
      .ZN(n_0_657_647));
   NAND3_X1 i_0_657_736 (.A1(n_0_179), .A2(n_0_657_649), .A3(n_0_657_964), 
      .ZN(n_0_657_648));
   INV_X1 i_0_657_737 (.A(n_0_656), .ZN(n_0_657_649));
   NAND2_X1 i_0_657_738 (.A1(n_0_657_651), .A2(n_0_657_652), .ZN(n_0_657_650));
   NAND2_X1 i_0_657_739 (.A1(n_0_179), .A2(n_0_657_964), .ZN(n_0_657_651));
   INV_X1 i_0_657_740 (.A(n_914), .ZN(n_0_657_652));
   OAI21_X1 i_0_657_741 (.A(n_0_657_657), .B1(n_0_657_655), .B2(n_0_657_653), 
      .ZN(n_0_903));
   OAI21_X1 i_0_657_742 (.A(n_0_657_959), .B1(n_0_657_654), .B2(n_1002), 
      .ZN(n_0_657_653));
   INV_X1 i_0_657_743 (.A(n_0_657_656), .ZN(n_0_657_654));
   NOR2_X1 i_0_657_744 (.A1(n_0_301), .A2(n_0_657_656), .ZN(n_0_657_655));
   NAND2_X1 i_0_657_745 (.A1(n_0_727), .A2(n_0_657_964), .ZN(n_0_657_656));
   OAI21_X1 i_0_657_746 (.A(n_0_657_658), .B1(n_0_659), .B2(n_0_657_660), 
      .ZN(n_0_657_657));
   AOI21_X1 i_0_657_747 (.A(n_0_657_959), .B1(n_0_657_660), .B2(n_0_657_659), 
      .ZN(n_0_657_658));
   INV_X1 i_0_657_748 (.A(n_1002), .ZN(n_0_657_659));
   NAND2_X1 i_0_657_749 (.A1(n_0_178), .A2(n_0_657_964), .ZN(n_0_657_660));
   OAI21_X1 i_0_657_750 (.A(n_0_657_665), .B1(n_0_657_663), .B2(n_0_657_661), 
      .ZN(n_0_904));
   OAI21_X1 i_0_657_751 (.A(n_0_657_959), .B1(n_0_657_662), .B2(n_1003), 
      .ZN(n_0_657_661));
   INV_X1 i_0_657_752 (.A(n_0_657_664), .ZN(n_0_657_662));
   NOR2_X1 i_0_657_753 (.A1(n_0_300), .A2(n_0_657_664), .ZN(n_0_657_663));
   NAND2_X1 i_0_657_754 (.A1(n_0_726), .A2(n_0_657_964), .ZN(n_0_657_664));
   OAI21_X1 i_0_657_755 (.A(n_0_657_666), .B1(n_0_660), .B2(n_0_657_668), 
      .ZN(n_0_657_665));
   AOI21_X1 i_0_657_756 (.A(n_0_657_959), .B1(n_0_657_667), .B2(n_0_657_668), 
      .ZN(n_0_657_666));
   INV_X1 i_0_657_757 (.A(n_1003), .ZN(n_0_657_667));
   NAND2_X1 i_0_657_758 (.A1(n_0_177), .A2(n_0_657_964), .ZN(n_0_657_668));
   OAI21_X1 i_0_657_759 (.A(n_0_657_673), .B1(n_0_657_671), .B2(n_0_657_669), 
      .ZN(n_0_905));
   OAI21_X1 i_0_657_760 (.A(n_0_657_959), .B1(n_0_657_670), .B2(n_1004), 
      .ZN(n_0_657_669));
   INV_X1 i_0_657_761 (.A(n_0_657_672), .ZN(n_0_657_670));
   NOR2_X1 i_0_657_762 (.A1(n_0_299), .A2(n_0_657_672), .ZN(n_0_657_671));
   NAND2_X1 i_0_657_763 (.A1(n_0_725), .A2(n_0_657_964), .ZN(n_0_657_672));
   OAI21_X1 i_0_657_764 (.A(n_0_657_674), .B1(n_0_661), .B2(n_0_657_676), 
      .ZN(n_0_657_673));
   AOI21_X1 i_0_657_765 (.A(n_0_657_959), .B1(n_0_657_675), .B2(n_0_657_676), 
      .ZN(n_0_657_674));
   INV_X1 i_0_657_766 (.A(n_1004), .ZN(n_0_657_675));
   NAND2_X1 i_0_657_767 (.A1(n_0_176), .A2(n_0_657_964), .ZN(n_0_657_676));
   NAND2_X1 i_0_657_768 (.A1(n_0_657_677), .A2(n_0_657_680), .ZN(n_0_906));
   OAI21_X1 i_0_657_769 (.A(n_0_657_678), .B1(n_0_298), .B2(n_0_657_679), 
      .ZN(n_0_657_677));
   AOI21_X1 i_0_657_770 (.A(n_0_806), .B1(n_0_657_679), .B2(n_0_657_682), 
      .ZN(n_0_657_678));
   NAND2_X1 i_0_657_771 (.A1(n_0_724), .A2(n_0_657_964), .ZN(n_0_657_679));
   OAI21_X1 i_0_657_772 (.A(n_0_657_681), .B1(n_0_662), .B2(n_0_657_683), 
      .ZN(n_0_657_680));
   AOI21_X1 i_0_657_773 (.A(n_0_657_959), .B1(n_0_657_683), .B2(n_0_657_682), 
      .ZN(n_0_657_681));
   INV_X1 i_0_657_774 (.A(n_915), .ZN(n_0_657_682));
   NAND2_X1 i_0_657_775 (.A1(n_0_175), .A2(n_0_657_964), .ZN(n_0_657_683));
   OAI21_X1 i_0_657_776 (.A(n_0_657_688), .B1(n_0_657_686), .B2(n_0_657_684), 
      .ZN(n_0_907));
   OAI21_X1 i_0_657_777 (.A(n_0_657_959), .B1(n_0_657_685), .B2(n_1005), 
      .ZN(n_0_657_684));
   INV_X1 i_0_657_778 (.A(n_0_657_687), .ZN(n_0_657_685));
   NOR2_X1 i_0_657_779 (.A1(n_0_297), .A2(n_0_657_687), .ZN(n_0_657_686));
   NAND2_X1 i_0_657_780 (.A1(n_0_723), .A2(n_0_657_964), .ZN(n_0_657_687));
   OAI21_X1 i_0_657_781 (.A(n_0_657_689), .B1(n_0_436), .B2(n_0_657_691), 
      .ZN(n_0_657_688));
   AOI21_X1 i_0_657_782 (.A(n_0_657_959), .B1(n_0_657_691), .B2(n_0_657_690), 
      .ZN(n_0_657_689));
   INV_X1 i_0_657_783 (.A(n_1005), .ZN(n_0_657_690));
   NAND2_X1 i_0_657_784 (.A1(n_0_174), .A2(n_0_657_964), .ZN(n_0_657_691));
   OAI21_X1 i_0_657_785 (.A(n_0_657_696), .B1(n_0_657_694), .B2(n_0_657_692), 
      .ZN(n_0_908));
   OAI21_X1 i_0_657_786 (.A(n_0_657_959), .B1(n_0_657_693), .B2(n_1006), 
      .ZN(n_0_657_692));
   INV_X1 i_0_657_787 (.A(n_0_657_695), .ZN(n_0_657_693));
   NOR2_X1 i_0_657_788 (.A1(n_0_296), .A2(n_0_657_695), .ZN(n_0_657_694));
   NAND2_X1 i_0_657_789 (.A1(n_0_722), .A2(n_0_657_964), .ZN(n_0_657_695));
   OAI21_X1 i_0_657_790 (.A(n_0_657_697), .B1(n_0_434), .B2(n_0_657_699), 
      .ZN(n_0_657_696));
   AOI21_X1 i_0_657_791 (.A(n_0_657_959), .B1(n_0_657_698), .B2(n_0_657_699), 
      .ZN(n_0_657_697));
   INV_X1 i_0_657_792 (.A(n_1006), .ZN(n_0_657_698));
   NAND2_X1 i_0_657_793 (.A1(n_0_173), .A2(n_0_657_964), .ZN(n_0_657_699));
   OAI21_X1 i_0_657_794 (.A(n_0_657_704), .B1(n_0_657_702), .B2(n_0_657_700), 
      .ZN(n_0_909));
   OAI21_X1 i_0_657_795 (.A(n_0_657_959), .B1(n_0_657_701), .B2(n_1007), 
      .ZN(n_0_657_700));
   INV_X1 i_0_657_796 (.A(n_0_657_703), .ZN(n_0_657_701));
   NOR2_X1 i_0_657_797 (.A1(n_0_295), .A2(n_0_657_703), .ZN(n_0_657_702));
   NAND2_X1 i_0_657_798 (.A1(n_0_721), .A2(n_0_657_964), .ZN(n_0_657_703));
   OAI21_X1 i_0_657_799 (.A(n_0_657_705), .B1(n_0_431), .B2(n_0_657_707), 
      .ZN(n_0_657_704));
   AOI21_X1 i_0_657_800 (.A(n_0_657_959), .B1(n_0_657_707), .B2(n_0_657_706), 
      .ZN(n_0_657_705));
   INV_X1 i_0_657_801 (.A(n_1007), .ZN(n_0_657_706));
   NAND2_X1 i_0_657_802 (.A1(n_0_172), .A2(n_0_657_964), .ZN(n_0_657_707));
   OAI21_X1 i_0_657_803 (.A(n_0_657_712), .B1(n_0_657_710), .B2(n_0_657_708), 
      .ZN(n_0_910));
   OAI21_X1 i_0_657_804 (.A(n_0_657_959), .B1(n_0_657_709), .B2(n_1008), 
      .ZN(n_0_657_708));
   INV_X1 i_0_657_805 (.A(n_0_657_711), .ZN(n_0_657_709));
   NOR2_X1 i_0_657_806 (.A1(n_0_294), .A2(n_0_657_711), .ZN(n_0_657_710));
   NAND2_X1 i_0_657_807 (.A1(n_0_720), .A2(n_0_657_964), .ZN(n_0_657_711));
   OAI21_X1 i_0_657_808 (.A(n_0_657_713), .B1(n_0_663), .B2(n_0_657_715), 
      .ZN(n_0_657_712));
   AOI21_X1 i_0_657_809 (.A(n_0_657_959), .B1(n_0_657_714), .B2(n_0_657_715), 
      .ZN(n_0_657_713));
   INV_X1 i_0_657_810 (.A(n_1008), .ZN(n_0_657_714));
   NAND2_X1 i_0_657_811 (.A1(n_0_171), .A2(n_0_657_964), .ZN(n_0_657_715));
   NAND2_X1 i_0_657_812 (.A1(n_0_657_716), .A2(n_0_657_719), .ZN(n_0_912));
   OAI21_X1 i_0_657_813 (.A(n_0_657_717), .B1(n_0_292), .B2(n_0_657_718), 
      .ZN(n_0_657_716));
   AOI21_X1 i_0_657_814 (.A(n_0_806), .B1(n_0_657_718), .B2(n_0_657_721), 
      .ZN(n_0_657_717));
   NAND2_X1 i_0_657_815 (.A1(n_0_718), .A2(n_0_657_964), .ZN(n_0_657_718));
   OAI21_X1 i_0_657_816 (.A(n_0_657_720), .B1(n_0_425), .B2(n_0_657_722), 
      .ZN(n_0_657_719));
   AOI21_X1 i_0_657_817 (.A(n_0_657_959), .B1(n_0_657_722), .B2(n_0_657_721), 
      .ZN(n_0_657_720));
   INV_X1 i_0_657_818 (.A(n_916), .ZN(n_0_657_721));
   NAND2_X1 i_0_657_819 (.A1(n_0_169), .A2(n_0_657_964), .ZN(n_0_657_722));
   NAND2_X1 i_0_657_820 (.A1(n_0_657_723), .A2(n_0_657_726), .ZN(n_0_913));
   OAI21_X1 i_0_657_821 (.A(n_0_657_724), .B1(n_0_291), .B2(n_0_657_725), 
      .ZN(n_0_657_723));
   AOI21_X1 i_0_657_822 (.A(n_0_806), .B1(n_0_657_725), .B2(n_0_657_728), 
      .ZN(n_0_657_724));
   NAND2_X1 i_0_657_823 (.A1(n_0_717), .A2(n_0_657_964), .ZN(n_0_657_725));
   OAI21_X1 i_0_657_824 (.A(n_0_657_727), .B1(n_0_666), .B2(n_0_657_729), 
      .ZN(n_0_657_726));
   AOI21_X1 i_0_657_825 (.A(n_0_657_959), .B1(n_0_657_729), .B2(n_0_657_728), 
      .ZN(n_0_657_727));
   INV_X1 i_0_657_826 (.A(n_917), .ZN(n_0_657_728));
   NAND2_X1 i_0_657_827 (.A1(n_0_168), .A2(n_0_657_964), .ZN(n_0_657_729));
   NAND2_X1 i_0_657_828 (.A1(n_0_657_735), .A2(n_0_657_730), .ZN(n_0_914));
   NAND3_X1 i_0_657_829 (.A1(n_0_657_733), .A2(n_0_657_731), .A3(n_0_657_959), 
      .ZN(n_0_657_730));
   OAI21_X1 i_0_657_830 (.A(n_0_657_740), .B1(n_0_657_732), .B2(n_0_657_813), 
      .ZN(n_0_657_731));
   INV_X1 i_0_657_831 (.A(n_0_716), .ZN(n_0_657_732));
   NAND3_X1 i_0_657_832 (.A1(n_0_657_734), .A2(n_0_716), .A3(n_0_657_964), 
      .ZN(n_0_657_733));
   INV_X1 i_0_657_833 (.A(n_0_290), .ZN(n_0_657_734));
   NAND3_X1 i_0_657_834 (.A1(n_0_657_738), .A2(n_0_806), .A3(n_0_657_736), 
      .ZN(n_0_657_735));
   NAND3_X1 i_0_657_835 (.A1(n_0_167), .A2(n_0_657_737), .A3(n_0_657_964), 
      .ZN(n_0_657_736));
   INV_X1 i_0_657_836 (.A(n_0_422), .ZN(n_0_657_737));
   NAND2_X1 i_0_657_837 (.A1(n_0_657_739), .A2(n_0_657_740), .ZN(n_0_657_738));
   NAND2_X1 i_0_657_838 (.A1(n_0_167), .A2(n_0_657_964), .ZN(n_0_657_739));
   INV_X1 i_0_657_839 (.A(n_918), .ZN(n_0_657_740));
   NAND2_X1 i_0_657_840 (.A1(n_0_657_746), .A2(n_0_657_741), .ZN(n_0_915));
   NAND3_X1 i_0_657_841 (.A1(n_0_657_744), .A2(n_0_657_742), .A3(n_0_657_959), 
      .ZN(n_0_657_741));
   OAI21_X1 i_0_657_842 (.A(n_0_657_751), .B1(n_0_657_743), .B2(n_0_657_813), 
      .ZN(n_0_657_742));
   INV_X1 i_0_657_843 (.A(n_0_715), .ZN(n_0_657_743));
   NAND3_X1 i_0_657_844 (.A1(n_0_657_745), .A2(n_0_715), .A3(n_0_657_964), 
      .ZN(n_0_657_744));
   INV_X1 i_0_657_845 (.A(n_0_289), .ZN(n_0_657_745));
   NAND3_X1 i_0_657_846 (.A1(n_0_657_749), .A2(n_0_806), .A3(n_0_657_747), 
      .ZN(n_0_657_746));
   NAND3_X1 i_0_657_847 (.A1(n_0_166), .A2(n_0_657_748), .A3(n_0_657_964), 
      .ZN(n_0_657_747));
   INV_X1 i_0_657_848 (.A(n_0_419), .ZN(n_0_657_748));
   NAND2_X1 i_0_657_849 (.A1(n_0_657_750), .A2(n_0_657_751), .ZN(n_0_657_749));
   NAND2_X1 i_0_657_850 (.A1(n_0_166), .A2(n_0_657_964), .ZN(n_0_657_750));
   INV_X1 i_0_657_851 (.A(n_919), .ZN(n_0_657_751));
   NAND2_X1 i_0_657_852 (.A1(n_0_657_752), .A2(n_0_657_757), .ZN(n_0_916));
   NAND3_X1 i_0_657_853 (.A1(n_0_657_755), .A2(n_0_657_753), .A3(n_0_657_959), 
      .ZN(n_0_657_752));
   OAI21_X1 i_0_657_854 (.A(n_0_657_762), .B1(n_0_657_754), .B2(n_0_657_813), 
      .ZN(n_0_657_753));
   INV_X1 i_0_657_855 (.A(n_0_714), .ZN(n_0_657_754));
   NAND3_X1 i_0_657_856 (.A1(n_0_657_756), .A2(n_0_714), .A3(n_0_657_964), 
      .ZN(n_0_657_755));
   INV_X1 i_0_657_857 (.A(n_0_288), .ZN(n_0_657_756));
   NAND3_X1 i_0_657_858 (.A1(n_0_657_760), .A2(n_0_806), .A3(n_0_657_758), 
      .ZN(n_0_657_757));
   NAND3_X1 i_0_657_859 (.A1(n_0_165), .A2(n_0_657_759), .A3(n_0_657_964), 
      .ZN(n_0_657_758));
   INV_X1 i_0_657_860 (.A(n_0_416), .ZN(n_0_657_759));
   NAND2_X1 i_0_657_861 (.A1(n_0_657_761), .A2(n_0_657_762), .ZN(n_0_657_760));
   NAND2_X1 i_0_657_862 (.A1(n_0_165), .A2(n_0_657_964), .ZN(n_0_657_761));
   INV_X1 i_0_657_863 (.A(n_920), .ZN(n_0_657_762));
   NAND2_X1 i_0_657_864 (.A1(n_0_657_763), .A2(n_0_657_768), .ZN(n_0_917));
   NAND3_X1 i_0_657_865 (.A1(n_0_657_766), .A2(n_0_657_764), .A3(n_0_657_959), 
      .ZN(n_0_657_763));
   OAI21_X1 i_0_657_866 (.A(n_0_657_773), .B1(n_0_657_765), .B2(n_0_657_813), 
      .ZN(n_0_657_764));
   INV_X1 i_0_657_867 (.A(n_0_713), .ZN(n_0_657_765));
   NAND3_X1 i_0_657_868 (.A1(n_0_657_767), .A2(n_0_713), .A3(n_0_657_964), 
      .ZN(n_0_657_766));
   INV_X1 i_0_657_869 (.A(n_0_287), .ZN(n_0_657_767));
   NAND3_X1 i_0_657_870 (.A1(n_0_657_771), .A2(n_0_806), .A3(n_0_657_769), 
      .ZN(n_0_657_768));
   NAND3_X1 i_0_657_871 (.A1(n_0_164), .A2(n_0_657_770), .A3(n_0_657_964), 
      .ZN(n_0_657_769));
   INV_X1 i_0_657_872 (.A(n_0_413), .ZN(n_0_657_770));
   NAND2_X1 i_0_657_873 (.A1(n_0_657_772), .A2(n_0_657_773), .ZN(n_0_657_771));
   NAND2_X1 i_0_657_874 (.A1(n_0_164), .A2(n_0_657_964), .ZN(n_0_657_772));
   INV_X1 i_0_657_875 (.A(n_921), .ZN(n_0_657_773));
   NAND2_X1 i_0_657_876 (.A1(n_0_657_774), .A2(n_0_657_777), .ZN(n_0_918));
   OAI211_X1 i_0_657_877 (.A(n_0_657_775), .B(n_0_657_959), .C1(n_0_286), 
      .C2(n_0_657_776), .ZN(n_0_657_774));
   NAND2_X1 i_0_657_878 (.A1(n_0_657_776), .A2(n_0_657_779), .ZN(n_0_657_775));
   NAND2_X1 i_0_657_879 (.A1(n_0_710), .A2(n_0_657_964), .ZN(n_0_657_776));
   OAI21_X1 i_0_657_880 (.A(n_0_657_778), .B1(n_0_410), .B2(n_0_657_780), 
      .ZN(n_0_657_777));
   AOI21_X1 i_0_657_881 (.A(n_0_657_959), .B1(n_0_657_780), .B2(n_0_657_779), 
      .ZN(n_0_657_778));
   INV_X1 i_0_657_882 (.A(n_922), .ZN(n_0_657_779));
   NAND2_X1 i_0_657_883 (.A1(n_0_163), .A2(n_0_657_964), .ZN(n_0_657_780));
   NAND2_X1 i_0_657_884 (.A1(n_0_657_781), .A2(n_0_657_784), .ZN(n_0_919));
   OAI21_X1 i_0_657_885 (.A(n_0_657_782), .B1(n_0_285), .B2(n_0_657_783), 
      .ZN(n_0_657_781));
   AOI21_X1 i_0_657_886 (.A(n_0_806), .B1(n_0_657_783), .B2(n_0_657_786), 
      .ZN(n_0_657_782));
   NAND2_X1 i_0_657_887 (.A1(n_0_707), .A2(n_0_657_964), .ZN(n_0_657_783));
   OAI211_X1 i_0_657_888 (.A(n_0_657_785), .B(n_0_806), .C1(n_0_407), .C2(
      n_0_657_787), .ZN(n_0_657_784));
   NAND2_X1 i_0_657_889 (.A1(n_0_657_787), .A2(n_0_657_786), .ZN(n_0_657_785));
   INV_X1 i_0_657_890 (.A(n_923), .ZN(n_0_657_786));
   NAND2_X1 i_0_657_891 (.A1(n_0_162), .A2(n_0_657_964), .ZN(n_0_657_787));
   NAND2_X1 i_0_657_892 (.A1(n_0_657_788), .A2(n_0_657_791), .ZN(n_0_921));
   OAI21_X1 i_0_657_893 (.A(n_0_657_789), .B1(n_0_284), .B2(n_0_657_790), 
      .ZN(n_0_657_788));
   AOI21_X1 i_0_657_894 (.A(n_0_806), .B1(n_0_657_790), .B2(n_0_657_793), 
      .ZN(n_0_657_789));
   NAND2_X1 i_0_657_895 (.A1(n_0_706), .A2(n_0_657_964), .ZN(n_0_657_790));
   OAI21_X1 i_0_657_896 (.A(n_0_657_792), .B1(n_0_669), .B2(n_0_657_794), 
      .ZN(n_0_657_791));
   AOI21_X1 i_0_657_897 (.A(n_0_657_959), .B1(n_0_657_794), .B2(n_0_657_793), 
      .ZN(n_0_657_792));
   INV_X1 i_0_657_898 (.A(n_925), .ZN(n_0_657_793));
   NAND2_X1 i_0_657_899 (.A1(n_0_160), .A2(n_0_657_964), .ZN(n_0_657_794));
   NAND2_X1 i_0_657_900 (.A1(n_0_657_795), .A2(n_0_657_798), .ZN(n_0_923));
   OAI21_X1 i_0_657_901 (.A(n_0_657_796), .B1(n_0_282), .B2(n_0_657_797), 
      .ZN(n_0_657_795));
   AOI21_X1 i_0_657_902 (.A(n_0_806), .B1(n_0_657_797), .B2(n_0_657_800), 
      .ZN(n_0_657_796));
   NAND2_X1 i_0_657_903 (.A1(n_0_704), .A2(n_0_657_964), .ZN(n_0_657_797));
   OAI21_X1 i_0_657_904 (.A(n_0_657_799), .B1(n_0_402), .B2(n_0_657_801), 
      .ZN(n_0_657_798));
   AOI21_X1 i_0_657_905 (.A(n_0_657_959), .B1(n_0_657_801), .B2(n_0_657_800), 
      .ZN(n_0_657_799));
   INV_X1 i_0_657_906 (.A(n_926), .ZN(n_0_657_800));
   NAND2_X1 i_0_657_907 (.A1(n_0_158), .A2(n_0_657_964), .ZN(n_0_657_801));
   OAI21_X1 i_0_657_908 (.A(n_0_657_806), .B1(n_0_657_804), .B2(n_0_657_802), 
      .ZN(n_0_924));
   OAI21_X1 i_0_657_909 (.A(n_0_657_959), .B1(n_0_657_803), .B2(n_927), .ZN(
      n_0_657_802));
   INV_X1 i_0_657_910 (.A(n_0_657_805), .ZN(n_0_657_803));
   NOR2_X1 i_0_657_911 (.A1(n_0_281), .A2(n_0_657_805), .ZN(n_0_657_804));
   NAND2_X1 i_0_657_912 (.A1(n_0_703), .A2(n_0_657_964), .ZN(n_0_657_805));
   OAI211_X1 i_0_657_913 (.A(n_0_657_807), .B(n_0_806), .C1(n_927), .C2(
      n_0_657_809), .ZN(n_0_657_806));
   NAND2_X1 i_0_657_914 (.A1(n_0_657_808), .A2(n_0_657_809), .ZN(n_0_657_807));
   INV_X1 i_0_657_915 (.A(n_0_671), .ZN(n_0_657_808));
   INV_X1 i_0_657_916 (.A(n_0_657_810), .ZN(n_0_657_809));
   NAND2_X1 i_0_657_917 (.A1(n_0_157), .A2(n_0_657_964), .ZN(n_0_657_810));
   NAND2_X1 i_0_657_918 (.A1(n_0_657_811), .A2(n_0_657_817), .ZN(n_0_925));
   NAND3_X1 i_0_657_919 (.A1(n_0_657_812), .A2(n_0_657_959), .A3(n_0_657_815), 
      .ZN(n_0_657_811));
   OAI21_X1 i_0_657_920 (.A(n_0_657_819), .B1(n_0_657_814), .B2(n_0_657_813), 
      .ZN(n_0_657_812));
   INV_X1 i_0_657_921 (.A(n_0_657_964), .ZN(n_0_657_813));
   INV_X1 i_0_657_922 (.A(n_0_700), .ZN(n_0_657_814));
   NAND3_X1 i_0_657_923 (.A1(n_0_700), .A2(n_0_657_816), .A3(n_0_657_964), 
      .ZN(n_0_657_815));
   INV_X1 i_0_657_924 (.A(n_0_280), .ZN(n_0_657_816));
   OAI21_X1 i_0_657_925 (.A(n_0_657_818), .B1(n_0_399), .B2(n_0_657_820), 
      .ZN(n_0_657_817));
   AOI21_X1 i_0_657_926 (.A(n_0_657_959), .B1(n_0_657_820), .B2(n_0_657_819), 
      .ZN(n_0_657_818));
   INV_X1 i_0_657_927 (.A(n_928), .ZN(n_0_657_819));
   NAND2_X1 i_0_657_928 (.A1(n_0_156), .A2(n_0_657_964), .ZN(n_0_657_820));
   NAND2_X1 i_0_657_929 (.A1(n_0_657_821), .A2(n_0_657_824), .ZN(n_0_926));
   OAI21_X1 i_0_657_930 (.A(n_0_657_822), .B1(n_0_279), .B2(n_0_657_823), 
      .ZN(n_0_657_821));
   AOI21_X1 i_0_657_931 (.A(n_0_806), .B1(n_0_657_823), .B2(n_0_657_826), 
      .ZN(n_0_657_822));
   NAND2_X1 i_0_657_932 (.A1(n_0_699), .A2(n_0_657_964), .ZN(n_0_657_823));
   OAI211_X1 i_0_657_933 (.A(n_0_657_825), .B(n_0_806), .C1(n_1269), .C2(
      n_0_657_827), .ZN(n_0_657_824));
   NAND2_X1 i_0_657_934 (.A1(n_0_657_827), .A2(n_0_657_826), .ZN(n_0_657_825));
   INV_X1 i_0_657_935 (.A(n_929), .ZN(n_0_657_826));
   NAND2_X1 i_0_657_936 (.A1(n_0_155), .A2(n_0_657_964), .ZN(n_0_657_827));
   NAND2_X1 i_0_657_937 (.A1(n_0_657_828), .A2(n_0_657_831), .ZN(n_0_927));
   OAI21_X1 i_0_657_938 (.A(n_0_657_829), .B1(n_0_278), .B2(n_0_657_830), 
      .ZN(n_0_657_828));
   AOI21_X1 i_0_657_939 (.A(n_0_806), .B1(n_0_657_830), .B2(n_0_657_833), 
      .ZN(n_0_657_829));
   NAND2_X1 i_0_657_940 (.A1(n_0_698), .A2(n_0_657_964), .ZN(n_0_657_830));
   OAI21_X1 i_0_657_941 (.A(n_0_657_832), .B1(n_0_396), .B2(n_0_657_834), 
      .ZN(n_0_657_831));
   AOI21_X1 i_0_657_942 (.A(n_0_657_959), .B1(n_0_657_834), .B2(n_0_657_833), 
      .ZN(n_0_657_832));
   INV_X1 i_0_657_943 (.A(n_930), .ZN(n_0_657_833));
   NAND2_X1 i_0_657_944 (.A1(n_0_154), .A2(n_0_657_964), .ZN(n_0_657_834));
   NAND2_X1 i_0_657_945 (.A1(n_0_657_835), .A2(n_0_657_838), .ZN(n_0_928));
   OAI21_X1 i_0_657_946 (.A(n_0_657_836), .B1(n_0_277), .B2(n_0_657_837), 
      .ZN(n_0_657_835));
   AOI21_X1 i_0_657_947 (.A(n_0_806), .B1(n_0_657_837), .B2(n_0_657_840), 
      .ZN(n_0_657_836));
   NAND2_X1 i_0_657_948 (.A1(n_0_697), .A2(n_0_657_964), .ZN(n_0_657_837));
   OAI211_X1 i_0_657_949 (.A(n_0_657_839), .B(n_0_806), .C1(n_0_394), .C2(
      n_0_657_841), .ZN(n_0_657_838));
   NAND2_X1 i_0_657_950 (.A1(n_0_657_841), .A2(n_0_657_840), .ZN(n_0_657_839));
   INV_X1 i_0_657_951 (.A(n_931), .ZN(n_0_657_840));
   NAND2_X1 i_0_657_952 (.A1(n_0_153), .A2(n_0_657_964), .ZN(n_0_657_841));
   NAND2_X1 i_0_657_953 (.A1(n_0_657_842), .A2(n_0_657_845), .ZN(n_0_929));
   OAI21_X1 i_0_657_954 (.A(n_0_657_843), .B1(n_0_276), .B2(n_0_657_844), 
      .ZN(n_0_657_842));
   AOI21_X1 i_0_657_955 (.A(n_0_806), .B1(n_0_657_844), .B2(n_0_657_847), 
      .ZN(n_0_657_843));
   NAND2_X1 i_0_657_956 (.A1(n_0_696), .A2(n_0_657_964), .ZN(n_0_657_844));
   OAI21_X1 i_0_657_957 (.A(n_0_657_846), .B1(n_0_391), .B2(n_0_657_848), 
      .ZN(n_0_657_845));
   AOI21_X1 i_0_657_958 (.A(n_0_657_959), .B1(n_0_657_848), .B2(n_0_657_847), 
      .ZN(n_0_657_846));
   INV_X1 i_0_657_959 (.A(n_932), .ZN(n_0_657_847));
   NAND2_X1 i_0_657_960 (.A1(n_0_152), .A2(n_0_657_964), .ZN(n_0_657_848));
   NAND2_X1 i_0_657_961 (.A1(n_0_657_849), .A2(n_0_657_852), .ZN(n_0_930));
   OAI21_X1 i_0_657_962 (.A(n_0_657_850), .B1(n_0_275), .B2(n_0_657_851), 
      .ZN(n_0_657_849));
   AOI21_X1 i_0_657_963 (.A(n_0_806), .B1(n_0_657_851), .B2(n_0_657_854), 
      .ZN(n_0_657_850));
   NAND2_X1 i_0_657_964 (.A1(n_0_695), .A2(n_0_657_964), .ZN(n_0_657_851));
   OAI21_X1 i_0_657_965 (.A(n_0_657_853), .B1(n_0_389), .B2(n_0_657_855), 
      .ZN(n_0_657_852));
   AOI21_X1 i_0_657_966 (.A(n_0_657_959), .B1(n_0_657_855), .B2(n_0_657_854), 
      .ZN(n_0_657_853));
   INV_X1 i_0_657_967 (.A(n_933), .ZN(n_0_657_854));
   NAND2_X1 i_0_657_968 (.A1(n_0_151), .A2(n_0_657_964), .ZN(n_0_657_855));
   NAND2_X1 i_0_657_969 (.A1(n_0_657_856), .A2(n_0_657_859), .ZN(n_0_931));
   OAI21_X1 i_0_657_970 (.A(n_0_657_857), .B1(n_0_274), .B2(n_0_657_858), 
      .ZN(n_0_657_856));
   AOI21_X1 i_0_657_971 (.A(n_0_806), .B1(n_0_657_858), .B2(n_0_657_861), 
      .ZN(n_0_657_857));
   NAND2_X1 i_0_657_972 (.A1(n_0_694), .A2(n_0_657_964), .ZN(n_0_657_858));
   OAI211_X1 i_0_657_973 (.A(n_0_657_860), .B(n_0_806), .C1(n_0_388), .C2(
      n_0_657_862), .ZN(n_0_657_859));
   NAND2_X1 i_0_657_974 (.A1(n_0_657_862), .A2(n_0_657_861), .ZN(n_0_657_860));
   INV_X1 i_0_657_975 (.A(n_934), .ZN(n_0_657_861));
   NAND2_X1 i_0_657_976 (.A1(n_0_150), .A2(n_0_657_964), .ZN(n_0_657_862));
   NAND2_X1 i_0_657_977 (.A1(n_0_657_863), .A2(n_0_657_866), .ZN(n_0_932));
   OAI21_X1 i_0_657_978 (.A(n_0_657_864), .B1(n_0_273), .B2(n_0_657_865), 
      .ZN(n_0_657_863));
   AOI21_X1 i_0_657_979 (.A(n_0_806), .B1(n_0_657_865), .B2(n_0_657_868), 
      .ZN(n_0_657_864));
   NAND2_X1 i_0_657_980 (.A1(n_0_693), .A2(n_0_657_964), .ZN(n_0_657_865));
   OAI211_X1 i_0_657_981 (.A(n_0_657_867), .B(n_0_806), .C1(n_0_387), .C2(
      n_0_657_869), .ZN(n_0_657_866));
   NAND2_X1 i_0_657_982 (.A1(n_0_657_869), .A2(n_0_657_868), .ZN(n_0_657_867));
   INV_X1 i_0_657_983 (.A(n_935), .ZN(n_0_657_868));
   NAND2_X1 i_0_657_984 (.A1(n_0_149), .A2(n_0_657_964), .ZN(n_0_657_869));
   NAND2_X1 i_0_657_985 (.A1(n_0_657_870), .A2(n_0_657_873), .ZN(n_0_933));
   OAI21_X1 i_0_657_986 (.A(n_0_657_871), .B1(n_0_272), .B2(n_0_657_872), 
      .ZN(n_0_657_870));
   AOI21_X1 i_0_657_987 (.A(n_0_806), .B1(n_0_657_872), .B2(n_0_657_875), 
      .ZN(n_0_657_871));
   NAND2_X1 i_0_657_988 (.A1(n_0_692), .A2(n_0_657_964), .ZN(n_0_657_872));
   OAI21_X1 i_0_657_989 (.A(n_0_657_874), .B1(n_0_674), .B2(n_0_657_876), 
      .ZN(n_0_657_873));
   AOI21_X1 i_0_657_990 (.A(n_0_657_959), .B1(n_0_657_876), .B2(n_0_657_875), 
      .ZN(n_0_657_874));
   INV_X1 i_0_657_991 (.A(n_936), .ZN(n_0_657_875));
   NAND2_X1 i_0_657_992 (.A1(n_0_148), .A2(n_0_657_964), .ZN(n_0_657_876));
   NAND2_X1 i_0_657_993 (.A1(n_0_657_877), .A2(n_0_657_878), .ZN(n_0_935));
   OAI221_X1 i_0_657_994 (.A(n_0_806), .B1(n_0_657_53), .B2(n_0_810), .C1(n_951), 
      .C2(n_0_657_52), .ZN(n_0_657_877));
   OAI21_X1 i_0_657_995 (.A(n_0_657_879), .B1(n_1282), .B2(n_0_657_881), 
      .ZN(n_0_657_878));
   AOI21_X1 i_0_657_996 (.A(n_0_806), .B1(n_0_657_881), .B2(n_0_657_880), 
      .ZN(n_0_657_879));
   INV_X1 i_0_657_997 (.A(n_951), .ZN(n_0_657_880));
   NAND2_X1 i_0_657_998 (.A1(n_1288), .A2(n_0_657_964), .ZN(n_0_657_881));
   NAND2_X1 i_0_657_999 (.A1(n_0_657_882), .A2(n_0_657_885), .ZN(n_0_936));
   OAI21_X1 i_0_657_1000 (.A(n_0_657_883), .B1(n_0_271), .B2(n_0_657_884), 
      .ZN(n_0_657_882));
   AOI21_X1 i_0_657_1001 (.A(n_0_806), .B1(n_0_657_884), .B2(n_0_657_887), 
      .ZN(n_0_657_883));
   NAND2_X1 i_0_657_1002 (.A1(n_0_691), .A2(n_0_657_964), .ZN(n_0_657_884));
   OAI211_X1 i_0_657_1003 (.A(n_0_657_886), .B(n_0_806), .C1(n_0_675), .C2(
      n_0_657_888), .ZN(n_0_657_885));
   NAND2_X1 i_0_657_1004 (.A1(n_0_657_888), .A2(n_0_657_887), .ZN(n_0_657_886));
   INV_X1 i_0_657_1005 (.A(n_978), .ZN(n_0_657_887));
   NAND2_X1 i_0_657_1006 (.A1(n_0_145), .A2(n_0_657_964), .ZN(n_0_657_888));
   NAND2_X1 i_0_657_1007 (.A1(n_0_657_889), .A2(n_0_657_895), .ZN(n_0_937));
   NAND3_X1 i_0_657_1008 (.A1(n_0_657_891), .A2(n_0_657_959), .A3(n_0_657_890), 
      .ZN(n_0_657_889));
   NAND2_X1 i_0_657_1009 (.A1(n_0_657_893), .A2(n_0_657_897), .ZN(n_0_657_890));
   NAND2_X1 i_0_657_1010 (.A1(n_0_657_892), .A2(n_0_657_894), .ZN(n_0_657_891));
   INV_X1 i_0_657_1011 (.A(n_0_657_893), .ZN(n_0_657_892));
   NAND2_X1 i_0_657_1012 (.A1(n_0_690), .A2(n_0_657_964), .ZN(n_0_657_893));
   INV_X1 i_0_657_1013 (.A(n_0_270), .ZN(n_0_657_894));
   OAI211_X1 i_0_657_1014 (.A(n_0_657_896), .B(n_0_806), .C1(n_0_386), .C2(
      n_0_657_898), .ZN(n_0_657_895));
   NAND2_X1 i_0_657_1015 (.A1(n_0_657_898), .A2(n_0_657_897), .ZN(n_0_657_896));
   INV_X1 i_0_657_1016 (.A(n_938), .ZN(n_0_657_897));
   NAND2_X1 i_0_657_1017 (.A1(n_0_144), .A2(n_0_657_964), .ZN(n_0_657_898));
   NAND2_X1 i_0_657_1018 (.A1(n_0_657_899), .A2(n_0_657_900), .ZN(n_0_938));
   OAI221_X1 i_0_657_1019 (.A(n_0_806), .B1(n_0_657_55), .B2(n_0_385), .C1(n_939), 
      .C2(n_0_657_54), .ZN(n_0_657_899));
   OAI21_X1 i_0_657_1020 (.A(n_0_657_901), .B1(n_1212), .B2(n_0_657_903), 
      .ZN(n_0_657_900));
   AOI21_X1 i_0_657_1021 (.A(n_0_806), .B1(n_0_657_903), .B2(n_0_657_902), 
      .ZN(n_0_657_901));
   INV_X1 i_0_657_1022 (.A(n_939), .ZN(n_0_657_902));
   NAND2_X1 i_0_657_1023 (.A1(n_1088), .A2(n_0_657_964), .ZN(n_0_657_903));
   NAND2_X1 i_0_657_1024 (.A1(n_0_657_904), .A2(n_0_657_910), .ZN(n_0_940));
   NAND3_X1 i_0_657_1025 (.A1(n_0_657_906), .A2(n_0_657_959), .A3(n_0_657_905), 
      .ZN(n_0_657_904));
   NAND2_X1 i_0_657_1026 (.A1(n_0_657_908), .A2(n_0_657_912), .ZN(n_0_657_905));
   NAND2_X1 i_0_657_1027 (.A1(n_0_657_907), .A2(n_0_657_909), .ZN(n_0_657_906));
   INV_X1 i_0_657_1028 (.A(n_0_657_908), .ZN(n_0_657_907));
   NAND2_X1 i_0_657_1029 (.A1(n_0_687), .A2(n_0_657_964), .ZN(n_0_657_908));
   INV_X1 i_0_657_1030 (.A(n_0_269), .ZN(n_0_657_909));
   OAI211_X1 i_0_657_1031 (.A(n_0_657_911), .B(n_0_806), .C1(n_0_384), .C2(
      n_0_657_913), .ZN(n_0_657_910));
   NAND2_X1 i_0_657_1032 (.A1(n_0_657_913), .A2(n_0_657_912), .ZN(n_0_657_911));
   INV_X1 i_0_657_1033 (.A(n_941), .ZN(n_0_657_912));
   NAND2_X1 i_0_657_1034 (.A1(n_0_141), .A2(n_0_657_964), .ZN(n_0_657_913));
   NAND2_X1 i_0_657_1035 (.A1(n_0_657_914), .A2(n_0_657_917), .ZN(n_0_942));
   OAI21_X1 i_0_657_1036 (.A(n_0_657_915), .B1(n_0_268), .B2(n_0_657_916), 
      .ZN(n_0_657_914));
   AOI21_X1 i_0_657_1037 (.A(n_0_806), .B1(n_0_657_916), .B2(n_0_657_919), 
      .ZN(n_0_657_915));
   NAND2_X1 i_0_657_1038 (.A1(n_1305), .A2(n_0_657_964), .ZN(n_0_657_916));
   OAI211_X1 i_0_657_1039 (.A(n_0_657_918), .B(n_0_806), .C1(n_0_813), .C2(
      n_0_657_920), .ZN(n_0_657_917));
   NAND2_X1 i_0_657_1040 (.A1(n_0_657_920), .A2(n_0_657_919), .ZN(n_0_657_918));
   INV_X1 i_0_657_1041 (.A(n_943), .ZN(n_0_657_919));
   NAND2_X1 i_0_657_1042 (.A1(n_0_139), .A2(n_0_657_964), .ZN(n_0_657_920));
   NAND2_X1 i_0_657_1043 (.A1(n_0_657_921), .A2(n_0_657_924), .ZN(n_0_943));
   OAI21_X1 i_0_657_1044 (.A(n_0_657_922), .B1(n_0_267), .B2(n_0_657_923), 
      .ZN(n_0_657_921));
   AOI21_X1 i_0_657_1045 (.A(n_0_806), .B1(n_0_657_923), .B2(n_0_657_926), 
      .ZN(n_0_657_922));
   NAND2_X1 i_0_657_1046 (.A1(n_1306), .A2(n_0_657_964), .ZN(n_0_657_923));
   OAI211_X1 i_0_657_1047 (.A(n_0_657_925), .B(n_0_806), .C1(n_0_814), .C2(
      n_0_657_927), .ZN(n_0_657_924));
   NAND2_X1 i_0_657_1048 (.A1(n_0_657_927), .A2(n_0_657_926), .ZN(n_0_657_925));
   INV_X1 i_0_657_1049 (.A(n_944), .ZN(n_0_657_926));
   NAND2_X1 i_0_657_1050 (.A1(n_0_138), .A2(n_0_657_964), .ZN(n_0_657_927));
   NAND2_X1 i_0_657_1051 (.A1(n_0_657_928), .A2(n_0_657_931), .ZN(n_0_944));
   OAI21_X1 i_0_657_1052 (.A(n_0_657_929), .B1(n_0_266), .B2(n_0_657_930), 
      .ZN(n_0_657_928));
   AOI21_X1 i_0_657_1053 (.A(n_0_806), .B1(n_0_657_930), .B2(n_0_657_933), 
      .ZN(n_0_657_929));
   NAND2_X1 i_0_657_1054 (.A1(n_0_686), .A2(n_0_657_964), .ZN(n_0_657_930));
   OAI21_X1 i_0_657_1055 (.A(n_0_657_932), .B1(n_0_383), .B2(n_0_657_934), 
      .ZN(n_0_657_931));
   AOI21_X1 i_0_657_1056 (.A(n_0_657_959), .B1(n_0_657_934), .B2(n_0_657_933), 
      .ZN(n_0_657_932));
   INV_X1 i_0_657_1057 (.A(n_945), .ZN(n_0_657_933));
   NAND2_X1 i_0_657_1058 (.A1(n_0_137), .A2(n_0_657_964), .ZN(n_0_657_934));
   NAND2_X1 i_0_657_1059 (.A1(n_0_657_935), .A2(n_0_657_938), .ZN(n_0_946));
   OAI21_X1 i_0_657_1060 (.A(n_0_657_936), .B1(n_0_265), .B2(n_0_657_937), 
      .ZN(n_0_657_935));
   AOI21_X1 i_0_657_1061 (.A(n_0_806), .B1(n_0_657_937), .B2(n_0_657_940), 
      .ZN(n_0_657_936));
   NAND2_X1 i_0_657_1062 (.A1(n_0_685), .A2(n_0_657_964), .ZN(n_0_657_937));
   OAI21_X1 i_0_657_1063 (.A(n_0_657_939), .B1(n_0_382), .B2(n_0_657_941), 
      .ZN(n_0_657_938));
   AOI21_X1 i_0_657_1064 (.A(n_0_657_959), .B1(n_0_657_941), .B2(n_0_657_940), 
      .ZN(n_0_657_939));
   INV_X1 i_0_657_1065 (.A(n_947), .ZN(n_0_657_940));
   NAND2_X1 i_0_657_1066 (.A1(n_0_135), .A2(n_0_657_964), .ZN(n_0_657_941));
   OAI21_X1 i_0_657_1067 (.A(n_0_657_942), .B1(n_0_806), .B2(n_0_657_946), 
      .ZN(n_0_947));
   OAI21_X1 i_0_657_1068 (.A(n_0_657_943), .B1(n_0_676), .B2(n_0_657_945), 
      .ZN(n_0_657_942));
   AOI21_X1 i_0_657_1069 (.A(n_0_657_959), .B1(n_0_657_944), .B2(n_0_657_945), 
      .ZN(n_0_657_943));
   INV_X1 i_0_657_1070 (.A(n_1010), .ZN(n_0_657_944));
   NAND2_X1 i_0_657_1071 (.A1(n_0_134), .A2(n_0_657_964), .ZN(n_0_657_945));
   AOI22_X1 i_0_657_1072 (.A1(n_0_264), .A2(n_0_657_74), .B1(n_0_657_75), 
      .B2(n_1010), .ZN(n_0_657_946));
   NAND2_X1 i_0_657_1073 (.A1(n_0_657_947), .A2(n_0_657_952), .ZN(n_0_948));
   NAND3_X1 i_0_657_1074 (.A1(n_0_657_948), .A2(n_0_657_959), .A3(n_0_657_950), 
      .ZN(n_0_657_947));
   NAND2_X1 i_0_657_1075 (.A1(n_0_657_949), .A2(n_0_657_954), .ZN(n_0_657_948));
   NAND2_X1 i_0_657_1076 (.A1(n_0_679), .A2(n_0_657_964), .ZN(n_0_657_949));
   NAND3_X1 i_0_657_1077 (.A1(n_0_679), .A2(n_0_657_951), .A3(n_0_657_964), 
      .ZN(n_0_657_950));
   INV_X1 i_0_657_1078 (.A(n_0_263), .ZN(n_0_657_951));
   OAI211_X1 i_0_657_1079 (.A(n_0_657_953), .B(n_0_806), .C1(n_0_381), .C2(
      n_0_657_955), .ZN(n_0_657_952));
   NAND2_X1 i_0_657_1080 (.A1(n_0_657_955), .A2(n_0_657_954), .ZN(n_0_657_953));
   INV_X1 i_0_657_1081 (.A(n_948), .ZN(n_0_657_954));
   NAND2_X1 i_0_657_1082 (.A1(n_0_133), .A2(n_0_657_964), .ZN(n_0_657_955));
   NAND2_X1 i_0_657_1083 (.A1(n_0_657_956), .A2(n_0_657_960), .ZN(n_0_949));
   OAI211_X1 i_0_657_1084 (.A(n_0_657_957), .B(n_0_657_959), .C1(n_0_259), 
      .C2(n_0_657_958), .ZN(n_0_657_956));
   NAND2_X1 i_0_657_1085 (.A1(n_0_657_958), .A2(n_0_657_962), .ZN(n_0_657_957));
   NAND2_X1 i_0_657_1086 (.A1(n_0_260), .A2(n_0_657_964), .ZN(n_0_657_958));
   INV_X1 i_0_657_1087 (.A(n_0_806), .ZN(n_0_657_959));
   OAI211_X1 i_0_657_1088 (.A(n_0_657_961), .B(n_0_806), .C1(n_0_128), .C2(
      n_0_657_963), .ZN(n_0_657_960));
   NAND2_X1 i_0_657_1089 (.A1(n_0_657_963), .A2(n_0_657_962), .ZN(n_0_657_961));
   INV_X1 i_0_657_1090 (.A(n_949), .ZN(n_0_657_962));
   NAND2_X1 i_0_657_1091 (.A1(n_0_132), .A2(n_0_657_964), .ZN(n_0_657_963));
   NOR2_X1 i_0_657_1092 (.A1(n_0_657_78), .A2(rst), .ZN(n_0_657_964));
   DFF_X1 \buf_reg[118]  (.D(n_0_825), .CK(clk), .Q(n_987), .QN());
   DFF_X1 \buf_reg[115]  (.D(n_0_828), .CK(clk), .Q(n_988), .QN());
   DFF_X1 \buf_reg[102]  (.D(n_0_841), .CK(clk), .Q(n_989), .QN());
   DFF_X1 \buf_reg[96]  (.D(n_0_847), .CK(clk), .Q(n_990), .QN());
   DFF_X1 \buf_reg[88]  (.D(n_0_855), .CK(clk), .Q(n_991), .QN());
   DFF_X1 \buf_reg[86]  (.D(n_0_857), .CK(clk), .Q(n_992), .QN());
   DFF_X1 \buf_reg[82]  (.D(n_0_861), .CK(clk), .Q(n_993), .QN());
   DFF_X1 \buf_reg[75]  (.D(n_0_868), .CK(clk), .Q(n_994), .QN());
   DFF_X1 \buf_reg[74]  (.D(n_0_869), .CK(clk), .Q(n_995), .QN());
   DFF_X1 \buf_reg[73]  (.D(n_0_870), .CK(clk), .Q(n_996), .QN());
   DFF_X1 \buf_reg[72]  (.D(n_0_871), .CK(clk), .Q(n_997), .QN());
   DFF_X1 \buf_reg[58]  (.D(n_0_885), .CK(clk), .Q(n_998), .QN());
   DFF_X1 \buf_reg[55]  (.D(n_0_888), .CK(clk), .Q(n_999), .QN());
   DFF_X1 \buf_reg[53]  (.D(n_0_890), .CK(clk), .Q(n_1000), .QN());
   DFF_X1 \buf_reg[52]  (.D(n_0_891), .CK(clk), .Q(n_1001), .QN());
   DFF_X1 \buf_reg[47]  (.D(n_0_903), .CK(clk), .Q(n_1002), .QN());
   DFF_X1 \buf_reg[46]  (.D(n_0_904), .CK(clk), .Q(n_1003), .QN());
   DFF_X1 \buf_reg[45]  (.D(n_0_905), .CK(clk), .Q(n_1004), .QN());
   DFF_X1 \buf_reg[43]  (.D(n_0_907), .CK(clk), .Q(n_1005), .QN());
   DFF_X1 \buf_reg[42]  (.D(n_0_908), .CK(clk), .Q(n_1006), .QN());
   DFF_X1 \buf_reg[41]  (.D(n_0_909), .CK(clk), .Q(n_1007), .QN());
   DFF_X1 \buf_reg[40]  (.D(n_0_910), .CK(clk), .Q(n_1008), .QN());
   DFF_X1 \buf_reg[56]  (.D(n_0_887), .CK(clk), .Q(n_1009), .QN());
   DFF_X1 \buf_reg[3]  (.D(n_0_947), .CK(clk), .Q(n_1010), .QN());
   BUF_X1 rt_shieldBuf__8 (.A(n_1089), .Z(n_1011));
   OAI21_X1 i_2_0_0 (.A(n_2_0_0), .B1(n_952), .B2(n_2_0_1), .ZN(n_1012));
   AOI21_X1 i_2_0_1 (.A(n_2_1), .B1(n_952), .B2(n_2_2), .ZN(n_2_0_0));
   INV_X1 i_2_0_2 (.A(n_2_3), .ZN(n_2_0_1));
   OAI21_X1 i_2_1_0 (.A(n_2_1_0), .B1(n_952), .B2(n_2_1_1), .ZN(n_1013));
   AOI21_X1 i_2_1_1 (.A(n_2_4), .B1(n_952), .B2(n_1199), .ZN(n_2_1_0));
   INV_X1 i_2_1_2 (.A(n_1200), .ZN(n_2_1_1));
   OAI21_X1 i_2_2_0 (.A(n_2_2_0), .B1(n_952), .B2(n_2_2_1), .ZN(n_1014));
   AOI21_X1 i_2_2_1 (.A(n_2_5), .B1(n_952), .B2(n_2_6), .ZN(n_2_2_0));
   INV_X1 i_2_2_2 (.A(n_2_7), .ZN(n_2_2_1));
   OAI21_X1 i_2_3_0 (.A(n_2_3_0), .B1(n_952), .B2(n_2_3_1), .ZN(n_1015));
   AOI21_X1 i_2_3_1 (.A(n_2_17), .B1(n_952), .B2(n_2_18), .ZN(n_2_3_0));
   INV_X1 i_2_3_2 (.A(n_2_19), .ZN(n_2_3_1));
   OAI21_X1 i_2_4_0 (.A(n_2_4_0), .B1(n_952), .B2(n_2_4_1), .ZN(n_1016));
   AOI21_X1 i_2_4_1 (.A(n_2_21), .B1(n_952), .B2(n_1201), .ZN(n_2_4_0));
   INV_X1 i_2_4_2 (.A(n_1202), .ZN(n_2_4_1));
   OAI21_X1 i_2_5_0 (.A(n_2_5_0), .B1(n_952), .B2(n_2_5_1), .ZN(n_1017));
   AOI21_X1 i_2_5_1 (.A(n_2_22), .B1(n_952), .B2(n_2_23), .ZN(n_2_5_0));
   INV_X1 i_2_5_2 (.A(n_2_24), .ZN(n_2_5_1));
   OAI21_X1 i_2_6_0 (.A(n_2_6_0), .B1(n_952), .B2(n_2_6_1), .ZN(n_1018));
   AOI21_X1 i_2_6_1 (.A(n_2_28), .B1(n_952), .B2(n_2_29), .ZN(n_2_6_0));
   INV_X1 i_2_6_2 (.A(n_2_30), .ZN(n_2_6_1));
   OAI21_X1 i_2_7_0 (.A(n_2_7_0), .B1(n_952), .B2(n_2_7_1), .ZN(n_1019));
   AOI21_X1 i_2_7_1 (.A(n_2_38), .B1(n_952), .B2(n_2_39), .ZN(n_2_7_0));
   INV_X1 i_2_7_2 (.A(n_2_40), .ZN(n_2_7_1));
   OAI21_X1 i_2_8_0 (.A(n_2_8_0), .B1(n_952), .B2(n_2_8_1), .ZN(n_1020));
   AOI21_X1 i_2_8_1 (.A(n_2_50), .B1(n_952), .B2(n_2_51), .ZN(n_2_8_0));
   INV_X1 i_2_8_2 (.A(n_2_52), .ZN(n_2_8_1));
   OAI21_X1 i_2_9_0 (.A(n_2_9_0), .B1(n_952), .B2(n_2_9_1), .ZN(n_1021));
   AOI21_X1 i_2_9_1 (.A(n_2_53), .B1(n_952), .B2(n_2_54), .ZN(n_2_9_0));
   INV_X1 i_2_9_2 (.A(n_2_55), .ZN(n_2_9_1));
   OAI21_X1 i_2_10_0 (.A(n_2_10_0), .B1(n_952), .B2(n_2_10_1), .ZN(n_1022));
   AOI21_X1 i_2_10_1 (.A(n_2_56), .B1(n_952), .B2(n_2_57), .ZN(n_2_10_0));
   INV_X1 i_2_10_2 (.A(n_2_58), .ZN(n_2_10_1));
   OAI21_X1 i_2_11_0 (.A(n_2_11_0), .B1(n_952), .B2(n_2_11_1), .ZN(n_1023));
   AOI21_X1 i_2_11_1 (.A(n_2_60), .B1(n_952), .B2(n_2_61), .ZN(n_2_11_0));
   INV_X1 i_2_11_2 (.A(n_2_62), .ZN(n_2_11_1));
   OAI21_X1 i_2_12_0 (.A(n_2_12_0), .B1(n_952), .B2(n_2_12_1), .ZN(n_1024));
   AOI21_X1 i_2_12_1 (.A(n_2_67), .B1(n_952), .B2(n_542), .ZN(n_2_12_0));
   INV_X1 i_2_12_2 (.A(n_543), .ZN(n_2_12_1));
   OAI21_X1 i_2_13_0 (.A(n_2_13_0), .B1(n_952), .B2(n_2_13_1), .ZN(n_1025));
   AOI21_X1 i_2_13_1 (.A(n_2_68), .B1(n_952), .B2(n_537), .ZN(n_2_13_0));
   INV_X1 i_2_13_2 (.A(n_538), .ZN(n_2_13_1));
   OAI21_X1 i_2_14_0 (.A(n_2_14_0), .B1(n_952), .B2(n_2_14_1), .ZN(n_1026));
   AOI21_X1 i_2_14_1 (.A(n_2_69), .B1(n_952), .B2(n_532), .ZN(n_2_14_0));
   INV_X1 i_2_14_2 (.A(n_533), .ZN(n_2_14_1));
   OAI21_X1 i_2_15_0 (.A(n_2_15_0), .B1(n_952), .B2(n_2_15_1), .ZN(n_1027));
   AOI21_X1 i_2_15_1 (.A(n_2_70), .B1(n_952), .B2(n_527), .ZN(n_2_15_0));
   INV_X1 i_2_15_2 (.A(n_528), .ZN(n_2_15_1));
   OAI21_X1 i_2_16_0 (.A(n_2_16_0), .B1(n_952), .B2(n_2_16_1), .ZN(n_1028));
   AOI21_X1 i_2_16_1 (.A(n_2_71), .B1(n_952), .B2(n_522), .ZN(n_2_16_0));
   INV_X1 i_2_16_2 (.A(n_523), .ZN(n_2_16_1));
   OAI21_X1 i_2_17_0 (.A(n_2_17_0), .B1(n_952), .B2(n_2_17_1), .ZN(n_1029));
   AOI21_X1 i_2_17_1 (.A(n_2_75), .B1(n_952), .B2(n_502), .ZN(n_2_17_0));
   INV_X1 i_2_17_2 (.A(n_503), .ZN(n_2_17_1));
   OAI21_X1 i_2_18_0 (.A(n_2_18_0), .B1(n_952), .B2(n_2_18_1), .ZN(n_1030));
   AOI21_X1 i_2_18_1 (.A(n_2_76), .B1(n_952), .B2(n_497), .ZN(n_2_18_0));
   INV_X1 i_2_18_2 (.A(n_498), .ZN(n_2_18_1));
   OAI21_X1 i_2_19_0 (.A(n_2_19_0), .B1(n_952), .B2(n_2_19_1), .ZN(n_1031));
   AOI21_X1 i_2_19_1 (.A(n_2_77), .B1(n_952), .B2(n_492), .ZN(n_2_19_0));
   INV_X1 i_2_19_2 (.A(n_493), .ZN(n_2_19_1));
   OAI21_X1 i_2_20_0 (.A(n_2_20_0), .B1(n_952), .B2(n_2_20_1), .ZN(n_1032));
   AOI21_X1 i_2_20_1 (.A(n_2_78), .B1(n_952), .B2(n_487), .ZN(n_2_20_0));
   INV_X1 i_2_20_2 (.A(n_488), .ZN(n_2_20_1));
   OAI21_X1 i_2_21_0 (.A(n_2_21_0), .B1(n_952), .B2(n_2_21_1), .ZN(n_1033));
   AOI21_X1 i_2_21_1 (.A(n_2_80), .B1(n_952), .B2(n_2_81), .ZN(n_2_21_0));
   INV_X1 i_2_21_2 (.A(n_2_82), .ZN(n_2_21_1));
   OAI21_X1 i_2_22_0 (.A(n_2_22_0), .B1(n_952), .B2(n_2_22_1), .ZN(n_1034));
   AOI21_X1 i_2_22_1 (.A(n_2_83), .B1(n_952), .B2(n_2_84), .ZN(n_2_22_0));
   INV_X1 i_2_22_2 (.A(n_2_85), .ZN(n_2_22_1));
   OAI21_X1 i_2_23_0 (.A(n_2_23_0), .B1(n_952), .B2(n_2_23_1), .ZN(n_1035));
   AOI21_X1 i_2_23_1 (.A(n_2_86), .B1(n_952), .B2(n_2_87), .ZN(n_2_23_0));
   INV_X1 i_2_23_2 (.A(n_2_88), .ZN(n_2_23_1));
   OAI21_X1 i_2_24_0 (.A(n_2_24_0), .B1(n_952), .B2(n_2_24_1), .ZN(n_1036));
   AOI21_X1 i_2_24_1 (.A(n_2_89), .B1(n_952), .B2(n_1203), .ZN(n_2_24_0));
   INV_X1 i_2_24_2 (.A(n_465), .ZN(n_2_24_1));
   OAI21_X1 i_2_25_0 (.A(n_2_25_0), .B1(n_952), .B2(n_2_25_1), .ZN(n_1037));
   AOI21_X1 i_2_25_1 (.A(n_2_90), .B1(n_952), .B2(n_460), .ZN(n_2_25_0));
   INV_X1 i_2_25_2 (.A(n_461), .ZN(n_2_25_1));
   OAI21_X1 i_2_26_0 (.A(n_2_26_0), .B1(n_952), .B2(n_2_26_1), .ZN(n_1038));
   AOI21_X1 i_2_26_1 (.A(n_2_91), .B1(n_952), .B2(n_455), .ZN(n_2_26_0));
   INV_X1 i_2_26_2 (.A(n_456), .ZN(n_2_26_1));
   OAI21_X1 i_2_27_0 (.A(n_2_27_0), .B1(n_952), .B2(n_2_27_1), .ZN(n_1039));
   AOI21_X1 i_2_27_1 (.A(n_2_93), .B1(n_952), .B2(n_445), .ZN(n_2_27_0));
   INV_X1 i_2_27_2 (.A(n_446), .ZN(n_2_27_1));
   OAI21_X1 i_2_28_0 (.A(n_2_28_0), .B1(n_952), .B2(n_2_28_1), .ZN(n_1040));
   AOI21_X1 i_2_28_1 (.A(n_2_94), .B1(n_952), .B2(n_2_95), .ZN(n_2_28_0));
   INV_X1 i_2_28_2 (.A(n_440), .ZN(n_2_28_1));
   OAI21_X1 i_2_29_0 (.A(n_2_29_0), .B1(n_952), .B2(n_2_29_1), .ZN(n_1041));
   AOI21_X1 i_2_29_1 (.A(n_2_97), .B1(n_952), .B2(n_2_98), .ZN(n_2_29_0));
   INV_X1 i_2_29_2 (.A(n_2_99), .ZN(n_2_29_1));
   OAI21_X1 i_2_30_0 (.A(n_2_30_0), .B1(n_952), .B2(n_2_30_1), .ZN(n_1042));
   AOI21_X1 i_2_30_1 (.A(n_2_100), .B1(n_952), .B2(n_426), .ZN(n_2_30_0));
   INV_X1 i_2_30_2 (.A(n_427), .ZN(n_2_30_1));
   OAI21_X1 i_2_31_0 (.A(n_2_31_0), .B1(n_952), .B2(n_2_31_1), .ZN(n_1043));
   AOI21_X1 i_2_31_1 (.A(n_2_102), .B1(n_952), .B2(n_416), .ZN(n_2_31_0));
   INV_X1 i_2_31_2 (.A(n_417), .ZN(n_2_31_1));
   OAI21_X1 i_2_32_0 (.A(n_2_32_0), .B1(n_952), .B2(n_2_32_1), .ZN(n_1044));
   AOI21_X1 i_2_32_1 (.A(n_2_104), .B1(n_952), .B2(n_406), .ZN(n_2_32_0));
   INV_X1 i_2_32_2 (.A(n_407), .ZN(n_2_32_1));
   OAI21_X1 i_2_33_0 (.A(n_2_33_0), .B1(n_952), .B2(n_2_33_1), .ZN(n_1045));
   AOI21_X1 i_2_33_1 (.A(n_2_112), .B1(n_952), .B2(n_378), .ZN(n_2_33_0));
   INV_X1 i_2_33_2 (.A(n_379), .ZN(n_2_33_1));
   OAI21_X1 i_2_34_0 (.A(n_2_34_0), .B1(n_952), .B2(n_2_34_1), .ZN(n_1046));
   AOI21_X1 i_2_34_1 (.A(n_2_113), .B1(n_952), .B2(n_2_114), .ZN(n_2_34_0));
   INV_X1 i_2_34_2 (.A(n_2_115), .ZN(n_2_34_1));
   OAI21_X1 i_2_35_0 (.A(n_2_35_0), .B1(n_952), .B2(n_2_35_1), .ZN(n_1047));
   AOI21_X1 i_2_35_1 (.A(n_2_116), .B1(n_952), .B2(n_2_117), .ZN(n_2_35_0));
   INV_X1 i_2_35_2 (.A(n_2_118), .ZN(n_2_35_1));
   OAI21_X1 i_2_36_0 (.A(n_2_36_0), .B1(n_952), .B2(n_2_36_1), .ZN(n_1048));
   AOI21_X1 i_2_36_1 (.A(n_2_119), .B1(n_952), .B2(n_367), .ZN(n_2_36_0));
   INV_X1 i_2_36_2 (.A(n_368), .ZN(n_2_36_1));
   OAI21_X1 i_2_37_0 (.A(n_2_37_0), .B1(n_952), .B2(n_2_37_1), .ZN(n_1049));
   AOI21_X1 i_2_37_1 (.A(n_2_120), .B1(n_952), .B2(n_362), .ZN(n_2_37_0));
   INV_X1 i_2_37_2 (.A(n_363), .ZN(n_2_37_1));
   OAI21_X1 i_2_38_0 (.A(n_2_38_0), .B1(n_952), .B2(n_2_38_1), .ZN(n_1050));
   AOI21_X1 i_2_38_1 (.A(n_2_121), .B1(n_952), .B2(n_357), .ZN(n_2_38_0));
   INV_X1 i_2_38_2 (.A(n_358), .ZN(n_2_38_1));
   OAI21_X1 i_2_39_0 (.A(n_2_39_0), .B1(n_952), .B2(n_2_39_1), .ZN(n_1051));
   AOI21_X1 i_2_39_1 (.A(n_2_122), .B1(n_952), .B2(n_352), .ZN(n_2_39_0));
   INV_X1 i_2_39_2 (.A(n_353), .ZN(n_2_39_1));
   OAI21_X1 i_2_40_0 (.A(n_2_40_0), .B1(n_952), .B2(n_2_40_1), .ZN(n_1052));
   AOI21_X1 i_2_40_1 (.A(n_2_123), .B1(n_952), .B2(n_2_124), .ZN(n_2_40_0));
   INV_X1 i_2_40_2 (.A(n_2_125), .ZN(n_2_40_1));
   OAI21_X1 i_2_41_0 (.A(n_2_41_0), .B1(n_952), .B2(n_2_41_1), .ZN(n_1053));
   AOI21_X1 i_2_41_1 (.A(n_2_126), .B1(n_952), .B2(n_344), .ZN(n_2_41_0));
   INV_X1 i_2_41_2 (.A(n_345), .ZN(n_2_41_1));
   OAI21_X1 i_2_42_0 (.A(n_2_42_0), .B1(n_952), .B2(n_2_42_1), .ZN(n_1054));
   AOI21_X1 i_2_42_1 (.A(n_2_127), .B1(n_952), .B2(n_339), .ZN(n_2_42_0));
   INV_X1 i_2_42_2 (.A(n_340), .ZN(n_2_42_1));
   OAI21_X1 i_2_43_0 (.A(n_2_43_0), .B1(n_952), .B2(n_2_43_1), .ZN(n_1055));
   AOI21_X1 i_2_43_1 (.A(n_2_128), .B1(n_952), .B2(n_334), .ZN(n_2_43_0));
   INV_X1 i_2_43_2 (.A(n_335), .ZN(n_2_43_1));
   OAI21_X1 i_2_44_0 (.A(n_2_44_0), .B1(n_952), .B2(n_2_44_1), .ZN(n_1056));
   AOI21_X1 i_2_44_1 (.A(n_2_129), .B1(n_952), .B2(n_2_130), .ZN(n_2_44_0));
   INV_X1 i_2_44_2 (.A(n_2_131), .ZN(n_2_44_1));
   OAI21_X1 i_2_45_0 (.A(n_2_45_0), .B1(n_952), .B2(n_2_45_1), .ZN(n_1057));
   AOI21_X1 i_2_45_1 (.A(n_2_138), .B1(n_952), .B2(n_320), .ZN(n_2_45_0));
   INV_X1 i_2_45_2 (.A(n_321), .ZN(n_2_45_1));
   OAI21_X1 i_2_46_0 (.A(n_2_46_0), .B1(n_952), .B2(n_2_46_1), .ZN(n_1058));
   AOI21_X1 i_2_46_1 (.A(n_2_142), .B1(n_952), .B2(n_312), .ZN(n_2_46_0));
   INV_X1 i_2_46_2 (.A(n_313), .ZN(n_2_46_1));
   OAI21_X1 i_2_47_0 (.A(n_2_47_0), .B1(n_952), .B2(n_2_47_1), .ZN(n_1059));
   AOI21_X1 i_2_47_1 (.A(n_2_150), .B1(n_952), .B2(n_2_151), .ZN(n_2_47_0));
   INV_X1 i_2_47_2 (.A(n_2_152), .ZN(n_2_47_1));
   OAI21_X1 i_2_48_0 (.A(n_2_48_0), .B1(n_952), .B2(n_2_48_1), .ZN(n_1060));
   AOI21_X1 i_2_48_1 (.A(n_2_153), .B1(n_952), .B2(n_2_154), .ZN(n_2_48_0));
   INV_X1 i_2_48_2 (.A(n_2_155), .ZN(n_2_48_1));
   OAI21_X1 i_2_49_0 (.A(n_2_49_0), .B1(n_952), .B2(n_2_49_1), .ZN(n_1061));
   AOI21_X1 i_2_49_1 (.A(n_2_156), .B1(n_952), .B2(n_290), .ZN(n_2_49_0));
   INV_X1 i_2_49_2 (.A(n_291), .ZN(n_2_49_1));
   OAI21_X1 i_2_50_0 (.A(n_2_50_0), .B1(n_952), .B2(n_2_50_1), .ZN(n_1062));
   AOI21_X1 i_2_50_1 (.A(n_2_157), .B1(n_952), .B2(n_2_158), .ZN(n_2_50_0));
   INV_X1 i_2_50_2 (.A(n_2_159), .ZN(n_2_50_1));
   OAI21_X1 i_2_51_0 (.A(n_2_51_0), .B1(n_952), .B2(n_2_51_1), .ZN(n_1063));
   AOI21_X1 i_2_51_1 (.A(n_2_160), .B1(n_952), .B2(n_282), .ZN(n_2_51_0));
   INV_X1 i_2_51_2 (.A(n_283), .ZN(n_2_51_1));
   OAI21_X1 i_2_52_0 (.A(n_2_52_0), .B1(n_952), .B2(n_2_52_1), .ZN(n_1064));
   AOI21_X1 i_2_52_1 (.A(n_2_161), .B1(n_952), .B2(n_1204), .ZN(n_2_52_0));
   INV_X1 i_2_52_2 (.A(n_1205), .ZN(n_2_52_1));
   OAI21_X1 i_2_53_0 (.A(n_2_53_0), .B1(n_952), .B2(n_2_53_1), .ZN(n_1065));
   AOI21_X1 i_2_53_1 (.A(n_2_162), .B1(n_952), .B2(n_271), .ZN(n_2_53_0));
   INV_X1 i_2_53_2 (.A(n_272), .ZN(n_2_53_1));
   OAI21_X1 i_2_54_0 (.A(n_2_54_0), .B1(n_952), .B2(n_2_54_1), .ZN(n_1066));
   AOI21_X1 i_2_54_1 (.A(n_2_163), .B1(n_952), .B2(n_266), .ZN(n_2_54_0));
   INV_X1 i_2_54_2 (.A(n_267), .ZN(n_2_54_1));
   OAI21_X1 i_2_55_0 (.A(n_2_55_0), .B1(n_952), .B2(n_2_55_1), .ZN(n_1067));
   AOI21_X1 i_2_55_1 (.A(n_2_167), .B1(n_952), .B2(n_255), .ZN(n_2_55_0));
   INV_X1 i_2_55_2 (.A(n_256), .ZN(n_2_55_1));
   OAI21_X1 i_2_56_0 (.A(n_2_56_0), .B1(n_952), .B2(n_2_56_1), .ZN(n_1068));
   AOI21_X1 i_2_56_1 (.A(n_2_168), .B1(n_952), .B2(n_2_169), .ZN(n_2_56_0));
   INV_X1 i_2_56_2 (.A(n_2_170), .ZN(n_2_56_1));
   OAI21_X1 i_2_57_0 (.A(n_2_57_0), .B1(n_952), .B2(n_2_57_1), .ZN(n_1069));
   AOI21_X1 i_2_57_1 (.A(n_2_172), .B1(n_952), .B2(n_242), .ZN(n_2_57_0));
   INV_X1 i_2_57_2 (.A(n_243), .ZN(n_2_57_1));
   OAI21_X1 i_2_58_0 (.A(n_2_58_0), .B1(n_952), .B2(n_2_58_1), .ZN(n_1070));
   AOI21_X1 i_2_58_1 (.A(n_2_173), .B1(n_952), .B2(n_237), .ZN(n_2_58_0));
   INV_X1 i_2_58_2 (.A(n_238), .ZN(n_2_58_1));
   OAI21_X1 i_2_59_0 (.A(n_2_59_0), .B1(n_952), .B2(n_2_59_1), .ZN(n_1071));
   AOI21_X1 i_2_59_1 (.A(n_2_174), .B1(n_952), .B2(n_232), .ZN(n_2_59_0));
   INV_X1 i_2_59_2 (.A(n_233), .ZN(n_2_59_1));
   OAI21_X1 i_2_60_0 (.A(n_2_60_0), .B1(n_952), .B2(n_2_60_1), .ZN(n_1072));
   AOI21_X1 i_2_60_1 (.A(n_2_180), .B1(n_952), .B2(n_2_181), .ZN(n_2_60_0));
   INV_X1 i_2_60_2 (.A(n_2_182), .ZN(n_2_60_1));
   OAI21_X1 i_2_61_0 (.A(n_2_61_0), .B1(n_952), .B2(n_2_61_1), .ZN(n_1073));
   AOI21_X1 i_2_61_1 (.A(n_2_184), .B1(n_952), .B2(n_1206), .ZN(n_2_61_0));
   INV_X1 i_2_61_2 (.A(n_1207), .ZN(n_2_61_1));
   OAI21_X1 i_2_62_0 (.A(n_2_62_0), .B1(n_952), .B2(n_2_62_1), .ZN(n_1074));
   AOI21_X1 i_2_62_1 (.A(n_2_185), .B1(n_952), .B2(n_2_186), .ZN(n_2_62_0));
   INV_X1 i_2_62_2 (.A(n_2_187), .ZN(n_2_62_1));
   OAI21_X1 i_2_63_0 (.A(n_2_63_0), .B1(n_952), .B2(n_2_63_1), .ZN(n_1075));
   AOI21_X1 i_2_63_1 (.A(n_2_188), .B1(n_952), .B2(n_2_189), .ZN(n_2_63_0));
   INV_X1 i_2_63_2 (.A(n_2_190), .ZN(n_2_63_1));
   OAI21_X1 i_2_64_0 (.A(n_2_64_0), .B1(n_952), .B2(n_2_64_1), .ZN(n_1076));
   AOI21_X1 i_2_64_1 (.A(n_2_194), .B1(n_952), .B2(n_179), .ZN(n_2_64_0));
   INV_X1 i_2_64_2 (.A(n_180), .ZN(n_2_64_1));
   OAI21_X1 i_2_65_0 (.A(n_2_65_0), .B1(n_952), .B2(n_2_65_1), .ZN(n_1077));
   AOI21_X1 i_2_65_1 (.A(n_2_196), .B1(n_952), .B2(n_169), .ZN(n_2_65_0));
   INV_X1 i_2_65_2 (.A(n_170), .ZN(n_2_65_1));
   OAI21_X1 i_2_66_0 (.A(n_2_66_0), .B1(n_952), .B2(n_2_66_1), .ZN(n_1078));
   AOI21_X1 i_2_66_1 (.A(n_2_197), .B1(n_952), .B2(n_164), .ZN(n_2_66_0));
   INV_X1 i_2_66_2 (.A(n_165), .ZN(n_2_66_1));
   OAI21_X1 i_2_67_0 (.A(n_2_67_0), .B1(n_952), .B2(n_2_67_1), .ZN(n_1079));
   AOI21_X1 i_2_67_1 (.A(n_2_198), .B1(n_952), .B2(n_2_199), .ZN(n_2_67_0));
   INV_X1 i_2_67_2 (.A(n_2_200), .ZN(n_2_67_1));
   OAI21_X1 i_2_68_0 (.A(n_2_68_0), .B1(n_952), .B2(n_2_68_1), .ZN(n_1080));
   AOI21_X1 i_2_68_1 (.A(n_2_201), .B1(n_952), .B2(n_153), .ZN(n_2_68_0));
   INV_X1 i_2_68_2 (.A(n_154), .ZN(n_2_68_1));
   OAI21_X1 i_2_69_0 (.A(n_2_69_0), .B1(n_952), .B2(n_2_69_1), .ZN(n_1081));
   AOI21_X1 i_2_69_1 (.A(n_2_202), .B1(n_952), .B2(n_1208), .ZN(n_2_69_0));
   INV_X1 i_2_69_2 (.A(n_1209), .ZN(n_2_69_1));
   OAI21_X1 i_2_70_0 (.A(n_2_70_0), .B1(n_952), .B2(n_2_70_1), .ZN(n_1082));
   AOI21_X1 i_2_70_1 (.A(n_2_203), .B1(n_952), .B2(n_1210), .ZN(n_2_70_0));
   INV_X1 i_2_70_2 (.A(n_1211), .ZN(n_2_70_1));
   OAI21_X1 i_2_71_0 (.A(n_2_71_0), .B1(n_952), .B2(n_2_71_1), .ZN(n_1083));
   AOI21_X1 i_2_71_1 (.A(n_2_205), .B1(n_952), .B2(n_138), .ZN(n_2_71_0));
   INV_X1 i_2_71_2 (.A(n_2_206), .ZN(n_2_71_1));
   OAI21_X1 i_2_72_0 (.A(n_2_72_0), .B1(n_2_72_3), .B2(n_2_72_1), .ZN(n_1084));
   NAND2_X1 i_2_72_1 (.A1(n_2_225), .A2(n_2_72_1), .ZN(n_2_72_0));
   OAI22_X1 i_2_72_2 (.A1(n_952), .A2(n_2_182), .B1(n_2_72_2), .B2(n_2_181), 
      .ZN(n_2_72_1));
   INV_X1 i_2_72_3 (.A(n_952), .ZN(n_2_72_2));
   INV_X1 i_2_72_4 (.A(in_data[4]), .ZN(n_2_72_3));
   OAI21_X1 i_2_73_0 (.A(n_2_73_0), .B1(n_2_73_3), .B2(n_2_73_1), .ZN(n_1085));
   NAND2_X1 i_2_73_1 (.A1(n_2_226), .A2(n_2_73_1), .ZN(n_2_73_0));
   OAI22_X1 i_2_73_2 (.A1(n_952), .A2(n_2_187), .B1(n_2_73_2), .B2(n_2_186), 
      .ZN(n_2_73_1));
   INV_X1 i_2_73_3 (.A(n_952), .ZN(n_2_73_2));
   INV_X1 i_2_73_4 (.A(in_data[4]), .ZN(n_2_73_3));
   OAI21_X1 i_2_74_0 (.A(n_2_74_0), .B1(n_2_74_3), .B2(n_2_74_1), .ZN(n_1086));
   NAND2_X1 i_2_74_1 (.A1(n_2_227), .A2(n_2_74_1), .ZN(n_2_74_0));
   OAI22_X1 i_2_74_2 (.A1(n_952), .A2(n_2_190), .B1(n_2_74_2), .B2(n_2_189), 
      .ZN(n_2_74_1));
   INV_X1 i_2_74_3 (.A(n_952), .ZN(n_2_74_2));
   INV_X1 i_2_74_4 (.A(in_data[4]), .ZN(n_2_74_3));
   OAI21_X1 i_2_75_0 (.A(n_2_75_0), .B1(n_2_75_3), .B2(n_2_75_1), .ZN(n_1087));
   NAND2_X1 i_2_75_1 (.A1(n_2_228), .A2(n_2_75_1), .ZN(n_2_75_0));
   OAI22_X1 i_2_75_2 (.A1(n_952), .A2(n_2_200), .B1(n_2_75_2), .B2(n_2_199), 
      .ZN(n_2_75_1));
   INV_X1 i_2_75_3 (.A(n_952), .ZN(n_2_75_2));
   INV_X1 i_2_75_4 (.A(in_data[4]), .ZN(n_2_75_3));
   OAI21_X1 i_2_76_0 (.A(n_2_76_0), .B1(n_2_339), .B2(n_2_76_1), .ZN(n_2_1));
   AOI21_X1 i_2_76_1 (.A(n_663), .B1(n_2_339), .B2(n_661), .ZN(n_2_76_0));
   INV_X1 i_2_76_2 (.A(n_662), .ZN(n_2_76_1));
   OAI21_X1 i_2_77_0 (.A(n_2_77_0), .B1(n_2_339), .B2(n_2_77_1), .ZN(n_2_4));
   AOI21_X1 i_2_77_1 (.A(n_658), .B1(n_2_339), .B2(n_656), .ZN(n_2_77_0));
   INV_X1 i_2_77_2 (.A(n_657), .ZN(n_2_77_1));
   OAI21_X1 i_2_78_0 (.A(n_2_78_0), .B1(n_2_339), .B2(n_2_78_1), .ZN(n_2_5));
   AOI21_X1 i_2_78_1 (.A(n_655), .B1(n_2_339), .B2(n_653), .ZN(n_2_78_0));
   INV_X1 i_2_78_2 (.A(n_654), .ZN(n_2_78_1));
   OAI21_X1 i_2_79_0 (.A(n_2_79_0), .B1(n_2_339), .B2(n_2_79_1), .ZN(n_2_17));
   AOI21_X1 i_2_79_1 (.A(n_631), .B1(n_2_339), .B2(n_629), .ZN(n_2_79_0));
   INV_X1 i_2_79_2 (.A(n_630), .ZN(n_2_79_1));
   OR2_X1 i_2_80_0 (.A1(n_1016), .A2(n_2_241), .ZN(n_1088));
   OAI21_X1 i_2_81_0 (.A(n_2_81_0), .B1(n_2_339), .B2(n_2_81_1), .ZN(n_2_21));
   AOI21_X1 i_2_81_1 (.A(n_623), .B1(n_2_339), .B2(n_621), .ZN(n_2_81_0));
   INV_X1 i_2_81_2 (.A(n_622), .ZN(n_2_81_1));
   OAI21_X1 i_2_82_0 (.A(n_2_82_0), .B1(n_2_339), .B2(n_2_82_1), .ZN(n_2_22));
   AOI21_X1 i_2_82_1 (.A(n_619), .B1(n_2_339), .B2(n_617), .ZN(n_2_82_0));
   INV_X1 i_2_82_2 (.A(n_618), .ZN(n_2_82_1));
   OAI21_X1 i_2_83_0 (.A(n_2_83_0), .B1(n_2_339), .B2(n_2_83_1), .ZN(n_2_28));
   AOI21_X1 i_2_83_1 (.A(n_604), .B1(n_2_339), .B2(n_602), .ZN(n_2_83_0));
   INV_X1 i_2_83_2 (.A(n_603), .ZN(n_2_83_1));
   OAI21_X1 i_2_84_0 (.A(n_2_84_0), .B1(n_2_339), .B2(n_2_84_1), .ZN(n_2_38));
   AOI21_X1 i_2_84_1 (.A(n_587), .B1(n_2_339), .B2(n_838), .ZN(n_2_84_0));
   INV_X1 i_2_84_2 (.A(n_832), .ZN(n_2_84_1));
   OAI21_X1 i_2_85_0 (.A(n_2_85_0), .B1(n_2_339), .B2(n_2_85_1), .ZN(n_2_50));
   AOI21_X1 i_2_85_1 (.A(n_573), .B1(n_2_339), .B2(n_571), .ZN(n_2_85_0));
   INV_X1 i_2_85_2 (.A(n_572), .ZN(n_2_85_1));
   OAI21_X1 i_2_86_0 (.A(n_2_86_0), .B1(n_2_339), .B2(n_2_86_1), .ZN(n_2_53));
   AOI21_X1 i_2_86_1 (.A(n_569), .B1(n_2_339), .B2(n_567), .ZN(n_2_86_0));
   INV_X1 i_2_86_2 (.A(n_568), .ZN(n_2_86_1));
   OAI21_X1 i_2_87_0 (.A(n_2_87_0), .B1(n_2_339), .B2(n_2_87_1), .ZN(n_2_56));
   AOI21_X1 i_2_87_1 (.A(n_565), .B1(n_2_339), .B2(n_563), .ZN(n_2_87_0));
   INV_X1 i_2_87_2 (.A(n_564), .ZN(n_2_87_1));
   OAI21_X1 i_2_88_0 (.A(n_2_88_0), .B1(n_2_339), .B2(n_2_88_1), .ZN(n_2_60));
   AOI21_X1 i_2_88_1 (.A(n_557), .B1(n_2_339), .B2(n_555), .ZN(n_2_88_0));
   INV_X1 i_2_88_2 (.A(n_556), .ZN(n_2_88_1));
   OAI21_X1 i_2_89_0 (.A(n_2_89_0), .B1(n_2_339), .B2(n_2_89_1), .ZN(n_2_67));
   AOI21_X1 i_2_89_1 (.A(n_546), .B1(n_2_339), .B2(n_544), .ZN(n_2_89_0));
   INV_X1 i_2_89_2 (.A(n_545), .ZN(n_2_89_1));
   OAI21_X1 i_2_90_0 (.A(n_2_90_0), .B1(n_2_339), .B2(n_2_90_1), .ZN(n_2_68));
   AOI21_X1 i_2_90_1 (.A(n_541), .B1(n_2_339), .B2(n_539), .ZN(n_2_90_0));
   INV_X1 i_2_90_2 (.A(n_540), .ZN(n_2_90_1));
   OAI21_X1 i_2_91_0 (.A(n_2_91_0), .B1(n_2_339), .B2(n_2_91_1), .ZN(n_2_69));
   AOI21_X1 i_2_91_1 (.A(n_536), .B1(n_2_339), .B2(n_534), .ZN(n_2_91_0));
   INV_X1 i_2_91_2 (.A(n_535), .ZN(n_2_91_1));
   OAI21_X1 i_2_92_0 (.A(n_2_92_0), .B1(n_2_339), .B2(n_2_92_1), .ZN(n_2_70));
   AOI21_X1 i_2_92_1 (.A(n_531), .B1(n_2_339), .B2(n_529), .ZN(n_2_92_0));
   INV_X1 i_2_92_2 (.A(n_530), .ZN(n_2_92_1));
   OAI21_X1 i_2_93_0 (.A(n_2_93_0), .B1(n_2_339), .B2(n_2_93_1), .ZN(n_2_71));
   AOI21_X1 i_2_93_1 (.A(n_526), .B1(n_2_339), .B2(n_524), .ZN(n_2_93_0));
   INV_X1 i_2_93_2 (.A(n_525), .ZN(n_2_93_1));
   OAI21_X1 i_2_94_0 (.A(n_2_94_0), .B1(n_2_339), .B2(n_2_94_1), .ZN(n_2_75));
   AOI21_X1 i_2_94_1 (.A(n_506), .B1(n_2_339), .B2(n_504), .ZN(n_2_94_0));
   INV_X1 i_2_94_2 (.A(n_505), .ZN(n_2_94_1));
   OAI21_X1 i_2_95_0 (.A(n_2_95_0), .B1(n_2_339), .B2(n_2_95_1), .ZN(n_2_76));
   AOI21_X1 i_2_95_1 (.A(n_501), .B1(n_2_339), .B2(n_499), .ZN(n_2_95_0));
   INV_X1 i_2_95_2 (.A(n_500), .ZN(n_2_95_1));
   OAI21_X1 i_2_96_0 (.A(n_2_96_0), .B1(n_2_339), .B2(n_2_96_1), .ZN(n_2_77));
   AOI21_X1 i_2_96_1 (.A(n_496), .B1(n_2_339), .B2(n_494), .ZN(n_2_96_0));
   INV_X1 i_2_96_2 (.A(n_495), .ZN(n_2_96_1));
   OAI21_X1 i_2_97_0 (.A(n_2_97_0), .B1(n_2_339), .B2(n_2_97_1), .ZN(n_2_78));
   AOI21_X1 i_2_97_1 (.A(n_491), .B1(n_2_339), .B2(n_489), .ZN(n_2_97_0));
   INV_X1 i_2_97_2 (.A(n_490), .ZN(n_2_97_1));
   OAI21_X1 i_2_98_0 (.A(n_2_98_0), .B1(n_2_339), .B2(n_2_98_1), .ZN(n_2_80));
   AOI21_X1 i_2_98_1 (.A(n_481), .B1(n_2_339), .B2(n_479), .ZN(n_2_98_0));
   INV_X1 i_2_98_2 (.A(n_480), .ZN(n_2_98_1));
   OAI21_X1 i_2_99_0 (.A(n_2_99_0), .B1(n_2_339), .B2(n_2_99_1), .ZN(n_2_83));
   AOI21_X1 i_2_99_1 (.A(n_477), .B1(n_2_339), .B2(n_475), .ZN(n_2_99_0));
   INV_X1 i_2_99_2 (.A(n_476), .ZN(n_2_99_1));
   OAI21_X1 i_2_100_0 (.A(n_2_100_0), .B1(n_2_339), .B2(n_2_100_1), .ZN(n_2_86));
   AOI21_X1 i_2_100_1 (.A(n_473), .B1(n_2_339), .B2(n_471), .ZN(n_2_100_0));
   INV_X1 i_2_100_2 (.A(n_472), .ZN(n_2_100_1));
   OAI21_X1 i_2_101_0 (.A(n_2_101_0), .B1(n_2_339), .B2(n_2_101_1), .ZN(n_2_89));
   AOI21_X1 i_2_101_1 (.A(n_469), .B1(n_2_339), .B2(n_467), .ZN(n_2_101_0));
   INV_X1 i_2_101_2 (.A(n_468), .ZN(n_2_101_1));
   OAI21_X1 i_2_102_0 (.A(n_2_102_0), .B1(n_2_339), .B2(n_2_102_1), .ZN(n_2_90));
   AOI21_X1 i_2_102_1 (.A(n_464), .B1(n_2_339), .B2(n_462), .ZN(n_2_102_0));
   INV_X1 i_2_102_2 (.A(n_463), .ZN(n_2_102_1));
   OAI21_X1 i_2_103_0 (.A(n_2_103_0), .B1(n_2_339), .B2(n_2_103_1), .ZN(n_2_91));
   AOI21_X1 i_2_103_1 (.A(n_459), .B1(n_2_339), .B2(n_457), .ZN(n_2_103_0));
   INV_X1 i_2_103_2 (.A(n_458), .ZN(n_2_103_1));
   OAI21_X1 i_2_104_0 (.A(n_2_104_0), .B1(n_2_339), .B2(n_2_104_1), .ZN(n_2_93));
   AOI21_X1 i_2_104_1 (.A(n_449), .B1(n_2_339), .B2(n_447), .ZN(n_2_104_0));
   INV_X1 i_2_104_2 (.A(n_448), .ZN(n_2_104_1));
   OAI21_X1 i_2_105_0 (.A(n_2_105_0), .B1(n_2_339), .B2(n_2_105_1), .ZN(n_2_94));
   AOI21_X1 i_2_105_1 (.A(n_444), .B1(n_2_339), .B2(n_442), .ZN(n_2_105_0));
   INV_X1 i_2_105_2 (.A(n_443), .ZN(n_2_105_1));
   OAI21_X1 i_2_106_0 (.A(n_2_106_0), .B1(n_2_339), .B2(n_2_106_1), .ZN(n_2_97));
   AOI21_X1 i_2_106_1 (.A(n_434), .B1(n_2_339), .B2(n_432), .ZN(n_2_106_0));
   INV_X1 i_2_106_2 (.A(n_433), .ZN(n_2_106_1));
   OAI21_X1 i_2_107_0 (.A(n_2_107_0), .B1(n_2_339), .B2(n_2_107_1), .ZN(n_2_100));
   AOI21_X1 i_2_107_1 (.A(n_430), .B1(n_2_339), .B2(n_428), .ZN(n_2_107_0));
   INV_X1 i_2_107_2 (.A(n_429), .ZN(n_2_107_1));
   OAI21_X1 i_2_108_0 (.A(n_2_108_0), .B1(n_2_339), .B2(n_2_108_1), .ZN(n_2_102));
   AOI21_X1 i_2_108_1 (.A(n_420), .B1(n_2_339), .B2(n_418), .ZN(n_2_108_0));
   INV_X1 i_2_108_2 (.A(n_419), .ZN(n_2_108_1));
   OAI21_X1 i_2_109_0 (.A(n_2_109_0), .B1(n_2_339), .B2(n_2_109_1), .ZN(n_2_104));
   AOI21_X1 i_2_109_1 (.A(n_410), .B1(n_2_339), .B2(n_408), .ZN(n_2_109_0));
   INV_X1 i_2_109_2 (.A(n_409), .ZN(n_2_109_1));
   OAI21_X1 i_2_110_0 (.A(n_2_110_0), .B1(n_2_339), .B2(n_2_110_1), .ZN(n_2_112));
   AOI21_X1 i_2_110_1 (.A(n_382), .B1(n_2_339), .B2(n_380), .ZN(n_2_110_0));
   INV_X1 i_2_110_2 (.A(n_381), .ZN(n_2_110_1));
   OAI21_X1 i_2_111_0 (.A(n_2_111_0), .B1(n_2_339), .B2(n_2_111_1), .ZN(n_2_113));
   AOI21_X1 i_2_111_1 (.A(n_377), .B1(n_2_339), .B2(n_375), .ZN(n_2_111_0));
   INV_X1 i_2_111_2 (.A(n_376), .ZN(n_2_111_1));
   OAI21_X1 i_2_112_0 (.A(n_2_112_0), .B1(n_2_339), .B2(n_2_112_1), .ZN(n_2_116));
   AOI21_X1 i_2_112_1 (.A(n_374), .B1(n_2_339), .B2(n_372), .ZN(n_2_112_0));
   INV_X1 i_2_112_2 (.A(n_373), .ZN(n_2_112_1));
   OAI21_X1 i_2_113_0 (.A(n_2_113_0), .B1(n_2_339), .B2(n_2_113_1), .ZN(n_2_119));
   AOI21_X1 i_2_113_1 (.A(n_371), .B1(n_2_339), .B2(n_369), .ZN(n_2_113_0));
   INV_X1 i_2_113_2 (.A(n_370), .ZN(n_2_113_1));
   OAI21_X1 i_2_114_0 (.A(n_2_114_0), .B1(n_2_339), .B2(n_2_114_1), .ZN(n_2_120));
   AOI21_X1 i_2_114_1 (.A(n_366), .B1(n_2_339), .B2(n_364), .ZN(n_2_114_0));
   INV_X1 i_2_114_2 (.A(n_365), .ZN(n_2_114_1));
   OAI21_X1 i_2_115_0 (.A(n_2_115_0), .B1(n_2_339), .B2(n_2_115_1), .ZN(n_2_121));
   AOI21_X1 i_2_115_1 (.A(n_361), .B1(n_2_339), .B2(n_359), .ZN(n_2_115_0));
   INV_X1 i_2_115_2 (.A(n_360), .ZN(n_2_115_1));
   OAI21_X1 i_2_116_0 (.A(n_2_116_0), .B1(n_2_339), .B2(n_2_116_1), .ZN(n_2_122));
   AOI21_X1 i_2_116_1 (.A(n_356), .B1(n_2_339), .B2(n_354), .ZN(n_2_116_0));
   INV_X1 i_2_116_2 (.A(n_355), .ZN(n_2_116_1));
   OAI21_X1 i_2_117_0 (.A(n_2_117_0), .B1(n_2_339), .B2(n_2_117_1), .ZN(n_2_123));
   AOI21_X1 i_2_117_1 (.A(n_351), .B1(n_2_339), .B2(n_349), .ZN(n_2_117_0));
   INV_X1 i_2_117_2 (.A(n_350), .ZN(n_2_117_1));
   OAI21_X1 i_2_118_0 (.A(n_2_118_0), .B1(n_2_339), .B2(n_2_118_1), .ZN(n_2_126));
   AOI21_X1 i_2_118_1 (.A(n_348), .B1(n_2_339), .B2(n_346), .ZN(n_2_118_0));
   INV_X1 i_2_118_2 (.A(n_347), .ZN(n_2_118_1));
   OAI21_X1 i_2_119_0 (.A(n_2_119_0), .B1(n_2_339), .B2(n_2_119_1), .ZN(n_2_127));
   AOI21_X1 i_2_119_1 (.A(n_343), .B1(n_2_339), .B2(n_341), .ZN(n_2_119_0));
   INV_X1 i_2_119_2 (.A(n_342), .ZN(n_2_119_1));
   OAI21_X1 i_2_120_0 (.A(n_2_120_0), .B1(n_2_339), .B2(n_2_120_1), .ZN(n_2_128));
   AOI21_X1 i_2_120_1 (.A(n_338), .B1(n_2_339), .B2(n_336), .ZN(n_2_120_0));
   INV_X1 i_2_120_2 (.A(n_337), .ZN(n_2_120_1));
   OAI21_X1 i_2_121_0 (.A(n_2_121_0), .B1(n_2_339), .B2(n_2_121_1), .ZN(n_2_129));
   AOI21_X1 i_2_121_1 (.A(n_333), .B1(n_2_339), .B2(n_331), .ZN(n_2_121_0));
   INV_X1 i_2_121_2 (.A(n_332), .ZN(n_2_121_1));
   OAI21_X1 i_2_122_0 (.A(n_2_122_0), .B1(n_2_339), .B2(n_2_122_1), .ZN(n_2_138));
   AOI21_X1 i_2_122_1 (.A(n_324), .B1(n_2_339), .B2(n_322), .ZN(n_2_122_0));
   INV_X1 i_2_122_2 (.A(n_323), .ZN(n_2_122_1));
   OAI21_X1 i_2_123_0 (.A(n_2_123_0), .B1(n_2_339), .B2(n_2_123_1), .ZN(n_2_142));
   AOI21_X1 i_2_123_1 (.A(n_316), .B1(n_2_339), .B2(n_314), .ZN(n_2_123_0));
   INV_X1 i_2_123_2 (.A(n_315), .ZN(n_2_123_1));
   OAI21_X1 i_2_124_0 (.A(n_2_124_0), .B1(n_2_339), .B2(n_2_124_1), .ZN(n_2_150));
   AOI21_X1 i_2_124_1 (.A(n_300), .B1(n_2_339), .B2(n_298), .ZN(n_2_124_0));
   INV_X1 i_2_124_2 (.A(n_299), .ZN(n_2_124_1));
   OAI21_X1 i_2_125_0 (.A(n_2_125_0), .B1(n_2_339), .B2(n_2_125_1), .ZN(n_2_153));
   AOI21_X1 i_2_125_1 (.A(n_297), .B1(n_2_339), .B2(n_295), .ZN(n_2_125_0));
   INV_X1 i_2_125_2 (.A(n_296), .ZN(n_2_125_1));
   OAI21_X1 i_2_126_0 (.A(n_2_126_0), .B1(n_2_339), .B2(n_2_126_1), .ZN(n_2_156));
   AOI21_X1 i_2_126_1 (.A(n_294), .B1(n_2_339), .B2(n_292), .ZN(n_2_126_0));
   INV_X1 i_2_126_2 (.A(n_293), .ZN(n_2_126_1));
   OAI21_X1 i_2_127_0 (.A(n_2_127_0), .B1(n_2_339), .B2(n_2_127_1), .ZN(n_2_157));
   AOI21_X1 i_2_127_1 (.A(n_289), .B1(n_2_339), .B2(n_287), .ZN(n_2_127_0));
   INV_X1 i_2_127_2 (.A(n_288), .ZN(n_2_127_1));
   OAI21_X1 i_2_128_0 (.A(n_2_128_0), .B1(n_2_339), .B2(n_2_128_1), .ZN(n_2_160));
   AOI21_X1 i_2_128_1 (.A(n_286), .B1(n_2_339), .B2(n_284), .ZN(n_2_128_0));
   INV_X1 i_2_128_2 (.A(n_285), .ZN(n_2_128_1));
   OAI21_X1 i_2_129_0 (.A(n_2_129_0), .B1(n_2_339), .B2(n_2_129_1), .ZN(n_2_161));
   AOI21_X1 i_2_129_1 (.A(n_281), .B1(n_2_339), .B2(n_279), .ZN(n_2_129_0));
   INV_X1 i_2_129_2 (.A(n_280), .ZN(n_2_129_1));
   OAI21_X1 i_2_130_0 (.A(n_2_130_0), .B1(n_2_339), .B2(n_2_130_1), .ZN(n_2_162));
   AOI21_X1 i_2_130_1 (.A(n_275), .B1(n_2_339), .B2(n_273), .ZN(n_2_130_0));
   INV_X1 i_2_130_2 (.A(n_274), .ZN(n_2_130_1));
   OAI21_X1 i_2_131_0 (.A(n_2_131_0), .B1(n_2_339), .B2(n_2_131_1), .ZN(n_2_163));
   AOI21_X1 i_2_131_1 (.A(n_270), .B1(n_2_339), .B2(n_268), .ZN(n_2_131_0));
   INV_X1 i_2_131_2 (.A(n_269), .ZN(n_2_131_1));
   OAI21_X1 i_2_132_0 (.A(n_2_132_0), .B1(n_2_339), .B2(n_2_132_1), .ZN(n_2_167));
   AOI21_X1 i_2_132_1 (.A(n_259), .B1(n_2_339), .B2(n_257), .ZN(n_2_132_0));
   INV_X1 i_2_132_2 (.A(n_258), .ZN(n_2_132_1));
   OAI21_X1 i_2_133_0 (.A(n_2_133_0), .B1(n_2_339), .B2(n_2_133_1), .ZN(n_2_168));
   AOI21_X1 i_2_133_1 (.A(n_254), .B1(n_2_339), .B2(n_252), .ZN(n_2_133_0));
   INV_X1 i_2_133_2 (.A(n_253), .ZN(n_2_133_1));
   OAI21_X1 i_2_134_0 (.A(n_2_134_0), .B1(n_2_339), .B2(n_2_134_1), .ZN(n_2_172));
   AOI21_X1 i_2_134_1 (.A(n_246), .B1(n_2_339), .B2(n_244), .ZN(n_2_134_0));
   INV_X1 i_2_134_2 (.A(n_245), .ZN(n_2_134_1));
   OAI21_X1 i_2_135_0 (.A(n_2_135_0), .B1(n_2_339), .B2(n_2_135_1), .ZN(n_2_173));
   AOI21_X1 i_2_135_1 (.A(n_241), .B1(n_2_339), .B2(n_239), .ZN(n_2_135_0));
   INV_X1 i_2_135_2 (.A(n_240), .ZN(n_2_135_1));
   OAI21_X1 i_2_136_0 (.A(n_2_136_0), .B1(n_2_339), .B2(n_2_136_1), .ZN(n_2_174));
   AOI21_X1 i_2_136_1 (.A(n_236), .B1(n_2_339), .B2(n_234), .ZN(n_2_136_0));
   INV_X1 i_2_136_2 (.A(n_235), .ZN(n_2_136_1));
   OAI21_X1 i_2_137_0 (.A(n_2_137_0), .B1(n_2_339), .B2(n_2_137_1), .ZN(n_2_180));
   AOI21_X1 i_2_137_1 (.A(n_215), .B1(n_2_339), .B2(n_213), .ZN(n_2_137_0));
   INV_X1 i_2_137_2 (.A(n_214), .ZN(n_2_137_1));
   OAI21_X1 i_2_138_0 (.A(n_2_138_0), .B1(n_2_339), .B2(n_2_138_1), .ZN(n_2_184));
   AOI21_X1 i_2_138_1 (.A(n_207), .B1(n_2_339), .B2(n_205), .ZN(n_2_138_0));
   INV_X1 i_2_138_2 (.A(n_206), .ZN(n_2_138_1));
   OAI21_X1 i_2_139_0 (.A(n_2_139_0), .B1(n_2_339), .B2(n_2_139_1), .ZN(n_2_185));
   AOI21_X1 i_2_139_1 (.A(n_204), .B1(n_2_339), .B2(n_202), .ZN(n_2_139_0));
   INV_X1 i_2_139_2 (.A(n_203), .ZN(n_2_139_1));
   OAI21_X1 i_2_140_0 (.A(n_2_140_0), .B1(n_2_339), .B2(n_2_140_1), .ZN(n_2_188));
   AOI21_X1 i_2_140_1 (.A(n_201), .B1(n_2_339), .B2(n_199), .ZN(n_2_140_0));
   INV_X1 i_2_140_2 (.A(n_200), .ZN(n_2_140_1));
   OAI21_X1 i_2_141_0 (.A(n_2_141_0), .B1(n_2_339), .B2(n_2_141_1), .ZN(n_2_194));
   AOI21_X1 i_2_141_1 (.A(n_183), .B1(n_2_339), .B2(n_181), .ZN(n_2_141_0));
   INV_X1 i_2_141_2 (.A(n_182), .ZN(n_2_141_1));
   OAI21_X1 i_2_142_0 (.A(n_2_142_0), .B1(n_2_339), .B2(n_2_142_1), .ZN(n_2_196));
   AOI21_X1 i_2_142_1 (.A(n_173), .B1(n_2_339), .B2(n_171), .ZN(n_2_142_0));
   INV_X1 i_2_142_2 (.A(n_172), .ZN(n_2_142_1));
   OAI21_X1 i_2_143_0 (.A(n_2_143_0), .B1(n_2_339), .B2(n_2_143_1), .ZN(n_2_197));
   AOI21_X1 i_2_143_1 (.A(n_168), .B1(n_2_339), .B2(n_166), .ZN(n_2_143_0));
   INV_X1 i_2_143_2 (.A(n_167), .ZN(n_2_143_1));
   OAI21_X1 i_2_144_0 (.A(n_2_144_0), .B1(n_2_339), .B2(n_2_144_1), .ZN(n_2_198));
   AOI21_X1 i_2_144_1 (.A(n_163), .B1(n_2_339), .B2(n_161), .ZN(n_2_144_0));
   INV_X1 i_2_144_2 (.A(n_162), .ZN(n_2_144_1));
   OAI21_X1 i_2_145_0 (.A(n_2_145_0), .B1(n_2_339), .B2(n_2_145_1), .ZN(n_2_201));
   AOI21_X1 i_2_145_1 (.A(n_157), .B1(n_2_339), .B2(n_155), .ZN(n_2_145_0));
   INV_X1 i_2_145_2 (.A(n_156), .ZN(n_2_145_1));
   OAI21_X1 i_2_146_0 (.A(n_2_146_0), .B1(n_2_339), .B2(n_2_146_1), .ZN(n_2_202));
   AOI21_X1 i_2_146_1 (.A(n_152), .B1(n_2_339), .B2(n_150), .ZN(n_2_146_0));
   INV_X1 i_2_146_2 (.A(n_151), .ZN(n_2_146_1));
   OAI21_X1 i_2_147_0 (.A(n_2_147_0), .B1(n_2_339), .B2(n_2_147_1), .ZN(n_2_203));
   AOI21_X1 i_2_147_1 (.A(n_149), .B1(n_2_339), .B2(n_147), .ZN(n_2_147_0));
   INV_X1 i_2_147_2 (.A(n_148), .ZN(n_2_147_1));
   OAI21_X1 i_2_148_0 (.A(n_2_148_0), .B1(n_2_339), .B2(n_2_148_1), .ZN(n_2_205));
   AOI21_X1 i_2_148_1 (.A(n_141), .B1(n_2_339), .B2(n_139), .ZN(n_2_148_0));
   INV_X1 i_2_148_2 (.A(n_140), .ZN(n_2_148_1));
   OAI21_X1 i_2_149_0 (.A(n_2_149_0), .B1(n_2_149_3), .B2(n_2_149_1), .ZN(
      n_2_225));
   NAND2_X1 i_2_149_1 (.A1(n_10), .A2(n_2_149_1), .ZN(n_2_149_0));
   OAI22_X1 i_2_149_2 (.A1(n_2_339), .A2(n_214), .B1(n_2_149_2), .B2(n_213), 
      .ZN(n_2_149_1));
   INV_X1 i_2_149_3 (.A(n_2_339), .ZN(n_2_149_2));
   INV_X1 i_2_149_4 (.A(in_data[8]), .ZN(n_2_149_3));
   OAI21_X1 i_2_150_0 (.A(n_2_150_0), .B1(n_2_150_3), .B2(n_2_150_1), .ZN(
      n_2_226));
   NAND2_X1 i_2_150_1 (.A1(n_8), .A2(n_2_150_1), .ZN(n_2_150_0));
   OAI22_X1 i_2_150_2 (.A1(n_2_339), .A2(n_203), .B1(n_2_150_2), .B2(n_202), 
      .ZN(n_2_150_1));
   INV_X1 i_2_150_3 (.A(n_2_339), .ZN(n_2_150_2));
   INV_X1 i_2_150_4 (.A(in_data[8]), .ZN(n_2_150_3));
   OAI21_X1 i_2_151_0 (.A(n_2_151_0), .B1(n_2_151_3), .B2(n_2_151_1), .ZN(
      n_2_227));
   NAND2_X1 i_2_151_1 (.A1(n_7), .A2(n_2_151_1), .ZN(n_2_151_0));
   OAI22_X1 i_2_151_2 (.A1(n_2_339), .A2(n_200), .B1(n_2_151_2), .B2(n_199), 
      .ZN(n_2_151_1));
   INV_X1 i_2_151_3 (.A(n_2_339), .ZN(n_2_151_2));
   INV_X1 i_2_151_4 (.A(in_data[8]), .ZN(n_2_151_3));
   OAI21_X1 i_2_152_0 (.A(n_2_152_0), .B1(n_2_152_3), .B2(n_2_152_1), .ZN(
      n_2_228));
   NAND2_X1 i_2_152_1 (.A1(n_6), .A2(n_2_152_1), .ZN(n_2_152_0));
   OAI22_X1 i_2_152_2 (.A1(n_2_339), .A2(n_162), .B1(n_2_152_2), .B2(n_161), 
      .ZN(n_2_152_1));
   INV_X1 i_2_152_3 (.A(n_2_339), .ZN(n_2_152_2));
   INV_X1 i_2_152_4 (.A(in_data[8]), .ZN(n_2_152_3));
   datapath__1_13509 i_2_153 (.\out_as[5] (\out_as[5] ), .\out_bs[5] ({n_844, 
      n_2_368, n_848, n_846, n_849, n_2_371, \out_bs[5] [0]}), .p_0(n_1089));
   OAI21_X1 i_2_154_0 (.A(n_2_154_0), .B1(n_2_154_3), .B2(n_2_154_1), .ZN(n_1090));
   NAND2_X1 i_2_154_1 (.A1(n_9), .A2(n_2_154_1), .ZN(n_2_154_0));
   OAI22_X1 i_2_154_2 (.A1(n_2_339), .A2(n_206), .B1(n_2_154_2), .B2(n_205), 
      .ZN(n_2_154_1));
   INV_X1 i_2_154_3 (.A(n_2_339), .ZN(n_2_154_2));
   INV_X1 i_2_154_4 (.A(in_data[8]), .ZN(n_2_154_3));
   OR2_X1 i_2_155_0 (.A1(n_852), .A2(n_727), .ZN(n_2_241));
   BUF_X1 rt_shieldBuf__5__5__0 (.A(n_1089), .Z(n_2_339));
   OAI21_X1 i_2_156_0 (.A(n_2_156_0), .B1(n_2_156_3), .B2(n_2_156_1), .ZN(n_1091));
   NAND2_X1 i_2_156_1 (.A1(n_127), .A2(n_2_156_1), .ZN(n_2_156_0));
   OAI22_X1 i_2_156_2 (.A1(n_952), .A2(n_2_3), .B1(n_2_156_2), .B2(n_2_2), 
      .ZN(n_2_156_1));
   INV_X1 i_2_156_3 (.A(n_952), .ZN(n_2_156_2));
   INV_X1 i_2_156_4 (.A(in_data[4]), .ZN(n_2_156_3));
   OAI21_X1 i_2_157_0 (.A(n_2_157_0), .B1(n_2_157_3), .B2(n_2_157_1), .ZN(n_1092));
   NAND2_X1 i_2_157_1 (.A1(n_125), .A2(n_2_157_1), .ZN(n_2_157_0));
   OAI22_X1 i_2_157_2 (.A1(n_952), .A2(n_2_7), .B1(n_2_157_2), .B2(n_2_6), 
      .ZN(n_2_157_1));
   INV_X1 i_2_157_3 (.A(n_952), .ZN(n_2_157_2));
   INV_X1 i_2_157_4 (.A(in_data[4]), .ZN(n_2_157_3));
   OAI21_X1 i_2_158_0 (.A(n_2_158_0), .B1(n_2_158_3), .B2(n_2_158_1), .ZN(n_1093));
   NAND2_X1 i_2_158_1 (.A1(n_123), .A2(n_2_158_1), .ZN(n_2_158_0));
   OAI22_X1 i_2_158_2 (.A1(n_952), .A2(n_644), .B1(n_2_158_2), .B2(n_643), 
      .ZN(n_2_158_1));
   INV_X1 i_2_158_3 (.A(n_952), .ZN(n_2_158_2));
   INV_X1 i_2_158_4 (.A(in_data[4]), .ZN(n_2_158_3));
   OAI21_X1 i_2_159_0 (.A(n_2_159_0), .B1(n_2_159_3), .B2(n_2_159_1), .ZN(n_1094));
   NAND2_X1 i_2_159_1 (.A1(n_122), .A2(n_2_159_1), .ZN(n_2_159_0));
   OAI22_X1 i_2_159_2 (.A1(n_952), .A2(n_2_12), .B1(n_2_159_2), .B2(n_2_11), 
      .ZN(n_2_159_1));
   INV_X1 i_2_159_3 (.A(n_952), .ZN(n_2_159_2));
   INV_X1 i_2_159_4 (.A(in_data[4]), .ZN(n_2_159_3));
   OAI21_X1 i_2_160_0 (.A(n_2_160_0), .B1(n_2_160_3), .B2(n_2_160_1), .ZN(n_1095));
   NAND2_X1 i_2_160_1 (.A1(n_121), .A2(n_2_160_1), .ZN(n_2_160_0));
   OAI22_X1 i_2_160_2 (.A1(n_952), .A2(n_2_15), .B1(n_2_160_2), .B2(n_2_14), 
      .ZN(n_2_160_1));
   INV_X1 i_2_160_3 (.A(n_952), .ZN(n_2_160_2));
   INV_X1 i_2_160_4 (.A(in_data[4]), .ZN(n_2_160_3));
   OAI21_X1 i_2_161_0 (.A(n_2_161_0), .B1(n_2_161_3), .B2(n_2_161_1), .ZN(n_1096));
   NAND2_X1 i_2_161_1 (.A1(n_119), .A2(n_2_161_1), .ZN(n_2_161_0));
   OAI22_X1 i_2_161_2 (.A1(n_952), .A2(n_2_19), .B1(n_2_161_2), .B2(n_2_18), 
      .ZN(n_2_161_1));
   INV_X1 i_2_161_3 (.A(n_952), .ZN(n_2_161_2));
   INV_X1 i_2_161_4 (.A(in_data[4]), .ZN(n_2_161_3));
   OAI21_X1 i_2_162_0 (.A(n_2_162_0), .B1(n_2_162_3), .B2(n_2_162_1), .ZN(n_1097));
   NAND2_X1 i_2_162_1 (.A1(n_116), .A2(n_2_162_1), .ZN(n_2_162_0));
   OAI22_X1 i_2_162_2 (.A1(n_952), .A2(n_2_24), .B1(n_2_162_2), .B2(n_2_23), 
      .ZN(n_2_162_1));
   INV_X1 i_2_162_3 (.A(n_952), .ZN(n_2_162_2));
   INV_X1 i_2_162_4 (.A(in_data[4]), .ZN(n_2_162_3));
   OAI21_X1 i_2_163_0 (.A(n_2_163_0), .B1(n_2_163_3), .B2(n_2_163_1), .ZN(n_1098));
   NAND2_X1 i_2_163_1 (.A1(n_114), .A2(n_2_163_1), .ZN(n_2_163_0));
   OAI22_X1 i_2_163_2 (.A1(n_952), .A2(n_597), .B1(n_2_163_2), .B2(n_596), 
      .ZN(n_2_163_1));
   INV_X1 i_2_163_3 (.A(n_952), .ZN(n_2_163_2));
   INV_X1 i_2_163_4 (.A(in_data[4]), .ZN(n_2_163_3));
   OAI21_X1 i_2_164_0 (.A(n_2_164_0), .B1(n_2_164_3), .B2(n_2_164_1), .ZN(n_1099));
   NAND2_X1 i_2_164_1 (.A1(n_113), .A2(n_2_164_1), .ZN(n_2_164_0));
   OAI22_X1 i_2_164_2 (.A1(n_952), .A2(n_2_34), .B1(n_2_164_2), .B2(n_2_33), 
      .ZN(n_2_164_1));
   INV_X1 i_2_164_3 (.A(n_952), .ZN(n_2_164_2));
   INV_X1 i_2_164_4 (.A(in_data[4]), .ZN(n_2_164_3));
   OAI21_X1 i_2_165_0 (.A(n_2_165_0), .B1(n_2_165_3), .B2(n_2_165_1), .ZN(n_1100));
   NAND2_X1 i_2_165_1 (.A1(n_112), .A2(n_2_165_1), .ZN(n_2_165_0));
   OAI22_X1 i_2_165_2 (.A1(n_952), .A2(n_2_37), .B1(n_2_165_2), .B2(n_2_36), 
      .ZN(n_2_165_1));
   INV_X1 i_2_165_3 (.A(n_952), .ZN(n_2_165_2));
   INV_X1 i_2_165_4 (.A(in_data[4]), .ZN(n_2_165_3));
   OAI21_X1 i_2_166_0 (.A(n_2_166_0), .B1(n_2_166_3), .B2(n_2_166_1), .ZN(n_1101));
   NAND2_X1 i_2_166_1 (.A1(n_833), .A2(n_2_166_1), .ZN(n_2_166_0));
   OAI22_X1 i_2_166_2 (.A1(n_952), .A2(n_2_40), .B1(n_2_166_2), .B2(n_2_39), 
      .ZN(n_2_166_1));
   INV_X1 i_2_166_3 (.A(n_952), .ZN(n_2_166_2));
   INV_X1 i_2_166_4 (.A(in_data[4]), .ZN(n_2_166_3));
   OAI21_X1 i_2_167_0 (.A(n_2_167_0), .B1(n_2_167_3), .B2(n_2_167_1), .ZN(n_1102));
   NAND2_X1 i_2_167_1 (.A1(n_111), .A2(n_2_167_1), .ZN(n_2_167_0));
   OAI22_X1 i_2_167_2 (.A1(n_952), .A2(n_2_43), .B1(n_2_167_2), .B2(n_2_42), 
      .ZN(n_2_167_1));
   INV_X1 i_2_167_3 (.A(n_952), .ZN(n_2_167_2));
   INV_X1 i_2_167_4 (.A(in_data[4]), .ZN(n_2_167_3));
   OAI21_X1 i_2_168_0 (.A(n_2_168_0), .B1(n_2_168_3), .B2(n_2_168_1), .ZN(n_1103));
   NAND2_X1 i_2_168_1 (.A1(n_110), .A2(n_2_168_1), .ZN(n_2_168_0));
   OAI22_X1 i_2_168_2 (.A1(n_952), .A2(n_2_46), .B1(n_2_168_2), .B2(n_2_45), 
      .ZN(n_2_168_1));
   INV_X1 i_2_168_3 (.A(n_952), .ZN(n_2_168_2));
   INV_X1 i_2_168_4 (.A(in_data[4]), .ZN(n_2_168_3));
   OAI21_X1 i_2_169_0 (.A(n_2_169_0), .B1(n_2_169_3), .B2(n_2_169_1), .ZN(n_1104));
   NAND2_X1 i_2_169_1 (.A1(n_109), .A2(n_2_169_1), .ZN(n_2_169_0));
   OAI22_X1 i_2_169_2 (.A1(n_952), .A2(n_2_52), .B1(n_2_169_2), .B2(n_2_51), 
      .ZN(n_2_169_1));
   INV_X1 i_2_169_3 (.A(n_952), .ZN(n_2_169_2));
   INV_X1 i_2_169_4 (.A(in_data[4]), .ZN(n_2_169_3));
   OAI21_X1 i_2_170_0 (.A(n_2_170_0), .B1(n_2_170_3), .B2(n_2_170_1), .ZN(n_1105));
   NAND2_X1 i_2_170_1 (.A1(n_108), .A2(n_2_170_1), .ZN(n_2_170_0));
   OAI22_X1 i_2_170_2 (.A1(n_952), .A2(n_2_58), .B1(n_2_170_2), .B2(n_2_57), 
      .ZN(n_2_170_1));
   INV_X1 i_2_170_3 (.A(n_952), .ZN(n_2_170_2));
   INV_X1 i_2_170_4 (.A(in_data[4]), .ZN(n_2_170_3));
   OAI21_X1 i_2_171_0 (.A(n_2_171_0), .B1(n_2_171_3), .B2(n_2_171_1), .ZN(n_1106));
   NAND2_X1 i_2_171_1 (.A1(n_106), .A2(n_2_171_1), .ZN(n_2_171_0));
   OAI22_X1 i_2_171_2 (.A1(n_952), .A2(n_2_66), .B1(n_2_171_2), .B2(n_2_65), 
      .ZN(n_2_171_1));
   INV_X1 i_2_171_3 (.A(n_952), .ZN(n_2_171_2));
   INV_X1 i_2_171_4 (.A(in_data[4]), .ZN(n_2_171_3));
   OAI21_X1 i_2_172_0 (.A(n_2_172_0), .B1(n_2_172_3), .B2(n_2_172_1), .ZN(n_1107));
   NAND2_X1 i_2_172_1 (.A1(n_105), .A2(n_2_172_1), .ZN(n_2_172_0));
   OAI22_X1 i_2_172_2 (.A1(n_952), .A2(n_543), .B1(n_2_172_2), .B2(n_542), 
      .ZN(n_2_172_1));
   INV_X1 i_2_172_3 (.A(n_952), .ZN(n_2_172_2));
   INV_X1 i_2_172_4 (.A(in_data[4]), .ZN(n_2_172_3));
   OAI21_X1 i_2_173_0 (.A(n_2_173_0), .B1(n_2_173_3), .B2(n_2_173_1), .ZN(n_1108));
   NAND2_X1 i_2_173_1 (.A1(n_104), .A2(n_2_173_1), .ZN(n_2_173_0));
   OAI22_X1 i_2_173_2 (.A1(n_952), .A2(n_538), .B1(n_2_173_2), .B2(n_537), 
      .ZN(n_2_173_1));
   INV_X1 i_2_173_3 (.A(n_952), .ZN(n_2_173_2));
   INV_X1 i_2_173_4 (.A(in_data[4]), .ZN(n_2_173_3));
   OAI21_X1 i_2_174_0 (.A(n_2_174_0), .B1(n_2_174_3), .B2(n_2_174_1), .ZN(n_1109));
   NAND2_X1 i_2_174_1 (.A1(n_103), .A2(n_2_174_1), .ZN(n_2_174_0));
   OAI22_X1 i_2_174_2 (.A1(n_952), .A2(n_533), .B1(n_2_174_2), .B2(n_532), 
      .ZN(n_2_174_1));
   INV_X1 i_2_174_3 (.A(n_952), .ZN(n_2_174_2));
   INV_X1 i_2_174_4 (.A(in_data[4]), .ZN(n_2_174_3));
   OAI21_X1 i_2_175_0 (.A(n_2_175_0), .B1(n_2_175_3), .B2(n_2_175_1), .ZN(n_1110));
   NAND2_X1 i_2_175_1 (.A1(n_100), .A2(n_2_175_1), .ZN(n_2_175_0));
   OAI22_X1 i_2_175_2 (.A1(n_952), .A2(n_513), .B1(n_2_175_2), .B2(n_512), 
      .ZN(n_2_175_1));
   INV_X1 i_2_175_3 (.A(n_952), .ZN(n_2_175_2));
   INV_X1 i_2_175_4 (.A(in_data[4]), .ZN(n_2_175_3));
   OAI21_X1 i_2_176_0 (.A(n_2_176_0), .B1(n_2_176_3), .B2(n_2_176_1), .ZN(n_1111));
   NAND2_X1 i_2_176_1 (.A1(n_98), .A2(n_2_176_1), .ZN(n_2_176_0));
   OAI22_X1 i_2_176_2 (.A1(n_952), .A2(n_498), .B1(n_2_176_2), .B2(n_497), 
      .ZN(n_2_176_1));
   INV_X1 i_2_176_3 (.A(n_952), .ZN(n_2_176_2));
   INV_X1 i_2_176_4 (.A(in_data[4]), .ZN(n_2_176_3));
   OAI21_X1 i_2_177_0 (.A(n_2_177_0), .B1(n_2_177_3), .B2(n_2_177_1), .ZN(n_1112));
   NAND2_X1 i_2_177_1 (.A1(n_97), .A2(n_2_177_1), .ZN(n_2_177_0));
   OAI22_X1 i_2_177_2 (.A1(n_952), .A2(n_493), .B1(n_2_177_2), .B2(n_492), 
      .ZN(n_2_177_1));
   INV_X1 i_2_177_3 (.A(n_952), .ZN(n_2_177_2));
   INV_X1 i_2_177_4 (.A(in_data[4]), .ZN(n_2_177_3));
   OAI21_X1 i_2_178_0 (.A(n_2_178_0), .B1(n_2_178_3), .B2(n_2_178_1), .ZN(n_1113));
   NAND2_X1 i_2_178_1 (.A1(n_96), .A2(n_2_178_1), .ZN(n_2_178_0));
   OAI22_X1 i_2_178_2 (.A1(n_952), .A2(n_488), .B1(n_2_178_2), .B2(n_487), 
      .ZN(n_2_178_1));
   INV_X1 i_2_178_3 (.A(n_952), .ZN(n_2_178_2));
   INV_X1 i_2_178_4 (.A(in_data[4]), .ZN(n_2_178_3));
   OAI21_X1 i_2_179_0 (.A(n_2_179_0), .B1(n_2_179_3), .B2(n_2_179_1), .ZN(n_1114));
   NAND2_X1 i_2_179_1 (.A1(n_94), .A2(n_2_179_1), .ZN(n_2_179_0));
   OAI22_X1 i_2_179_2 (.A1(n_952), .A2(n_456), .B1(n_2_179_2), .B2(n_455), 
      .ZN(n_2_179_1));
   INV_X1 i_2_179_3 (.A(n_952), .ZN(n_2_179_2));
   INV_X1 i_2_179_4 (.A(in_data[4]), .ZN(n_2_179_3));
   OAI21_X1 i_2_180_0 (.A(n_2_180_0), .B1(n_2_180_3), .B2(n_2_180_1), .ZN(n_1115));
   NAND2_X1 i_2_180_1 (.A1(n_93), .A2(n_2_180_1), .ZN(n_2_180_0));
   OAI22_X1 i_2_180_2 (.A1(n_952), .A2(n_451), .B1(n_2_180_2), .B2(n_450), 
      .ZN(n_2_180_1));
   INV_X1 i_2_180_3 (.A(n_952), .ZN(n_2_180_2));
   INV_X1 i_2_180_4 (.A(in_data[4]), .ZN(n_2_180_3));
   OAI21_X1 i_2_181_0 (.A(n_2_181_0), .B1(n_2_181_3), .B2(n_2_181_1), .ZN(n_1116));
   NAND2_X1 i_2_181_1 (.A1(n_92), .A2(n_2_181_1), .ZN(n_2_181_0));
   OAI22_X1 i_2_181_2 (.A1(n_952), .A2(n_446), .B1(n_2_181_2), .B2(n_445), 
      .ZN(n_2_181_1));
   INV_X1 i_2_181_3 (.A(n_952), .ZN(n_2_181_2));
   INV_X1 i_2_181_4 (.A(in_data[4]), .ZN(n_2_181_3));
   OAI21_X1 i_2_182_0 (.A(n_2_182_0), .B1(n_2_182_3), .B2(n_2_182_1), .ZN(n_1117));
   NAND2_X1 i_2_182_1 (.A1(n_91), .A2(n_2_182_1), .ZN(n_2_182_0));
   OAI22_X1 i_2_182_2 (.A1(n_952), .A2(n_440), .B1(n_2_182_2), .B2(n_2_95), 
      .ZN(n_2_182_1));
   INV_X1 i_2_182_3 (.A(n_952), .ZN(n_2_182_2));
   INV_X1 i_2_182_4 (.A(in_data[4]), .ZN(n_2_182_3));
   OAI21_X1 i_2_183_0 (.A(n_2_183_0), .B1(n_2_183_3), .B2(n_2_183_1), .ZN(n_1118));
   NAND2_X1 i_2_183_1 (.A1(n_90), .A2(n_2_183_1), .ZN(n_2_183_0));
   OAI22_X1 i_2_183_2 (.A1(n_952), .A2(n_436), .B1(n_2_183_2), .B2(n_435), 
      .ZN(n_2_183_1));
   INV_X1 i_2_183_3 (.A(n_952), .ZN(n_2_183_2));
   INV_X1 i_2_183_4 (.A(in_data[4]), .ZN(n_2_183_3));
   OAI21_X1 i_2_184_0 (.A(n_2_184_0), .B1(n_2_184_3), .B2(n_2_184_1), .ZN(n_1119));
   NAND2_X1 i_2_184_1 (.A1(n_89), .A2(n_2_184_1), .ZN(n_2_184_0));
   OAI22_X1 i_2_184_2 (.A1(n_952), .A2(n_2_99), .B1(n_2_184_2), .B2(n_2_98), 
      .ZN(n_2_184_1));
   INV_X1 i_2_184_3 (.A(n_952), .ZN(n_2_184_2));
   INV_X1 i_2_184_4 (.A(in_data[4]), .ZN(n_2_184_3));
   OAI21_X1 i_2_185_0 (.A(n_2_185_0), .B1(n_2_185_3), .B2(n_2_185_1), .ZN(n_1120));
   NAND2_X1 i_2_185_1 (.A1(n_88), .A2(n_2_185_1), .ZN(n_2_185_0));
   OAI22_X1 i_2_185_2 (.A1(n_952), .A2(n_427), .B1(n_2_185_2), .B2(n_426), 
      .ZN(n_2_185_1));
   INV_X1 i_2_185_3 (.A(n_952), .ZN(n_2_185_2));
   INV_X1 i_2_185_4 (.A(in_data[4]), .ZN(n_2_185_3));
   OAI21_X1 i_2_186_0 (.A(n_2_186_0), .B1(n_2_186_3), .B2(n_2_186_1), .ZN(n_1121));
   NAND2_X1 i_2_186_1 (.A1(n_87), .A2(n_2_186_1), .ZN(n_2_186_0));
   OAI22_X1 i_2_186_2 (.A1(n_952), .A2(n_422), .B1(n_2_186_2), .B2(n_421), 
      .ZN(n_2_186_1));
   INV_X1 i_2_186_3 (.A(n_952), .ZN(n_2_186_2));
   INV_X1 i_2_186_4 (.A(in_data[4]), .ZN(n_2_186_3));
   OAI21_X1 i_2_187_0 (.A(n_2_187_0), .B1(n_2_187_3), .B2(n_2_187_1), .ZN(n_1122));
   NAND2_X1 i_2_187_1 (.A1(n_86), .A2(n_2_187_1), .ZN(n_2_187_0));
   OAI22_X1 i_2_187_2 (.A1(n_952), .A2(n_417), .B1(n_2_187_2), .B2(n_416), 
      .ZN(n_2_187_1));
   INV_X1 i_2_187_3 (.A(n_952), .ZN(n_2_187_2));
   INV_X1 i_2_187_4 (.A(in_data[4]), .ZN(n_2_187_3));
   OAI21_X1 i_2_188_0 (.A(n_2_188_0), .B1(n_2_188_3), .B2(n_2_188_1), .ZN(n_1123));
   NAND2_X1 i_2_188_1 (.A1(n_85), .A2(n_2_188_1), .ZN(n_2_188_0));
   OAI22_X1 i_2_188_2 (.A1(n_952), .A2(n_412), .B1(n_2_188_2), .B2(n_411), 
      .ZN(n_2_188_1));
   INV_X1 i_2_188_3 (.A(n_952), .ZN(n_2_188_2));
   INV_X1 i_2_188_4 (.A(in_data[4]), .ZN(n_2_188_3));
   OAI21_X1 i_2_189_0 (.A(n_2_189_0), .B1(n_2_189_3), .B2(n_2_189_1), .ZN(n_1124));
   NAND2_X1 i_2_189_1 (.A1(n_83), .A2(n_2_189_1), .ZN(n_2_189_0));
   OAI22_X1 i_2_189_2 (.A1(n_952), .A2(n_402), .B1(n_2_189_2), .B2(n_401), 
      .ZN(n_2_189_1));
   INV_X1 i_2_189_3 (.A(n_952), .ZN(n_2_189_2));
   INV_X1 i_2_189_4 (.A(in_data[4]), .ZN(n_2_189_3));
   OAI21_X1 i_2_190_0 (.A(n_2_190_0), .B1(n_2_190_3), .B2(n_2_190_1), .ZN(n_1125));
   NAND2_X1 i_2_190_1 (.A1(n_82), .A2(n_2_190_1), .ZN(n_2_190_0));
   OAI22_X1 i_2_190_2 (.A1(n_952), .A2(n_397), .B1(n_2_190_2), .B2(n_396), 
      .ZN(n_2_190_1));
   INV_X1 i_2_190_3 (.A(n_952), .ZN(n_2_190_2));
   INV_X1 i_2_190_4 (.A(in_data[4]), .ZN(n_2_190_3));
   OAI21_X1 i_2_191_0 (.A(n_2_191_0), .B1(n_2_191_3), .B2(n_2_191_1), .ZN(n_1126));
   NAND2_X1 i_2_191_1 (.A1(n_81), .A2(n_2_191_1), .ZN(n_2_191_0));
   OAI22_X1 i_2_191_2 (.A1(n_952), .A2(n_2_111), .B1(n_2_191_2), .B2(n_2_110), 
      .ZN(n_2_191_1));
   INV_X1 i_2_191_3 (.A(n_952), .ZN(n_2_191_2));
   INV_X1 i_2_191_4 (.A(in_data[4]), .ZN(n_2_191_3));
   OAI21_X1 i_2_192_0 (.A(n_2_192_0), .B1(n_2_192_3), .B2(n_2_192_1), .ZN(n_1127));
   NAND2_X1 i_2_192_1 (.A1(n_80), .A2(n_2_192_1), .ZN(n_2_192_0));
   OAI22_X1 i_2_192_2 (.A1(n_952), .A2(n_379), .B1(n_2_192_2), .B2(n_378), 
      .ZN(n_2_192_1));
   INV_X1 i_2_192_3 (.A(n_952), .ZN(n_2_192_2));
   INV_X1 i_2_192_4 (.A(in_data[4]), .ZN(n_2_192_3));
   OAI21_X1 i_2_193_0 (.A(n_2_193_0), .B1(n_2_193_3), .B2(n_2_193_1), .ZN(n_1128));
   NAND2_X1 i_2_193_1 (.A1(n_79), .A2(n_2_193_1), .ZN(n_2_193_0));
   OAI22_X1 i_2_193_2 (.A1(n_952), .A2(n_2_115), .B1(n_2_193_2), .B2(n_2_114), 
      .ZN(n_2_193_1));
   INV_X1 i_2_193_3 (.A(n_952), .ZN(n_2_193_2));
   INV_X1 i_2_193_4 (.A(in_data[4]), .ZN(n_2_193_3));
   OAI21_X1 i_2_194_0 (.A(n_2_194_0), .B1(n_2_194_3), .B2(n_2_194_1), .ZN(n_1129));
   NAND2_X1 i_2_194_1 (.A1(n_78), .A2(n_2_194_1), .ZN(n_2_194_0));
   OAI22_X1 i_2_194_2 (.A1(n_952), .A2(n_368), .B1(n_2_194_2), .B2(n_367), 
      .ZN(n_2_194_1));
   INV_X1 i_2_194_3 (.A(n_952), .ZN(n_2_194_2));
   INV_X1 i_2_194_4 (.A(in_data[4]), .ZN(n_2_194_3));
   OAI21_X1 i_2_195_0 (.A(n_2_195_0), .B1(n_2_195_3), .B2(n_2_195_1), .ZN(n_1130));
   NAND2_X1 i_2_195_1 (.A1(n_77), .A2(n_2_195_1), .ZN(n_2_195_0));
   OAI22_X1 i_2_195_2 (.A1(n_952), .A2(n_363), .B1(n_2_195_2), .B2(n_362), 
      .ZN(n_2_195_1));
   INV_X1 i_2_195_3 (.A(n_952), .ZN(n_2_195_2));
   INV_X1 i_2_195_4 (.A(in_data[4]), .ZN(n_2_195_3));
   OAI21_X1 i_2_196_0 (.A(n_2_196_0), .B1(n_2_196_3), .B2(n_2_196_1), .ZN(n_1131));
   NAND2_X1 i_2_196_1 (.A1(n_76), .A2(n_2_196_1), .ZN(n_2_196_0));
   OAI22_X1 i_2_196_2 (.A1(n_952), .A2(n_358), .B1(n_2_196_2), .B2(n_357), 
      .ZN(n_2_196_1));
   INV_X1 i_2_196_3 (.A(n_952), .ZN(n_2_196_2));
   INV_X1 i_2_196_4 (.A(in_data[4]), .ZN(n_2_196_3));
   OAI21_X1 i_2_197_0 (.A(n_2_197_0), .B1(n_2_197_3), .B2(n_2_197_1), .ZN(n_1132));
   NAND2_X1 i_2_197_1 (.A1(n_75), .A2(n_2_197_1), .ZN(n_2_197_0));
   OAI22_X1 i_2_197_2 (.A1(n_952), .A2(n_353), .B1(n_2_197_2), .B2(n_352), 
      .ZN(n_2_197_1));
   INV_X1 i_2_197_3 (.A(n_952), .ZN(n_2_197_2));
   INV_X1 i_2_197_4 (.A(in_data[4]), .ZN(n_2_197_3));
   OAI21_X1 i_2_198_0 (.A(n_2_198_0), .B1(n_2_198_3), .B2(n_2_198_1), .ZN(n_1133));
   NAND2_X1 i_2_198_1 (.A1(n_74), .A2(n_2_198_1), .ZN(n_2_198_0));
   OAI22_X1 i_2_198_2 (.A1(n_952), .A2(n_2_125), .B1(n_2_198_2), .B2(n_2_124), 
      .ZN(n_2_198_1));
   INV_X1 i_2_198_3 (.A(n_952), .ZN(n_2_198_2));
   INV_X1 i_2_198_4 (.A(in_data[4]), .ZN(n_2_198_3));
   OAI21_X1 i_2_199_0 (.A(n_2_199_0), .B1(n_2_199_3), .B2(n_2_199_1), .ZN(n_1134));
   NAND2_X1 i_2_199_1 (.A1(n_73), .A2(n_2_199_1), .ZN(n_2_199_0));
   OAI22_X1 i_2_199_2 (.A1(n_952), .A2(n_345), .B1(n_2_199_2), .B2(n_344), 
      .ZN(n_2_199_1));
   INV_X1 i_2_199_3 (.A(n_952), .ZN(n_2_199_2));
   INV_X1 i_2_199_4 (.A(in_data[4]), .ZN(n_2_199_3));
   OAI21_X1 i_2_200_0 (.A(n_2_200_0), .B1(n_2_200_3), .B2(n_2_200_1), .ZN(n_1135));
   NAND2_X1 i_2_200_1 (.A1(n_72), .A2(n_2_200_1), .ZN(n_2_200_0));
   OAI22_X1 i_2_200_2 (.A1(n_952), .A2(n_340), .B1(n_2_200_2), .B2(n_339), 
      .ZN(n_2_200_1));
   INV_X1 i_2_200_3 (.A(n_952), .ZN(n_2_200_2));
   INV_X1 i_2_200_4 (.A(in_data[4]), .ZN(n_2_200_3));
   OAI21_X1 i_2_201_0 (.A(n_2_201_0), .B1(n_2_201_3), .B2(n_2_201_1), .ZN(n_1136));
   NAND2_X1 i_2_201_1 (.A1(n_71), .A2(n_2_201_1), .ZN(n_2_201_0));
   OAI22_X1 i_2_201_2 (.A1(n_952), .A2(n_2_131), .B1(n_2_201_2), .B2(n_2_130), 
      .ZN(n_2_201_1));
   INV_X1 i_2_201_3 (.A(n_952), .ZN(n_2_201_2));
   INV_X1 i_2_201_4 (.A(in_data[4]), .ZN(n_2_201_3));
   OAI21_X1 i_2_202_0 (.A(n_2_202_0), .B1(n_2_202_3), .B2(n_2_202_1), .ZN(n_1137));
   NAND2_X1 i_2_202_1 (.A1(n_70), .A2(n_2_202_1), .ZN(n_2_202_0));
   OAI22_X1 i_2_202_2 (.A1(n_952), .A2(n_2_134), .B1(n_2_202_2), .B2(n_2_133), 
      .ZN(n_2_202_1));
   INV_X1 i_2_202_3 (.A(n_952), .ZN(n_2_202_2));
   INV_X1 i_2_202_4 (.A(in_data[4]), .ZN(n_2_202_3));
   OAI21_X1 i_2_203_0 (.A(n_2_203_0), .B1(n_2_203_3), .B2(n_2_203_1), .ZN(n_1138));
   NAND2_X1 i_2_203_1 (.A1(n_69), .A2(n_2_203_1), .ZN(n_2_203_0));
   OAI22_X1 i_2_203_2 (.A1(n_952), .A2(n_2_137), .B1(n_2_203_2), .B2(n_2_136), 
      .ZN(n_2_203_1));
   INV_X1 i_2_203_3 (.A(n_952), .ZN(n_2_203_2));
   INV_X1 i_2_203_4 (.A(in_data[4]), .ZN(n_2_203_3));
   OAI21_X1 i_2_204_0 (.A(n_2_204_0), .B1(n_2_204_3), .B2(n_2_204_1), .ZN(n_1139));
   NAND2_X1 i_2_204_1 (.A1(n_68), .A2(n_2_204_1), .ZN(n_2_204_0));
   OAI22_X1 i_2_204_2 (.A1(n_952), .A2(n_321), .B1(n_2_204_2), .B2(n_320), 
      .ZN(n_2_204_1));
   INV_X1 i_2_204_3 (.A(n_952), .ZN(n_2_204_2));
   INV_X1 i_2_204_4 (.A(in_data[4]), .ZN(n_2_204_3));
   OAI21_X1 i_2_205_0 (.A(n_2_205_0), .B1(n_2_205_3), .B2(n_2_205_1), .ZN(n_1140));
   NAND2_X1 i_2_205_1 (.A1(n_67), .A2(n_2_205_1), .ZN(n_2_205_0));
   OAI22_X1 i_2_205_2 (.A1(n_952), .A2(n_2_141), .B1(n_2_205_2), .B2(n_2_140), 
      .ZN(n_2_205_1));
   INV_X1 i_2_205_3 (.A(n_952), .ZN(n_2_205_2));
   INV_X1 i_2_205_4 (.A(in_data[4]), .ZN(n_2_205_3));
   OAI21_X1 i_2_206_0 (.A(n_2_206_0), .B1(n_2_206_3), .B2(n_2_206_1), .ZN(n_1141));
   NAND2_X1 i_2_206_1 (.A1(n_66), .A2(n_2_206_1), .ZN(n_2_206_0));
   OAI22_X1 i_2_206_2 (.A1(n_952), .A2(n_313), .B1(n_2_206_2), .B2(n_312), 
      .ZN(n_2_206_1));
   INV_X1 i_2_206_3 (.A(n_952), .ZN(n_2_206_2));
   INV_X1 i_2_206_4 (.A(in_data[4]), .ZN(n_2_206_3));
   OAI21_X1 i_2_207_0 (.A(n_2_207_0), .B1(n_2_207_3), .B2(n_2_207_1), .ZN(n_1142));
   NAND2_X1 i_2_207_1 (.A1(n_65), .A2(n_2_207_1), .ZN(n_2_207_0));
   OAI22_X1 i_2_207_2 (.A1(n_952), .A2(n_2_145), .B1(n_2_207_2), .B2(n_2_144), 
      .ZN(n_2_207_1));
   INV_X1 i_2_207_3 (.A(n_952), .ZN(n_2_207_2));
   INV_X1 i_2_207_4 (.A(in_data[4]), .ZN(n_2_207_3));
   OAI21_X1 i_2_208_0 (.A(n_2_208_0), .B1(n_2_208_3), .B2(n_2_208_1), .ZN(n_1143));
   NAND2_X1 i_2_208_1 (.A1(n_64), .A2(n_2_208_1), .ZN(n_2_208_0));
   OAI22_X1 i_2_208_2 (.A1(n_952), .A2(n_305), .B1(n_2_208_2), .B2(n_304), 
      .ZN(n_2_208_1));
   INV_X1 i_2_208_3 (.A(n_952), .ZN(n_2_208_2));
   INV_X1 i_2_208_4 (.A(in_data[4]), .ZN(n_2_208_3));
   OAI21_X1 i_2_209_0 (.A(n_2_209_0), .B1(n_2_209_3), .B2(n_2_209_1), .ZN(n_1144));
   NAND2_X1 i_2_209_1 (.A1(n_63), .A2(n_2_209_1), .ZN(n_2_209_0));
   OAI22_X1 i_2_209_2 (.A1(n_952), .A2(n_2_149), .B1(n_2_209_2), .B2(n_2_148), 
      .ZN(n_2_209_1));
   INV_X1 i_2_209_3 (.A(n_952), .ZN(n_2_209_2));
   INV_X1 i_2_209_4 (.A(in_data[4]), .ZN(n_2_209_3));
   OAI21_X1 i_2_210_0 (.A(n_2_210_0), .B1(n_2_210_3), .B2(n_2_210_1), .ZN(n_1145));
   NAND2_X1 i_2_210_1 (.A1(n_62), .A2(n_2_210_1), .ZN(n_2_210_0));
   OAI22_X1 i_2_210_2 (.A1(n_952), .A2(n_2_152), .B1(n_2_210_2), .B2(n_2_151), 
      .ZN(n_2_210_1));
   INV_X1 i_2_210_3 (.A(n_952), .ZN(n_2_210_2));
   INV_X1 i_2_210_4 (.A(in_data[4]), .ZN(n_2_210_3));
   OAI21_X1 i_2_211_0 (.A(n_2_211_0), .B1(n_2_211_3), .B2(n_2_211_1), .ZN(n_1146));
   NAND2_X1 i_2_211_1 (.A1(n_61), .A2(n_2_211_1), .ZN(n_2_211_0));
   OAI22_X1 i_2_211_2 (.A1(n_952), .A2(n_2_155), .B1(n_2_211_2), .B2(n_2_154), 
      .ZN(n_2_211_1));
   INV_X1 i_2_211_3 (.A(n_952), .ZN(n_2_211_2));
   INV_X1 i_2_211_4 (.A(in_data[4]), .ZN(n_2_211_3));
   OAI21_X1 i_2_212_0 (.A(n_2_212_0), .B1(n_2_212_3), .B2(n_2_212_1), .ZN(n_1147));
   NAND2_X1 i_2_212_1 (.A1(n_60), .A2(n_2_212_1), .ZN(n_2_212_0));
   OAI22_X1 i_2_212_2 (.A1(n_952), .A2(n_291), .B1(n_2_212_2), .B2(n_290), 
      .ZN(n_2_212_1));
   INV_X1 i_2_212_3 (.A(n_952), .ZN(n_2_212_2));
   INV_X1 i_2_212_4 (.A(in_data[4]), .ZN(n_2_212_3));
   OAI21_X1 i_2_213_0 (.A(n_2_213_0), .B1(n_2_213_3), .B2(n_2_213_1), .ZN(n_1148));
   NAND2_X1 i_2_213_1 (.A1(n_59), .A2(n_2_213_1), .ZN(n_2_213_0));
   OAI22_X1 i_2_213_2 (.A1(n_952), .A2(n_2_159), .B1(n_2_213_2), .B2(n_2_158), 
      .ZN(n_2_213_1));
   INV_X1 i_2_213_3 (.A(n_952), .ZN(n_2_213_2));
   INV_X1 i_2_213_4 (.A(in_data[4]), .ZN(n_2_213_3));
   OAI21_X1 i_2_214_0 (.A(n_2_214_0), .B1(n_2_214_3), .B2(n_2_214_1), .ZN(n_1149));
   NAND2_X1 i_2_214_1 (.A1(n_58), .A2(n_2_214_1), .ZN(n_2_214_0));
   OAI22_X1 i_2_214_2 (.A1(n_952), .A2(n_277), .B1(n_2_214_2), .B2(n_276), 
      .ZN(n_2_214_1));
   INV_X1 i_2_214_3 (.A(n_952), .ZN(n_2_214_2));
   INV_X1 i_2_214_4 (.A(in_data[4]), .ZN(n_2_214_3));
   OAI21_X1 i_2_215_0 (.A(n_2_215_0), .B1(n_2_215_3), .B2(n_2_215_1), .ZN(n_1150));
   NAND2_X1 i_2_215_1 (.A1(n_57), .A2(n_2_215_1), .ZN(n_2_215_0));
   OAI22_X1 i_2_215_2 (.A1(n_952), .A2(n_267), .B1(n_2_215_2), .B2(n_266), 
      .ZN(n_2_215_1));
   INV_X1 i_2_215_3 (.A(n_952), .ZN(n_2_215_2));
   INV_X1 i_2_215_4 (.A(in_data[4]), .ZN(n_2_215_3));
   OAI21_X1 i_2_216_0 (.A(n_2_216_0), .B1(n_2_216_3), .B2(n_2_216_1), .ZN(n_1151));
   NAND2_X1 i_2_216_1 (.A1(n_56), .A2(n_2_216_1), .ZN(n_2_216_0));
   OAI22_X1 i_2_216_2 (.A1(n_952), .A2(n_256), .B1(n_2_216_2), .B2(n_255), 
      .ZN(n_2_216_1));
   INV_X1 i_2_216_3 (.A(n_952), .ZN(n_2_216_2));
   INV_X1 i_2_216_4 (.A(in_data[4]), .ZN(n_2_216_3));
   OAI21_X1 i_2_217_0 (.A(n_2_217_0), .B1(n_2_217_3), .B2(n_2_217_1), .ZN(n_1152));
   NAND2_X1 i_2_217_1 (.A1(n_55), .A2(n_2_217_1), .ZN(n_2_217_0));
   OAI22_X1 i_2_217_2 (.A1(n_952), .A2(n_248), .B1(n_2_217_2), .B2(n_247), 
      .ZN(n_2_217_1));
   INV_X1 i_2_217_3 (.A(n_952), .ZN(n_2_217_2));
   INV_X1 i_2_217_4 (.A(in_data[4]), .ZN(n_2_217_3));
   OAI21_X1 i_2_218_0 (.A(n_2_218_0), .B1(n_2_218_3), .B2(n_2_218_1), .ZN(n_1153));
   NAND2_X1 i_2_218_1 (.A1(n_54), .A2(n_2_218_1), .ZN(n_2_218_0));
   OAI22_X1 i_2_218_2 (.A1(n_952), .A2(n_238), .B1(n_2_218_2), .B2(n_237), 
      .ZN(n_2_218_1));
   INV_X1 i_2_218_3 (.A(n_952), .ZN(n_2_218_2));
   INV_X1 i_2_218_4 (.A(in_data[4]), .ZN(n_2_218_3));
   OAI21_X1 i_2_219_0 (.A(n_2_219_0), .B1(n_2_219_3), .B2(n_2_219_1), .ZN(n_1154));
   NAND2_X1 i_2_219_1 (.A1(n_53), .A2(n_2_219_1), .ZN(n_2_219_0));
   OAI22_X1 i_2_219_2 (.A1(n_952), .A2(n_233), .B1(n_2_219_2), .B2(n_232), 
      .ZN(n_2_219_1));
   INV_X1 i_2_219_3 (.A(n_952), .ZN(n_2_219_2));
   INV_X1 i_2_219_4 (.A(in_data[4]), .ZN(n_2_219_3));
   OAI21_X1 i_2_220_0 (.A(n_2_220_0), .B1(n_2_220_3), .B2(n_2_220_1), .ZN(n_1155));
   NAND2_X1 i_2_220_1 (.A1(n_52), .A2(n_2_220_1), .ZN(n_2_220_0));
   OAI22_X1 i_2_220_2 (.A1(n_952), .A2(n_228), .B1(n_2_220_2), .B2(n_227), 
      .ZN(n_2_220_1));
   INV_X1 i_2_220_3 (.A(n_952), .ZN(n_2_220_2));
   INV_X1 i_2_220_4 (.A(in_data[4]), .ZN(n_2_220_3));
   OAI21_X1 i_2_221_0 (.A(n_2_221_0), .B1(n_2_221_3), .B2(n_2_221_1), .ZN(n_1156));
   NAND2_X1 i_2_221_1 (.A1(n_51), .A2(n_2_221_1), .ZN(n_2_221_0));
   OAI22_X1 i_2_221_2 (.A1(n_952), .A2(n_222), .B1(n_2_221_2), .B2(n_221), 
      .ZN(n_2_221_1));
   INV_X1 i_2_221_3 (.A(n_952), .ZN(n_2_221_2));
   INV_X1 i_2_221_4 (.A(in_data[4]), .ZN(n_2_221_3));
   OAI21_X1 i_2_222_0 (.A(n_2_222_0), .B1(n_2_222_3), .B2(n_2_222_1), .ZN(n_1157));
   NAND2_X1 i_2_222_1 (.A1(n_50), .A2(n_2_222_1), .ZN(n_2_222_0));
   OAI22_X1 i_2_222_2 (.A1(n_952), .A2(n_217), .B1(n_2_222_2), .B2(n_216), 
      .ZN(n_2_222_1));
   INV_X1 i_2_222_3 (.A(n_952), .ZN(n_2_222_2));
   INV_X1 i_2_222_4 (.A(in_data[4]), .ZN(n_2_222_3));
   OAI21_X1 i_2_223_0 (.A(n_2_223_0), .B1(n_2_223_3), .B2(n_2_223_1), .ZN(n_1158));
   NAND2_X1 i_2_223_1 (.A1(n_49), .A2(n_2_223_1), .ZN(n_2_223_0));
   OAI22_X1 i_2_223_2 (.A1(n_952), .A2(n_209), .B1(n_2_223_2), .B2(n_208), 
      .ZN(n_2_223_1));
   INV_X1 i_2_223_3 (.A(n_952), .ZN(n_2_223_2));
   INV_X1 i_2_223_4 (.A(in_data[4]), .ZN(n_2_223_3));
   OAI21_X1 i_2_224_0 (.A(n_2_224_0), .B1(n_2_224_3), .B2(n_2_224_1), .ZN(n_1159));
   NAND2_X1 i_2_224_1 (.A1(n_48), .A2(n_2_224_1), .ZN(n_2_224_0));
   OAI22_X1 i_2_224_2 (.A1(n_952), .A2(n_195), .B1(n_2_224_2), .B2(n_194), 
      .ZN(n_2_224_1));
   INV_X1 i_2_224_3 (.A(n_952), .ZN(n_2_224_2));
   INV_X1 i_2_224_4 (.A(in_data[4]), .ZN(n_2_224_3));
   OAI21_X1 i_2_225_0 (.A(n_2_225_0), .B1(n_2_225_3), .B2(n_2_225_1), .ZN(n_1160));
   NAND2_X1 i_2_225_1 (.A1(n_47), .A2(n_2_225_1), .ZN(n_2_225_0));
   OAI22_X1 i_2_225_2 (.A1(n_952), .A2(n_190), .B1(n_2_225_2), .B2(n_189), 
      .ZN(n_2_225_1));
   INV_X1 i_2_225_3 (.A(n_952), .ZN(n_2_225_2));
   INV_X1 i_2_225_4 (.A(in_data[4]), .ZN(n_2_225_3));
   OAI21_X1 i_2_226_0 (.A(n_2_226_0), .B1(n_2_226_3), .B2(n_2_226_1), .ZN(n_1161));
   NAND2_X1 i_2_226_1 (.A1(n_46), .A2(n_2_226_1), .ZN(n_2_226_0));
   OAI22_X1 i_2_226_2 (.A1(n_952), .A2(n_185), .B1(n_2_226_2), .B2(n_184), 
      .ZN(n_2_226_1));
   INV_X1 i_2_226_3 (.A(n_952), .ZN(n_2_226_2));
   INV_X1 i_2_226_4 (.A(in_data[4]), .ZN(n_2_226_3));
   OAI21_X1 i_2_227_0 (.A(n_2_227_0), .B1(n_2_227_3), .B2(n_2_227_1), .ZN(n_1162));
   NAND2_X1 i_2_227_1 (.A1(n_45), .A2(n_2_227_1), .ZN(n_2_227_0));
   OAI22_X1 i_2_227_2 (.A1(n_952), .A2(n_180), .B1(n_2_227_2), .B2(n_179), 
      .ZN(n_2_227_1));
   INV_X1 i_2_227_3 (.A(n_952), .ZN(n_2_227_2));
   INV_X1 i_2_227_4 (.A(in_data[4]), .ZN(n_2_227_3));
   OAI21_X1 i_2_228_0 (.A(n_2_228_0), .B1(n_2_228_3), .B2(n_2_228_1), .ZN(n_1163));
   NAND2_X1 i_2_228_1 (.A1(n_44), .A2(n_2_228_1), .ZN(n_2_228_0));
   OAI22_X1 i_2_228_2 (.A1(n_952), .A2(n_175), .B1(n_2_228_2), .B2(n_174), 
      .ZN(n_2_228_1));
   INV_X1 i_2_228_3 (.A(n_952), .ZN(n_2_228_2));
   INV_X1 i_2_228_4 (.A(in_data[4]), .ZN(n_2_228_3));
   OAI21_X1 i_2_229_0 (.A(n_2_229_0), .B1(n_2_229_3), .B2(n_2_229_1), .ZN(n_1164));
   NAND2_X1 i_2_229_1 (.A1(n_43), .A2(n_2_229_1), .ZN(n_2_229_0));
   OAI22_X1 i_2_229_2 (.A1(n_952), .A2(n_170), .B1(n_2_229_2), .B2(n_169), 
      .ZN(n_2_229_1));
   INV_X1 i_2_229_3 (.A(n_952), .ZN(n_2_229_2));
   INV_X1 i_2_229_4 (.A(in_data[4]), .ZN(n_2_229_3));
   OAI21_X1 i_2_230_0 (.A(n_2_230_0), .B1(n_2_230_3), .B2(n_2_230_1), .ZN(n_1165));
   NAND2_X1 i_2_230_1 (.A1(n_42), .A2(n_2_230_1), .ZN(n_2_230_0));
   OAI22_X1 i_2_230_2 (.A1(n_952), .A2(n_165), .B1(n_2_230_2), .B2(n_164), 
      .ZN(n_2_230_1));
   INV_X1 i_2_230_3 (.A(n_952), .ZN(n_2_230_2));
   INV_X1 i_2_230_4 (.A(in_data[4]), .ZN(n_2_230_3));
   OAI21_X1 i_2_231_0 (.A(n_2_231_0), .B1(n_2_231_3), .B2(n_2_231_1), .ZN(n_1166));
   NAND2_X1 i_2_231_1 (.A1(n_41), .A2(n_2_231_1), .ZN(n_2_231_0));
   OAI22_X1 i_2_231_2 (.A1(n_952), .A2(n_159), .B1(n_2_231_2), .B2(n_158), 
      .ZN(n_2_231_1));
   INV_X1 i_2_231_3 (.A(n_952), .ZN(n_2_231_2));
   INV_X1 i_2_231_4 (.A(in_data[4]), .ZN(n_2_231_3));
   OAI21_X1 i_2_232_0 (.A(n_2_232_0), .B1(n_2_232_3), .B2(n_2_232_1), .ZN(n_1167));
   NAND2_X1 i_2_232_1 (.A1(n_40), .A2(n_2_232_1), .ZN(n_2_232_0));
   OAI22_X1 i_2_232_2 (.A1(n_952), .A2(n_154), .B1(n_2_232_2), .B2(n_153), 
      .ZN(n_2_232_1));
   INV_X1 i_2_232_3 (.A(n_952), .ZN(n_2_232_2));
   INV_X1 i_2_232_4 (.A(in_data[4]), .ZN(n_2_232_3));
   OAI21_X1 i_2_233_0 (.A(n_2_233_0), .B1(n_2_233_3), .B2(n_2_233_1), .ZN(n_1168));
   NAND2_X1 i_2_233_1 (.A1(n_39), .A2(n_2_233_1), .ZN(n_2_233_0));
   OAI22_X1 i_2_233_2 (.A1(n_952), .A2(n_143), .B1(n_2_233_2), .B2(n_142), 
      .ZN(n_2_233_1));
   INV_X1 i_2_233_3 (.A(n_952), .ZN(n_2_233_2));
   INV_X1 i_2_233_4 (.A(in_data[4]), .ZN(n_2_233_3));
   OAI21_X1 i_2_234_0 (.A(n_2_234_0), .B1(n_2_234_3), .B2(n_2_234_1), .ZN(n_1169));
   NAND2_X1 i_2_234_1 (.A1(n_38), .A2(n_2_234_1), .ZN(n_2_234_0));
   OAI22_X1 i_2_234_2 (.A1(n_952), .A2(n_2_206), .B1(n_2_234_2), .B2(n_138), 
      .ZN(n_2_234_1));
   INV_X1 i_2_234_3 (.A(n_952), .ZN(n_2_234_2));
   INV_X1 i_2_234_4 (.A(in_data[4]), .ZN(n_2_234_3));
   OAI21_X1 i_2_235_0 (.A(n_2_235_0), .B1(n_2_235_3), .B2(n_2_235_1), .ZN(n_1170));
   NAND2_X1 i_2_235_1 (.A1(n_37), .A2(n_2_235_1), .ZN(n_2_235_0));
   OAI22_X1 i_2_235_2 (.A1(n_952), .A2(n_134), .B1(n_2_235_2), .B2(n_133), 
      .ZN(n_2_235_1));
   INV_X1 i_2_235_3 (.A(n_952), .ZN(n_2_235_2));
   INV_X1 i_2_235_4 (.A(in_data[4]), .ZN(n_2_235_3));
   OAI21_X1 i_2_236_0 (.A(n_2_236_0), .B1(n_2_236_3), .B2(n_2_236_1), .ZN(n_2_0));
   NAND2_X1 i_2_236_1 (.A1(n_3), .A2(n_2_236_1), .ZN(n_2_236_0));
   NOR2_X1 i_2_236_2 (.A1(n_2_236_2), .A2(n_130), .ZN(n_2_236_1));
   INV_X1 i_2_236_3 (.A(n_952), .ZN(n_2_236_2));
   INV_X1 i_2_236_4 (.A(in_data[4]), .ZN(n_2_236_3));
   OAI21_X1 i_2_237_0 (.A(n_2_237_0), .B1(n_2_237_3), .B2(n_2_237_1), .ZN(n_1171));
   NAND2_X1 i_2_237_1 (.A1(n_11), .A2(n_2_237_1), .ZN(n_2_237_0));
   OAI22_X1 i_2_237_2 (.A1(n_952), .A2(n_2_177), .B1(n_2_237_2), .B2(n_2_176), 
      .ZN(n_2_237_1));
   INV_X1 i_2_237_3 (.A(n_952), .ZN(n_2_237_2));
   INV_X1 i_2_237_4 (.A(in_data[4]), .ZN(n_2_237_3));
   OAI21_X1 i_2_238_0 (.A(n_2_238_0), .B1(n_2_238_3), .B2(n_2_238_1), .ZN(n_1172));
   NAND2_X1 i_2_238_1 (.A1(n_2_224), .A2(n_2_238_1), .ZN(n_2_238_0));
   OAI22_X1 i_2_238_2 (.A1(n_952), .A2(n_243), .B1(n_2_238_2), .B2(n_242), 
      .ZN(n_2_238_1));
   INV_X1 i_2_238_3 (.A(n_952), .ZN(n_2_238_2));
   INV_X1 i_2_238_4 (.A(in_data[4]), .ZN(n_2_238_3));
   OAI21_X1 i_2_239_0 (.A(n_2_239_0), .B1(n_2_239_3), .B2(n_2_239_1), .ZN(n_1173));
   NAND2_X1 i_2_239_1 (.A1(n_2_223), .A2(n_2_239_1), .ZN(n_2_239_0));
   OAI22_X1 i_2_239_2 (.A1(n_952), .A2(n_2_170), .B1(n_2_239_2), .B2(n_2_169), 
      .ZN(n_2_239_1));
   INV_X1 i_2_239_3 (.A(n_952), .ZN(n_2_239_2));
   INV_X1 i_2_239_4 (.A(in_data[4]), .ZN(n_2_239_3));
   OAI21_X1 i_2_240_0 (.A(n_2_240_0), .B1(n_2_240_3), .B2(n_2_240_1), .ZN(n_1174));
   NAND2_X1 i_2_240_1 (.A1(n_14), .A2(n_2_240_1), .ZN(n_2_240_0));
   OAI22_X1 i_2_240_2 (.A1(n_952), .A2(n_2_166), .B1(n_2_240_2), .B2(n_2_165), 
      .ZN(n_2_240_1));
   INV_X1 i_2_240_3 (.A(n_952), .ZN(n_2_240_2));
   INV_X1 i_2_240_4 (.A(in_data[4]), .ZN(n_2_240_3));
   OAI21_X1 i_2_241_0 (.A(n_2_241_0), .B1(n_2_241_3), .B2(n_2_241_1), .ZN(n_1175));
   NAND2_X1 i_2_241_1 (.A1(n_2_222), .A2(n_2_241_1), .ZN(n_2_241_0));
   OAI22_X1 i_2_241_2 (.A1(n_952), .A2(n_272), .B1(n_2_241_2), .B2(n_271), 
      .ZN(n_2_241_1));
   INV_X1 i_2_241_3 (.A(n_952), .ZN(n_2_241_2));
   INV_X1 i_2_241_4 (.A(in_data[4]), .ZN(n_2_241_3));
   OAI21_X1 i_2_242_0 (.A(n_2_242_0), .B1(n_2_242_3), .B2(n_2_242_1), .ZN(n_1176));
   NAND2_X1 i_2_242_1 (.A1(n_2_221), .A2(n_2_242_1), .ZN(n_2_242_0));
   OAI22_X1 i_2_242_2 (.A1(n_952), .A2(n_283), .B1(n_2_242_2), .B2(n_282), 
      .ZN(n_2_242_1));
   INV_X1 i_2_242_3 (.A(n_952), .ZN(n_2_242_2));
   INV_X1 i_2_242_4 (.A(in_data[4]), .ZN(n_2_242_3));
   OAI21_X1 i_2_243_0 (.A(n_2_243_0), .B1(n_2_243_3), .B2(n_2_243_1), .ZN(n_1177));
   NAND2_X1 i_2_243_1 (.A1(n_2_220), .A2(n_2_243_1), .ZN(n_2_243_0));
   OAI22_X1 i_2_243_2 (.A1(n_952), .A2(n_335), .B1(n_2_243_2), .B2(n_334), 
      .ZN(n_2_243_1));
   INV_X1 i_2_243_3 (.A(n_952), .ZN(n_2_243_2));
   INV_X1 i_2_243_4 (.A(in_data[4]), .ZN(n_2_243_3));
   OAI21_X1 i_2_244_0 (.A(n_2_244_0), .B1(n_2_244_3), .B2(n_2_244_1), .ZN(n_1178));
   NAND2_X1 i_2_244_1 (.A1(n_2_219), .A2(n_2_244_1), .ZN(n_2_244_0));
   OAI22_X1 i_2_244_2 (.A1(n_952), .A2(n_2_118), .B1(n_2_244_2), .B2(n_2_117), 
      .ZN(n_2_244_1));
   INV_X1 i_2_244_3 (.A(n_952), .ZN(n_2_244_2));
   INV_X1 i_2_244_4 (.A(in_data[4]), .ZN(n_2_244_3));
   OAI21_X1 i_2_245_0 (.A(n_2_245_0), .B1(n_2_245_3), .B2(n_2_245_1), .ZN(n_1179));
   NAND2_X1 i_2_245_1 (.A1(n_2_218), .A2(n_2_245_1), .ZN(n_2_245_0));
   OAI22_X1 i_2_245_2 (.A1(n_952), .A2(n_392), .B1(n_2_245_2), .B2(n_391), 
      .ZN(n_2_245_1));
   INV_X1 i_2_245_3 (.A(n_952), .ZN(n_2_245_2));
   INV_X1 i_2_245_4 (.A(in_data[4]), .ZN(n_2_245_3));
   OAI21_X1 i_2_246_0 (.A(n_2_246_0), .B1(n_2_246_3), .B2(n_2_246_1), .ZN(n_1180));
   NAND2_X1 i_2_246_1 (.A1(n_2_217), .A2(n_2_246_1), .ZN(n_2_246_0));
   OAI22_X1 i_2_246_2 (.A1(n_952), .A2(n_2_88), .B1(n_2_246_2), .B2(n_2_87), 
      .ZN(n_2_246_1));
   INV_X1 i_2_246_3 (.A(n_952), .ZN(n_2_246_2));
   INV_X1 i_2_246_4 (.A(in_data[4]), .ZN(n_2_246_3));
   OAI21_X1 i_2_247_0 (.A(n_2_247_0), .B1(n_2_247_3), .B2(n_2_247_1), .ZN(n_1181));
   NAND2_X1 i_2_247_1 (.A1(n_2_216), .A2(n_2_247_1), .ZN(n_2_247_0));
   OAI22_X1 i_2_247_2 (.A1(n_952), .A2(n_2_85), .B1(n_2_247_2), .B2(n_2_84), 
      .ZN(n_2_247_1));
   INV_X1 i_2_247_3 (.A(n_952), .ZN(n_2_247_2));
   INV_X1 i_2_247_4 (.A(in_data[4]), .ZN(n_2_247_3));
   OAI21_X1 i_2_248_0 (.A(n_2_248_0), .B1(n_2_248_3), .B2(n_2_248_1), .ZN(n_1182));
   NAND2_X1 i_2_248_1 (.A1(n_2_215), .A2(n_2_248_1), .ZN(n_2_248_0));
   OAI22_X1 i_2_248_2 (.A1(n_952), .A2(n_2_82), .B1(n_2_248_2), .B2(n_2_81), 
      .ZN(n_2_248_1));
   INV_X1 i_2_248_3 (.A(n_952), .ZN(n_2_248_2));
   INV_X1 i_2_248_4 (.A(in_data[4]), .ZN(n_2_248_3));
   OAI21_X1 i_2_249_0 (.A(n_2_249_0), .B1(n_2_249_3), .B2(n_2_249_1), .ZN(n_1183));
   NAND2_X1 i_2_249_1 (.A1(n_2_214), .A2(n_2_249_1), .ZN(n_2_249_0));
   OAI22_X1 i_2_249_2 (.A1(n_952), .A2(n_483), .B1(n_2_249_2), .B2(n_482), 
      .ZN(n_2_249_1));
   INV_X1 i_2_249_3 (.A(n_952), .ZN(n_2_249_2));
   INV_X1 i_2_249_4 (.A(in_data[4]), .ZN(n_2_249_3));
   OAI21_X1 i_2_250_0 (.A(n_2_250_0), .B1(n_2_250_3), .B2(n_2_250_1), .ZN(n_1184));
   NAND2_X1 i_2_250_1 (.A1(n_2_213), .A2(n_2_250_1), .ZN(n_2_250_0));
   OAI22_X1 i_2_250_2 (.A1(n_952), .A2(n_503), .B1(n_2_250_2), .B2(n_502), 
      .ZN(n_2_250_1));
   INV_X1 i_2_250_3 (.A(n_952), .ZN(n_2_250_2));
   INV_X1 i_2_250_4 (.A(in_data[4]), .ZN(n_2_250_3));
   OAI21_X1 i_2_251_0 (.A(n_2_251_0), .B1(n_2_251_3), .B2(n_2_251_1), .ZN(n_1185));
   NAND2_X1 i_2_251_1 (.A1(n_2_212), .A2(n_2_251_1), .ZN(n_2_251_0));
   OAI22_X1 i_2_251_2 (.A1(n_952), .A2(n_518), .B1(n_2_251_2), .B2(n_517), 
      .ZN(n_2_251_1));
   INV_X1 i_2_251_3 (.A(n_952), .ZN(n_2_251_2));
   INV_X1 i_2_251_4 (.A(in_data[4]), .ZN(n_2_251_3));
   OAI21_X1 i_2_252_0 (.A(n_2_252_0), .B1(n_2_252_3), .B2(n_2_252_1), .ZN(n_1186));
   NAND2_X1 i_2_252_1 (.A1(n_2_211), .A2(n_2_252_1), .ZN(n_2_252_0));
   OAI22_X1 i_2_252_2 (.A1(n_952), .A2(n_2_62), .B1(n_2_252_2), .B2(n_2_61), 
      .ZN(n_2_252_1));
   INV_X1 i_2_252_3 (.A(n_952), .ZN(n_2_252_2));
   INV_X1 i_2_252_4 (.A(in_data[4]), .ZN(n_2_252_3));
   OAI21_X1 i_2_253_0 (.A(n_2_253_0), .B1(n_2_253_3), .B2(n_2_253_1), .ZN(n_1187));
   NAND2_X1 i_2_253_1 (.A1(n_2_210), .A2(n_2_253_1), .ZN(n_2_253_0));
   OAI22_X1 i_2_253_2 (.A1(n_952), .A2(n_2_55), .B1(n_2_253_2), .B2(n_2_54), 
      .ZN(n_2_253_1));
   INV_X1 i_2_253_3 (.A(n_952), .ZN(n_2_253_2));
   INV_X1 i_2_253_4 (.A(in_data[4]), .ZN(n_2_253_3));
   OAI21_X1 i_2_254_0 (.A(n_2_254_0), .B1(n_2_254_3), .B2(n_2_254_1), .ZN(n_1188));
   NAND2_X1 i_2_254_1 (.A1(n_2_209), .A2(n_2_254_1), .ZN(n_2_254_0));
   OAI22_X1 i_2_254_2 (.A1(n_952), .A2(n_2_49), .B1(n_2_254_2), .B2(n_2_48), 
      .ZN(n_2_254_1));
   INV_X1 i_2_254_3 (.A(n_952), .ZN(n_2_254_2));
   INV_X1 i_2_254_4 (.A(in_data[4]), .ZN(n_2_254_3));
   OAI21_X1 i_2_255_0 (.A(n_2_255_0), .B1(n_2_255_3), .B2(n_2_255_1), .ZN(n_1189));
   NAND2_X1 i_2_255_1 (.A1(n_2_208), .A2(n_2_255_1), .ZN(n_2_255_0));
   OAI22_X1 i_2_255_2 (.A1(n_952), .A2(n_2_30), .B1(n_2_255_2), .B2(n_2_29), 
      .ZN(n_2_255_1));
   INV_X1 i_2_255_3 (.A(n_952), .ZN(n_2_255_2));
   INV_X1 i_2_255_4 (.A(in_data[4]), .ZN(n_2_255_3));
   OAI21_X1 i_2_256_0 (.A(n_2_256_0), .B1(n_2_256_3), .B2(n_2_256_1), .ZN(n_1190));
   NAND2_X1 i_2_256_1 (.A1(n_36), .A2(n_2_256_1), .ZN(n_2_256_0));
   OAI22_X1 i_2_256_2 (.A1(n_2_369), .A2(n_614), .B1(n_2_256_2), .B2(n_613), 
      .ZN(n_2_256_1));
   INV_X1 i_2_256_3 (.A(n_2_369), .ZN(n_2_256_2));
   INV_X1 i_2_256_4 (.A(in_data[8]), .ZN(n_2_256_3));
   OAI21_X1 i_2_257_0 (.A(n_2_257_0), .B1(n_2_257_3), .B2(n_2_257_1), .ZN(n_1191));
   NAND2_X1 i_2_257_1 (.A1(n_35), .A2(n_2_257_1), .ZN(n_2_257_0));
   OAI22_X1 i_2_257_2 (.A1(n_2_369), .A2(n_607), .B1(n_2_257_2), .B2(n_606), 
      .ZN(n_2_257_1));
   INV_X1 i_2_257_3 (.A(n_2_369), .ZN(n_2_257_2));
   INV_X1 i_2_257_4 (.A(in_data[8]), .ZN(n_2_257_3));
   OAI21_X1 i_2_258_0 (.A(n_2_258_0), .B1(n_2_258_3), .B2(n_2_258_1), .ZN(
      n_2_208));
   NAND2_X1 i_2_258_1 (.A1(n_34), .A2(n_2_258_1), .ZN(n_2_258_0));
   OAI22_X1 i_2_258_2 (.A1(n_2_369), .A2(n_603), .B1(n_2_258_2), .B2(n_602), 
      .ZN(n_2_258_1));
   INV_X1 i_2_258_3 (.A(n_2_369), .ZN(n_2_258_2));
   INV_X1 i_2_258_4 (.A(in_data[8]), .ZN(n_2_258_3));
   OAI21_X1 i_2_259_0 (.A(n_2_259_0), .B1(n_2_259_3), .B2(n_2_259_1), .ZN(
      n_2_209));
   NAND2_X1 i_2_259_1 (.A1(n_33), .A2(n_2_259_1), .ZN(n_2_259_0));
   OAI22_X1 i_2_259_2 (.A1(n_2_369), .A2(n_576), .B1(n_2_259_2), .B2(n_575), 
      .ZN(n_2_259_1));
   INV_X1 i_2_259_3 (.A(n_2_369), .ZN(n_2_259_2));
   INV_X1 i_2_259_4 (.A(in_data[8]), .ZN(n_2_259_3));
   OAI21_X1 i_2_260_0 (.A(n_2_260_0), .B1(n_2_260_3), .B2(n_2_260_1), .ZN(
      n_2_210));
   NAND2_X1 i_2_260_1 (.A1(n_32), .A2(n_2_260_1), .ZN(n_2_260_0));
   OAI22_X1 i_2_260_2 (.A1(n_2_369), .A2(n_568), .B1(n_2_260_2), .B2(n_567), 
      .ZN(n_2_260_1));
   INV_X1 i_2_260_3 (.A(n_2_369), .ZN(n_2_260_2));
   INV_X1 i_2_260_4 (.A(in_data[8]), .ZN(n_2_260_3));
   OAI21_X1 i_2_261_0 (.A(n_2_261_0), .B1(n_2_261_3), .B2(n_2_261_1), .ZN(n_1192));
   NAND2_X1 i_2_261_1 (.A1(n_31), .A2(n_2_261_1), .ZN(n_2_261_0));
   OAI22_X1 i_2_261_2 (.A1(n_2_369), .A2(n_560), .B1(n_2_261_2), .B2(n_559), 
      .ZN(n_2_261_1));
   INV_X1 i_2_261_3 (.A(n_2_369), .ZN(n_2_261_2));
   INV_X1 i_2_261_4 (.A(in_data[8]), .ZN(n_2_261_3));
   OAI21_X1 i_2_262_0 (.A(n_2_262_0), .B1(n_2_262_3), .B2(n_2_262_1), .ZN(
      n_2_211));
   NAND2_X1 i_2_262_1 (.A1(n_30), .A2(n_2_262_1), .ZN(n_2_262_0));
   OAI22_X1 i_2_262_2 (.A1(n_2_369), .A2(n_556), .B1(n_2_262_2), .B2(n_555), 
      .ZN(n_2_262_1));
   INV_X1 i_2_262_3 (.A(n_2_369), .ZN(n_2_262_2));
   INV_X1 i_2_262_4 (.A(in_data[8]), .ZN(n_2_262_3));
   OAI21_X1 i_2_263_0 (.A(n_2_263_0), .B1(n_2_263_3), .B2(n_2_263_1), .ZN(
      n_2_212));
   NAND2_X1 i_2_263_1 (.A1(n_29), .A2(n_2_263_1), .ZN(n_2_263_0));
   OAI22_X1 i_2_263_2 (.A1(n_2_369), .A2(n_520), .B1(n_2_263_2), .B2(n_519), 
      .ZN(n_2_263_1));
   INV_X1 i_2_263_3 (.A(n_2_369), .ZN(n_2_263_2));
   INV_X1 i_2_263_4 (.A(in_data[8]), .ZN(n_2_263_3));
   OAI21_X1 i_2_264_0 (.A(n_2_264_0), .B1(n_2_264_3), .B2(n_2_264_1), .ZN(
      n_2_213));
   NAND2_X1 i_2_264_1 (.A1(n_28), .A2(n_2_264_1), .ZN(n_2_264_0));
   OAI22_X1 i_2_264_2 (.A1(n_2_369), .A2(n_505), .B1(n_2_264_2), .B2(n_504), 
      .ZN(n_2_264_1));
   INV_X1 i_2_264_3 (.A(n_2_369), .ZN(n_2_264_2));
   INV_X1 i_2_264_4 (.A(in_data[8]), .ZN(n_2_264_3));
   OAI21_X1 i_2_265_0 (.A(n_2_265_0), .B1(n_2_265_3), .B2(n_2_265_1), .ZN(
      n_2_214));
   NAND2_X1 i_2_265_1 (.A1(n_27), .A2(n_2_265_1), .ZN(n_2_265_0));
   OAI22_X1 i_2_265_2 (.A1(n_2_369), .A2(n_485), .B1(n_2_265_2), .B2(n_484), 
      .ZN(n_2_265_1));
   INV_X1 i_2_265_3 (.A(n_2_369), .ZN(n_2_265_2));
   INV_X1 i_2_265_4 (.A(in_data[8]), .ZN(n_2_265_3));
   OAI21_X1 i_2_266_0 (.A(n_2_266_0), .B1(n_2_266_3), .B2(n_2_266_1), .ZN(
      n_2_215));
   NAND2_X1 i_2_266_1 (.A1(n_26), .A2(n_2_266_1), .ZN(n_2_266_0));
   OAI22_X1 i_2_266_2 (.A1(n_2_369), .A2(n_480), .B1(n_2_266_2), .B2(n_479), 
      .ZN(n_2_266_1));
   INV_X1 i_2_266_3 (.A(n_2_369), .ZN(n_2_266_2));
   INV_X1 i_2_266_4 (.A(in_data[8]), .ZN(n_2_266_3));
   OAI21_X1 i_2_267_0 (.A(n_2_267_0), .B1(n_2_267_3), .B2(n_2_267_1), .ZN(
      n_2_216));
   NAND2_X1 i_2_267_1 (.A1(n_25), .A2(n_2_267_1), .ZN(n_2_267_0));
   OAI22_X1 i_2_267_2 (.A1(n_2_369), .A2(n_476), .B1(n_2_267_2), .B2(n_475), 
      .ZN(n_2_267_1));
   INV_X1 i_2_267_3 (.A(n_2_369), .ZN(n_2_267_2));
   INV_X1 i_2_267_4 (.A(in_data[8]), .ZN(n_2_267_3));
   OAI21_X1 i_2_268_0 (.A(n_2_268_0), .B1(n_2_268_3), .B2(n_2_268_1), .ZN(
      n_2_217));
   NAND2_X1 i_2_268_1 (.A1(n_24), .A2(n_2_268_1), .ZN(n_2_268_0));
   OAI22_X1 i_2_268_2 (.A1(n_2_369), .A2(n_472), .B1(n_2_268_2), .B2(n_471), 
      .ZN(n_2_268_1));
   INV_X1 i_2_268_3 (.A(n_2_369), .ZN(n_2_268_2));
   INV_X1 i_2_268_4 (.A(in_data[8]), .ZN(n_2_268_3));
   OAI21_X1 i_2_269_0 (.A(n_2_269_0), .B1(n_2_269_3), .B2(n_2_269_1), .ZN(n_1193));
   NAND2_X1 i_2_269_1 (.A1(n_23), .A2(n_2_269_1), .ZN(n_2_269_0));
   OAI22_X1 i_2_269_2 (.A1(n_2_369), .A2(n_468), .B1(n_2_269_2), .B2(n_467), 
      .ZN(n_2_269_1));
   INV_X1 i_2_269_3 (.A(n_2_369), .ZN(n_2_269_2));
   INV_X1 i_2_269_4 (.A(in_data[8]), .ZN(n_2_269_3));
   OAI21_X1 i_2_270_0 (.A(n_2_270_0), .B1(n_2_270_3), .B2(n_2_270_1), .ZN(
      n_2_218));
   NAND2_X1 i_2_270_1 (.A1(n_22), .A2(n_2_270_1), .ZN(n_2_270_0));
   OAI22_X1 i_2_270_2 (.A1(n_2_369), .A2(n_394), .B1(n_2_270_2), .B2(n_393), 
      .ZN(n_2_270_1));
   INV_X1 i_2_270_3 (.A(n_2_369), .ZN(n_2_270_2));
   INV_X1 i_2_270_4 (.A(in_data[8]), .ZN(n_2_270_3));
   OAI21_X1 i_2_271_0 (.A(n_2_271_0), .B1(n_2_271_3), .B2(n_2_271_1), .ZN(n_1194));
   NAND2_X1 i_2_271_1 (.A1(n_21), .A2(n_2_271_1), .ZN(n_2_271_0));
   OAI22_X1 i_2_271_2 (.A1(n_2_369), .A2(n_389), .B1(n_2_271_2), .B2(n_388), 
      .ZN(n_2_271_1));
   INV_X1 i_2_271_3 (.A(n_2_369), .ZN(n_2_271_2));
   INV_X1 i_2_271_4 (.A(in_data[8]), .ZN(n_2_271_3));
   OAI21_X1 i_2_272_0 (.A(n_2_272_0), .B1(n_2_272_3), .B2(n_2_272_1), .ZN(
      n_2_219));
   NAND2_X1 i_2_272_1 (.A1(n_20), .A2(n_2_272_1), .ZN(n_2_272_0));
   OAI22_X1 i_2_272_2 (.A1(n_2_369), .A2(n_373), .B1(n_2_272_2), .B2(n_372), 
      .ZN(n_2_272_1));
   INV_X1 i_2_272_3 (.A(n_2_369), .ZN(n_2_272_2));
   INV_X1 i_2_272_4 (.A(in_data[8]), .ZN(n_2_272_3));
   OAI21_X1 i_2_273_0 (.A(n_2_273_0), .B1(n_2_273_3), .B2(n_2_273_1), .ZN(
      n_2_220));
   NAND2_X1 i_2_273_1 (.A1(n_19), .A2(n_2_273_1), .ZN(n_2_273_0));
   OAI22_X1 i_2_273_2 (.A1(n_2_369), .A2(n_337), .B1(n_2_273_2), .B2(n_336), 
      .ZN(n_2_273_1));
   INV_X1 i_2_273_3 (.A(n_2_369), .ZN(n_2_273_2));
   INV_X1 i_2_273_4 (.A(in_data[8]), .ZN(n_2_273_3));
   OAI21_X1 i_2_274_0 (.A(n_2_274_0), .B1(n_2_274_3), .B2(n_2_274_1), .ZN(
      n_2_221));
   NAND2_X1 i_2_274_1 (.A1(n_18), .A2(n_2_274_1), .ZN(n_2_274_0));
   OAI22_X1 i_2_274_2 (.A1(n_2_369), .A2(n_285), .B1(n_2_274_2), .B2(n_284), 
      .ZN(n_2_274_1));
   INV_X1 i_2_274_3 (.A(n_2_369), .ZN(n_2_274_2));
   INV_X1 i_2_274_4 (.A(in_data[8]), .ZN(n_2_274_3));
   OAI21_X1 i_2_275_0 (.A(n_2_275_0), .B1(n_2_275_3), .B2(n_2_275_1), .ZN(n_1195));
   NAND2_X1 i_2_275_1 (.A1(n_17), .A2(n_2_275_1), .ZN(n_2_275_0));
   OAI22_X1 i_2_275_2 (.A1(n_2_369), .A2(n_280), .B1(n_2_275_2), .B2(n_279), 
      .ZN(n_2_275_1));
   INV_X1 i_2_275_3 (.A(n_2_369), .ZN(n_2_275_2));
   INV_X1 i_2_275_4 (.A(in_data[8]), .ZN(n_2_275_3));
   OAI21_X1 i_2_276_0 (.A(n_2_276_0), .B1(n_2_276_3), .B2(n_2_276_1), .ZN(
      n_2_222));
   NAND2_X1 i_2_276_1 (.A1(n_16), .A2(n_2_276_1), .ZN(n_2_276_0));
   OAI22_X1 i_2_276_2 (.A1(n_2_369), .A2(n_274), .B1(n_2_276_2), .B2(n_273), 
      .ZN(n_2_276_1));
   INV_X1 i_2_276_3 (.A(n_2_369), .ZN(n_2_276_2));
   INV_X1 i_2_276_4 (.A(in_data[8]), .ZN(n_2_276_3));
   OAI21_X1 i_2_277_0 (.A(n_2_277_0), .B1(n_2_277_3), .B2(n_2_277_1), .ZN(n_1196));
   NAND2_X1 i_2_277_1 (.A1(n_15), .A2(n_2_277_1), .ZN(n_2_277_0));
   OAI22_X1 i_2_277_2 (.A1(n_2_369), .A2(n_264), .B1(n_2_277_2), .B2(n_263), 
      .ZN(n_2_277_1));
   INV_X1 i_2_277_3 (.A(n_2_369), .ZN(n_2_277_2));
   INV_X1 i_2_277_4 (.A(in_data[8]), .ZN(n_2_277_3));
   OAI21_X1 i_2_278_0 (.A(n_2_278_0), .B1(n_2_278_3), .B2(n_2_278_1), .ZN(
      n_2_223));
   NAND2_X1 i_2_278_1 (.A1(n_13), .A2(n_2_278_1), .ZN(n_2_278_0));
   OAI22_X1 i_2_278_2 (.A1(n_2_369), .A2(n_253), .B1(n_2_278_2), .B2(n_252), 
      .ZN(n_2_278_1));
   INV_X1 i_2_278_3 (.A(n_2_369), .ZN(n_2_278_2));
   INV_X1 i_2_278_4 (.A(in_data[8]), .ZN(n_2_278_3));
   OAI21_X1 i_2_279_0 (.A(n_2_279_0), .B1(n_2_279_3), .B2(n_2_279_1), .ZN(
      n_2_224));
   NAND2_X1 i_2_279_1 (.A1(n_12), .A2(n_2_279_1), .ZN(n_2_279_0));
   OAI22_X1 i_2_279_2 (.A1(n_2_369), .A2(n_245), .B1(n_2_279_2), .B2(n_244), 
      .ZN(n_2_279_1));
   INV_X1 i_2_279_3 (.A(n_2_369), .ZN(n_2_279_2));
   INV_X1 i_2_279_4 (.A(in_data[8]), .ZN(n_2_279_3));
   OAI21_X1 i_2_280_0 (.A(n_2_280_0), .B1(n_2_280_3), .B2(n_2_280_1), .ZN(n_1197));
   NAND2_X1 i_2_280_1 (.A1(n_5), .A2(n_2_280_1), .ZN(n_2_280_0));
   OAI22_X1 i_2_280_2 (.A1(n_2_369), .A2(n_151), .B1(n_2_280_2), .B2(n_150), 
      .ZN(n_2_280_1));
   INV_X1 i_2_280_3 (.A(n_2_369), .ZN(n_2_280_2));
   INV_X1 i_2_280_4 (.A(in_data[8]), .ZN(n_2_280_3));
   OAI21_X1 i_2_281_0 (.A(n_2_281_0), .B1(n_2_281_3), .B2(n_2_281_1), .ZN(n_1198));
   NAND2_X1 i_2_281_1 (.A1(n_4), .A2(n_2_281_1), .ZN(n_2_281_0));
   OAI22_X1 i_2_281_2 (.A1(n_2_369), .A2(n_148), .B1(n_2_281_2), .B2(n_147), 
      .ZN(n_2_281_1));
   INV_X1 i_2_281_3 (.A(n_2_369), .ZN(n_2_281_2));
   INV_X1 i_2_281_4 (.A(in_data[8]), .ZN(n_2_281_3));
   AND2_X1 i_2_282_0 (.A1(n_659), .A2(n_2_229), .ZN(n_2_2));
   OR2_X1 i_2_283_0 (.A1(n_2_229), .A2(n_659), .ZN(n_2_3));
   AND2_X1 i_2_284_0 (.A1(n_660), .A2(n_2_230), .ZN(n_1199));
   OR2_X1 i_2_285_0 (.A1(n_2_230), .A2(n_660), .ZN(n_1200));
   AND2_X1 i_2_286_0 (.A1(n_652), .A2(n_2_231), .ZN(n_2_6));
   OR2_X1 i_2_287_0 (.A1(n_2_231), .A2(n_652), .ZN(n_2_7));
   AND2_X1 i_2_288_0 (.A1(n_628), .A2(n_2_238), .ZN(n_2_18));
   OR2_X1 i_2_289_0 (.A1(n_2_238), .A2(n_628), .ZN(n_2_19));
   AND2_X1 i_2_290_0 (.A1(n_620), .A2(n_2_242), .ZN(n_1201));
   OR2_X1 i_2_291_0 (.A1(n_2_242), .A2(n_620), .ZN(n_1202));
   AND2_X1 i_2_292_0 (.A1(n_616), .A2(n_2_243), .ZN(n_2_23));
   OR2_X1 i_2_293_0 (.A1(n_2_243), .A2(n_616), .ZN(n_2_24));
   AND2_X1 i_2_294_0 (.A1(n_601), .A2(n_2_249), .ZN(n_2_29));
   OR2_X1 i_2_295_0 (.A1(n_2_249), .A2(n_601), .ZN(n_2_30));
   AND2_X1 i_2_296_0 (.A1(n_586), .A2(n_2_252), .ZN(n_2_39));
   OR2_X1 i_2_297_0 (.A1(n_2_252), .A2(n_586), .ZN(n_2_40));
   AND2_X1 i_2_298_0 (.A1(n_570), .A2(n_2_256), .ZN(n_2_51));
   OR2_X1 i_2_299_0 (.A1(n_2_256), .A2(n_570), .ZN(n_2_52));
   AND2_X1 i_2_300_0 (.A1(n_566), .A2(n_2_257), .ZN(n_2_54));
   OR2_X1 i_2_301_0 (.A1(n_2_257), .A2(n_566), .ZN(n_2_55));
   AND2_X1 i_2_302_0 (.A1(n_562), .A2(n_2_258), .ZN(n_2_57));
   OR2_X1 i_2_303_0 (.A1(n_2_258), .A2(n_562), .ZN(n_2_58));
   AND2_X1 i_2_304_0 (.A1(n_554), .A2(n_2_260), .ZN(n_2_61));
   OR2_X1 i_2_305_0 (.A1(n_2_260), .A2(n_554), .ZN(n_2_62));
   AND2_X1 i_2_306_0 (.A1(n_478), .A2(n_2_264), .ZN(n_2_81));
   OR2_X1 i_2_307_0 (.A1(n_2_264), .A2(n_478), .ZN(n_2_82));
   AND2_X1 i_2_308_0 (.A1(n_474), .A2(n_2_265), .ZN(n_2_84));
   OR2_X1 i_2_309_0 (.A1(n_2_265), .A2(n_474), .ZN(n_2_85));
   AND2_X1 i_2_310_0 (.A1(n_470), .A2(n_2_266), .ZN(n_2_87));
   OR2_X1 i_2_311_0 (.A1(n_2_266), .A2(n_470), .ZN(n_2_88));
   AND2_X1 i_2_312_0 (.A1(n_466), .A2(n_1270), .ZN(n_1203));
   AND2_X1 i_2_313_0 (.A1(n_441), .A2(n_1271), .ZN(n_2_95));
   AND2_X1 i_2_314_0 (.A1(n_431), .A2(n_2_267), .ZN(n_2_98));
   OR2_X1 i_2_315_0 (.A1(n_2_267), .A2(n_431), .ZN(n_2_99));
   AND2_X1 i_2_316_0 (.A1(n_769), .A2(n_2_269), .ZN(n_2_114));
   OR2_X1 i_2_317_0 (.A1(n_2_269), .A2(n_769), .ZN(n_2_115));
   AND2_X1 i_2_318_0 (.A1(n_768), .A2(n_2_270), .ZN(n_2_117));
   OR2_X1 i_2_319_0 (.A1(n_2_270), .A2(n_768), .ZN(n_2_118));
   AND2_X1 i_2_320_0 (.A1(n_767), .A2(n_2_271), .ZN(n_2_124));
   OR2_X1 i_2_321_0 (.A1(n_2_271), .A2(n_767), .ZN(n_2_125));
   AND2_X1 i_2_322_0 (.A1(n_766), .A2(n_2_272), .ZN(n_2_130));
   OR2_X1 i_2_323_0 (.A1(n_2_272), .A2(n_766), .ZN(n_2_131));
   AND2_X1 i_2_324_0 (.A1(n_760), .A2(n_2_278), .ZN(n_2_151));
   OR2_X1 i_2_325_0 (.A1(n_2_278), .A2(n_760), .ZN(n_2_152));
   AND2_X1 i_2_326_0 (.A1(n_759), .A2(n_2_279), .ZN(n_2_154));
   OR2_X1 i_2_327_0 (.A1(n_2_279), .A2(n_759), .ZN(n_2_155));
   AND2_X1 i_2_328_0 (.A1(n_758), .A2(n_2_280), .ZN(n_2_158));
   OR2_X1 i_2_329_0 (.A1(n_2_280), .A2(n_758), .ZN(n_2_159));
   AND2_X1 i_2_330_0 (.A1(n_757), .A2(n_2_281), .ZN(n_1204));
   OR2_X1 i_2_331_0 (.A1(n_2_281), .A2(n_757), .ZN(n_1205));
   AND2_X1 i_2_332_0 (.A1(n_755), .A2(n_2_283), .ZN(n_2_169));
   OR2_X1 i_2_333_0 (.A1(n_2_283), .A2(n_755), .ZN(n_2_170));
   AND2_X1 i_2_334_0 (.A1(n_753), .A2(n_2_285), .ZN(n_2_181));
   OR2_X1 i_2_335_0 (.A1(n_2_285), .A2(n_753), .ZN(n_2_182));
   AND2_X1 i_2_336_0 (.A1(n_752), .A2(n_2_286), .ZN(n_1206));
   OR2_X1 i_2_337_0 (.A1(n_2_286), .A2(n_752), .ZN(n_1207));
   AND2_X1 i_2_338_0 (.A1(n_751), .A2(n_2_287), .ZN(n_2_186));
   OR2_X1 i_2_339_0 (.A1(n_2_287), .A2(n_751), .ZN(n_2_187));
   AND2_X1 i_2_340_0 (.A1(n_750), .A2(n_2_288), .ZN(n_2_189));
   OR2_X1 i_2_341_0 (.A1(n_2_288), .A2(n_750), .ZN(n_2_190));
   AND2_X1 i_2_342_0 (.A1(n_749), .A2(n_2_289), .ZN(n_2_199));
   OR2_X1 i_2_343_0 (.A1(n_2_289), .A2(n_749), .ZN(n_2_200));
   AND2_X1 i_2_344_0 (.A1(n_748), .A2(n_2_290), .ZN(n_1208));
   OR2_X1 i_2_345_0 (.A1(n_2_290), .A2(n_748), .ZN(n_1209));
   AND2_X1 i_2_346_0 (.A1(n_747), .A2(n_2_291), .ZN(n_1210));
   OR2_X1 i_2_347_0 (.A1(n_2_291), .A2(n_747), .ZN(n_1211));
   OR2_X1 i_2_348_0 (.A1(n_1272), .A2(n_746), .ZN(n_2_206));
   OAI21_X1 i_2_349_0 (.A(n_2_349_0), .B1(n_2_369), .B2(n_2_349_1), .ZN(n_2_8));
   AOI21_X1 i_2_349_1 (.A(n_651), .B1(n_2_369), .B2(n_649), .ZN(n_2_349_0));
   INV_X1 i_2_349_2 (.A(n_650), .ZN(n_2_349_1));
   OAI21_X1 i_2_350_0 (.A(n_2_350_0), .B1(n_2_369), .B2(n_2_350_1), .ZN(n_2_16));
   AOI21_X1 i_2_350_1 (.A(n_635), .B1(n_2_369), .B2(n_633), .ZN(n_2_350_0));
   INV_X1 i_2_350_2 (.A(n_634), .ZN(n_2_350_1));
   OAI21_X1 i_2_351_0 (.A(n_2_351_0), .B1(n_2_369), .B2(n_2_351_1), .ZN(n_2_20));
   AOI21_X1 i_2_351_1 (.A(n_627), .B1(n_2_369), .B2(n_625), .ZN(n_2_351_0));
   INV_X1 i_2_351_2 (.A(n_626), .ZN(n_2_351_1));
   OAI21_X1 i_2_352_0 (.A(n_2_352_0), .B1(n_2_369), .B2(n_2_352_1), .ZN(n_2_26));
   AOI21_X1 i_2_352_1 (.A(n_611), .B1(n_2_369), .B2(n_609), .ZN(n_2_352_0));
   INV_X1 i_2_352_2 (.A(n_610), .ZN(n_2_352_1));
   OAI21_X1 i_2_353_0 (.A(n_2_353_0), .B1(n_2_369), .B2(n_2_353_1), .ZN(n_2_27));
   AOI21_X1 i_2_353_1 (.A(n_608), .B1(n_2_369), .B2(n_606), .ZN(n_2_353_0));
   INV_X1 i_2_353_2 (.A(n_607), .ZN(n_2_353_1));
   OAI21_X1 i_2_354_0 (.A(n_2_354_0), .B1(n_2_369), .B2(n_2_354_1), .ZN(n_2_59));
   AOI21_X1 i_2_354_1 (.A(n_561), .B1(n_2_369), .B2(n_559), .ZN(n_2_354_0));
   INV_X1 i_2_354_2 (.A(n_560), .ZN(n_2_354_1));
   OAI21_X1 i_2_355_0 (.A(n_2_355_0), .B1(n_2_369), .B2(n_2_355_1), .ZN(n_2_63));
   AOI21_X1 i_2_355_1 (.A(n_553), .B1(n_2_369), .B2(n_551), .ZN(n_2_355_0));
   INV_X1 i_2_355_2 (.A(n_552), .ZN(n_2_355_1));
   OAI21_X1 i_2_356_0 (.A(n_2_356_0), .B1(n_2_369), .B2(n_2_356_1), .ZN(n_2_74));
   AOI21_X1 i_2_356_1 (.A(n_511), .B1(n_2_369), .B2(n_509), .ZN(n_2_356_0));
   INV_X1 i_2_356_2 (.A(n_510), .ZN(n_2_356_1));
   OAI21_X1 i_2_357_0 (.A(n_2_357_0), .B1(n_2_369), .B2(n_2_357_1), .ZN(n_2_108));
   AOI21_X1 i_2_357_1 (.A(n_390), .B1(n_2_369), .B2(n_388), .ZN(n_2_357_0));
   INV_X1 i_2_357_2 (.A(n_389), .ZN(n_2_357_1));
   OAI21_X1 i_2_358_0 (.A(n_2_358_0), .B1(n_2_369), .B2(n_2_358_1), .ZN(n_2_109));
   AOI21_X1 i_2_358_1 (.A(n_385), .B1(n_2_369), .B2(n_383), .ZN(n_2_358_0));
   INV_X1 i_2_358_2 (.A(n_384), .ZN(n_2_358_1));
   OAI21_X1 i_2_359_0 (.A(n_2_359_0), .B1(n_2_369), .B2(n_2_359_1), .ZN(n_2_164));
   AOI21_X1 i_2_359_1 (.A(n_265), .B1(n_2_369), .B2(n_263), .ZN(n_2_359_0));
   INV_X1 i_2_359_2 (.A(n_264), .ZN(n_2_359_1));
   OAI21_X1 i_2_360_0 (.A(n_2_360_0), .B1(n_2_360_1), .B2(n_2_241), .ZN(n_1212));
   NAND2_X1 i_2_360_1 (.A1(n_2_241), .A2(in_data[0]), .ZN(n_2_360_0));
   INV_X1 i_2_360_2 (.A(n_974), .ZN(n_2_360_1));
   OAI21_X1 i_2_361_0 (.A(n_2_361_0), .B1(n_2_339), .B2(n_2_361_1), .ZN(n_2_204));
   AOI21_X1 i_2_361_1 (.A(n_146), .B1(n_2_339), .B2(n_144), .ZN(n_2_361_0));
   INV_X1 i_2_361_2 (.A(n_145), .ZN(n_2_361_1));
   OAI21_X1 i_2_362_0 (.A(n_2_362_0), .B1(n_2_339), .B2(n_2_362_1), .ZN(n_2_195));
   AOI21_X1 i_2_362_1 (.A(n_178), .B1(n_2_339), .B2(n_176), .ZN(n_2_362_0));
   INV_X1 i_2_362_2 (.A(n_177), .ZN(n_2_362_1));
   OAI21_X1 i_2_363_0 (.A(n_2_363_0), .B1(n_2_339), .B2(n_2_363_1), .ZN(n_2_193));
   AOI21_X1 i_2_363_1 (.A(n_188), .B1(n_2_339), .B2(n_186), .ZN(n_2_363_0));
   INV_X1 i_2_363_2 (.A(n_187), .ZN(n_2_363_1));
   OAI21_X1 i_2_364_0 (.A(n_2_364_0), .B1(n_2_339), .B2(n_2_364_1), .ZN(n_2_178));
   AOI21_X1 i_2_364_1 (.A(n_225), .B1(n_2_339), .B2(n_223), .ZN(n_2_364_0));
   INV_X1 i_2_364_2 (.A(n_224), .ZN(n_2_364_1));
   OAI21_X1 i_2_365_0 (.A(n_2_365_0), .B1(n_2_339), .B2(n_2_365_1), .ZN(n_2_175));
   AOI21_X1 i_2_365_1 (.A(n_231), .B1(n_2_339), .B2(n_229), .ZN(n_2_365_0));
   INV_X1 i_2_365_2 (.A(n_230), .ZN(n_2_365_1));
   OAI21_X1 i_2_366_0 (.A(n_2_366_0), .B1(n_2_339), .B2(n_2_366_1), .ZN(n_2_171));
   AOI21_X1 i_2_366_1 (.A(n_251), .B1(n_2_339), .B2(n_249), .ZN(n_2_366_0));
   INV_X1 i_2_366_2 (.A(n_250), .ZN(n_2_366_1));
   OAI21_X1 i_2_367_0 (.A(n_2_367_0), .B1(n_2_339), .B2(n_2_367_1), .ZN(n_2_147));
   AOI21_X1 i_2_367_1 (.A(n_303), .B1(n_2_339), .B2(n_301), .ZN(n_2_367_0));
   INV_X1 i_2_367_2 (.A(n_302), .ZN(n_2_367_1));
   OAI21_X1 i_2_368_0 (.A(n_2_368_0), .B1(n_2_339), .B2(n_2_368_1), .ZN(n_2_143));
   AOI21_X1 i_2_368_1 (.A(n_311), .B1(n_2_339), .B2(n_309), .ZN(n_2_368_0));
   INV_X1 i_2_368_2 (.A(n_310), .ZN(n_2_368_1));
   OAI21_X1 i_2_369_0 (.A(n_2_369_0), .B1(n_2_339), .B2(n_2_369_1), .ZN(n_2_139));
   AOI21_X1 i_2_369_1 (.A(n_319), .B1(n_2_339), .B2(n_317), .ZN(n_2_369_0));
   INV_X1 i_2_369_2 (.A(n_318), .ZN(n_2_369_1));
   OAI21_X1 i_2_370_0 (.A(n_2_370_0), .B1(n_2_339), .B2(n_2_370_1), .ZN(n_2_135));
   AOI21_X1 i_2_370_1 (.A(n_327), .B1(n_2_339), .B2(n_325), .ZN(n_2_370_0));
   INV_X1 i_2_370_2 (.A(n_326), .ZN(n_2_370_1));
   OAI21_X1 i_2_371_0 (.A(n_2_371_0), .B1(n_2_339), .B2(n_2_371_1), .ZN(n_2_132));
   AOI21_X1 i_2_371_1 (.A(n_330), .B1(n_2_339), .B2(n_328), .ZN(n_2_371_0));
   INV_X1 i_2_371_2 (.A(n_329), .ZN(n_2_371_1));
   OAI21_X1 i_2_372_0 (.A(n_2_372_0), .B1(n_2_339), .B2(n_2_372_1), .ZN(n_2_107));
   AOI21_X1 i_2_372_1 (.A(n_395), .B1(n_2_339), .B2(n_393), .ZN(n_2_372_0));
   INV_X1 i_2_372_2 (.A(n_394), .ZN(n_2_372_1));
   OAI21_X1 i_2_373_0 (.A(n_2_373_0), .B1(n_2_339), .B2(n_2_373_1), .ZN(n_2_105));
   AOI21_X1 i_2_373_1 (.A(n_405), .B1(n_2_339), .B2(n_403), .ZN(n_2_373_0));
   INV_X1 i_2_373_2 (.A(n_404), .ZN(n_2_373_1));
   OAI21_X1 i_2_374_0 (.A(n_2_374_0), .B1(n_2_339), .B2(n_2_374_1), .ZN(n_2_103));
   AOI21_X1 i_2_374_1 (.A(n_415), .B1(n_2_339), .B2(n_413), .ZN(n_2_374_0));
   INV_X1 i_2_374_2 (.A(n_414), .ZN(n_2_374_1));
   OAI21_X1 i_2_375_0 (.A(n_2_375_0), .B1(n_2_339), .B2(n_2_375_1), .ZN(n_2_101));
   AOI21_X1 i_2_375_1 (.A(n_425), .B1(n_2_339), .B2(n_423), .ZN(n_2_375_0));
   INV_X1 i_2_375_2 (.A(n_424), .ZN(n_2_375_1));
   OAI21_X1 i_2_376_0 (.A(n_2_376_0), .B1(n_2_339), .B2(n_2_376_1), .ZN(n_2_96));
   AOI21_X1 i_2_376_1 (.A(n_439), .B1(n_2_339), .B2(n_437), .ZN(n_2_376_0));
   INV_X1 i_2_376_2 (.A(n_438), .ZN(n_2_376_1));
   OAI21_X1 i_2_377_0 (.A(n_2_377_0), .B1(n_2_339), .B2(n_2_377_1), .ZN(n_2_92));
   AOI21_X1 i_2_377_1 (.A(n_454), .B1(n_2_339), .B2(n_452), .ZN(n_2_377_0));
   INV_X1 i_2_377_2 (.A(n_453), .ZN(n_2_377_1));
   OAI21_X1 i_2_378_0 (.A(n_2_378_0), .B1(n_2_339), .B2(n_2_378_1), .ZN(n_2_79));
   AOI21_X1 i_2_378_1 (.A(n_486), .B1(n_2_339), .B2(n_484), .ZN(n_2_378_0));
   INV_X1 i_2_378_2 (.A(n_485), .ZN(n_2_378_1));
   OAI21_X1 i_2_379_0 (.A(n_2_379_0), .B1(n_2_339), .B2(n_2_379_1), .ZN(n_2_73));
   AOI21_X1 i_2_379_1 (.A(n_516), .B1(n_2_339), .B2(n_514), .ZN(n_2_379_0));
   INV_X1 i_2_379_2 (.A(n_515), .ZN(n_2_379_1));
   OAI21_X1 i_2_380_0 (.A(n_2_380_0), .B1(n_2_339), .B2(n_2_380_1), .ZN(n_2_72));
   AOI21_X1 i_2_380_1 (.A(n_521), .B1(n_2_339), .B2(n_519), .ZN(n_2_380_0));
   INV_X1 i_2_380_2 (.A(n_520), .ZN(n_2_380_1));
   OAI21_X1 i_2_381_0 (.A(n_2_381_0), .B1(n_2_339), .B2(n_2_381_1), .ZN(n_2_44));
   AOI21_X1 i_2_381_1 (.A(n_581), .B1(n_2_339), .B2(n_579), .ZN(n_2_381_0));
   INV_X1 i_2_381_2 (.A(n_580), .ZN(n_2_381_1));
   OAI21_X1 i_2_382_0 (.A(n_2_382_0), .B1(n_2_339), .B2(n_2_382_1), .ZN(n_2_35));
   AOI21_X1 i_2_382_1 (.A(n_591), .B1(n_2_339), .B2(n_589), .ZN(n_2_382_0));
   INV_X1 i_2_382_2 (.A(n_590), .ZN(n_2_382_1));
   OAI21_X1 i_2_383_0 (.A(n_2_383_0), .B1(n_2_339), .B2(n_2_383_1), .ZN(n_2_9));
   AOI21_X1 i_2_383_1 (.A(n_647), .B1(n_2_339), .B2(n_645), .ZN(n_2_383_0));
   INV_X1 i_2_383_2 (.A(n_646), .ZN(n_2_383_1));
   OAI21_X1 i_2_384_0 (.A(n_2_384_0), .B1(n_2_339), .B2(n_2_384_1), .ZN(n_2_146));
   AOI21_X1 i_2_384_1 (.A(n_308), .B1(n_2_339), .B2(n_306), .ZN(n_2_384_0));
   INV_X1 i_2_384_2 (.A(n_307), .ZN(n_2_384_1));
   OAI21_X1 i_2_385_0 (.A(n_2_385_0), .B1(n_2_339), .B2(n_2_385_1), .ZN(n_2_64));
   AOI21_X1 i_2_385_1 (.A(n_549), .B1(n_2_339), .B2(n_547), .ZN(n_2_385_0));
   INV_X1 i_2_385_2 (.A(n_548), .ZN(n_2_385_1));
   OAI21_X1 i_2_386_0 (.A(n_2_386_0), .B1(n_2_339), .B2(n_2_386_1), .ZN(n_2_47));
   AOI21_X1 i_2_386_1 (.A(n_577), .B1(n_2_339), .B2(n_575), .ZN(n_2_386_0));
   INV_X1 i_2_386_2 (.A(n_576), .ZN(n_2_386_1));
   OAI21_X1 i_2_387_0 (.A(n_2_387_0), .B1(n_2_339), .B2(n_2_387_1), .ZN(n_2_41));
   AOI21_X1 i_2_387_1 (.A(n_585), .B1(n_2_339), .B2(n_583), .ZN(n_2_387_0));
   INV_X1 i_2_387_2 (.A(n_584), .ZN(n_2_387_1));
   OAI21_X1 i_2_388_0 (.A(n_2_388_0), .B1(n_2_339), .B2(n_2_388_1), .ZN(n_2_32));
   AOI21_X1 i_2_388_1 (.A(n_595), .B1(n_2_339), .B2(n_593), .ZN(n_2_388_0));
   INV_X1 i_2_388_2 (.A(n_594), .ZN(n_2_388_1));
   OAI21_X1 i_2_389_0 (.A(n_2_389_0), .B1(n_2_339), .B2(n_2_389_1), .ZN(n_2_31));
   AOI21_X1 i_2_389_1 (.A(n_600), .B1(n_2_339), .B2(n_598), .ZN(n_2_389_0));
   INV_X1 i_2_389_2 (.A(n_599), .ZN(n_2_389_1));
   OAI21_X1 i_2_390_0 (.A(n_2_390_0), .B1(n_2_339), .B2(n_2_390_1), .ZN(n_2_25));
   AOI21_X1 i_2_390_1 (.A(n_615), .B1(n_2_339), .B2(n_613), .ZN(n_2_390_0));
   INV_X1 i_2_390_2 (.A(n_614), .ZN(n_2_390_1));
   OAI21_X1 i_2_391_0 (.A(n_2_391_0), .B1(n_2_339), .B2(n_2_391_1), .ZN(n_2_192));
   AOI21_X1 i_2_391_1 (.A(n_193), .B1(n_2_339), .B2(n_191), .ZN(n_2_391_0));
   INV_X1 i_2_391_2 (.A(n_192), .ZN(n_2_391_1));
   OAI21_X1 i_2_392_0 (.A(n_2_392_0), .B1(n_2_339), .B2(n_2_392_1), .ZN(n_2_191));
   AOI21_X1 i_2_392_1 (.A(n_198), .B1(n_2_339), .B2(n_196), .ZN(n_2_392_0));
   INV_X1 i_2_392_2 (.A(n_197), .ZN(n_2_392_1));
   OAI21_X1 i_2_393_0 (.A(n_2_393_0), .B1(n_2_339), .B2(n_2_393_1), .ZN(n_2_183));
   AOI21_X1 i_2_393_1 (.A(n_212), .B1(n_2_339), .B2(n_210), .ZN(n_2_393_0));
   INV_X1 i_2_393_2 (.A(n_211), .ZN(n_2_393_1));
   OAI21_X1 i_2_394_0 (.A(n_2_394_0), .B1(n_2_339), .B2(n_2_394_1), .ZN(n_2_106));
   AOI21_X1 i_2_394_1 (.A(n_400), .B1(n_2_339), .B2(n_398), .ZN(n_2_394_0));
   INV_X1 i_2_394_2 (.A(n_399), .ZN(n_2_394_1));
   OAI21_X1 i_2_395_0 (.A(n_2_395_0), .B1(n_2_339), .B2(n_2_395_1), .ZN(n_2_13));
   AOI21_X1 i_2_395_1 (.A(n_639), .B1(n_2_339), .B2(n_637), .ZN(n_2_395_0));
   INV_X1 i_2_395_2 (.A(n_638), .ZN(n_2_395_1));
   OAI21_X1 i_2_396_0 (.A(n_2_396_0), .B1(n_2_339), .B2(n_2_396_1), .ZN(n_2_10));
   AOI21_X1 i_2_396_1 (.A(n_642), .B1(n_2_339), .B2(n_640), .ZN(n_2_396_0));
   INV_X1 i_2_396_2 (.A(n_641), .ZN(n_2_396_1));
   OAI21_X1 i_2_397_0 (.A(n_2_397_0), .B1(n_2_339), .B2(n_2_397_1), .ZN(n_2_207));
   AOI21_X1 i_2_397_1 (.A(n_137), .B1(n_2_339), .B2(n_135), .ZN(n_2_397_0));
   INV_X1 i_2_397_2 (.A(n_136), .ZN(n_2_397_1));
   OAI21_X1 i_2_398_0 (.A(n_2_398_0), .B1(n_2_339), .B2(n_2_398_1), .ZN(n_2_179));
   AOI21_X1 i_2_398_1 (.A(n_220), .B1(n_2_339), .B2(n_218), .ZN(n_2_398_0));
   INV_X1 i_2_398_2 (.A(n_219), .ZN(n_2_398_1));
   CLKGATETST_X1 clk_gate_buf_fill_i_reg (.CK(clk), .E(enbl_in), .SE(1'b0), 
      .GCK(n_2_298));
   range_extractor__3_149 range_extr_0 (.in_a(buf_fill_i), .in_size({in_data[31], 
      in_data[30], in_data[29]}), .out_a(\out_as[0] ), .out_b({n_2_345, n_2_344, 
      n_2_343, n_2_342, n_2_341, n_2_340, n_2_360}));
   range_extractor__3_201 ranges_1_range_extr_i (.in_a({n_2_345, n_2_344, 
      n_2_343, n_2_342, n_2_341, n_2_340, n_2_360}), .in_size({in_data[27], 
      in_data[26], in_data[25]}), .out_a(\out_as[1] ), .out_b({n_2_348, n_2_362, 
      n_2_372, n_2_370, n_2_347, n_2_346, n_2_361}));
   range_extractor__3_253 ranges_2_range_extr_i (.in_a({n_2_348, n_2_362, 
      n_2_372, n_2_370, n_2_347, n_2_346, n_2_361}), .in_size({in_data[23], 
      in_data[22], in_data[21]}), .out_a(\out_as[2] ), .out_b({n_2_354, n_2_353, 
      n_2_352, n_2_351, n_2_350, n_2_349, \out_bs[2] [0]}));
   range_extractor__3_305 ranges_3_range_extr_i (.in_a({n_2_354, n_2_353, 
      n_2_352, n_2_351, n_2_350, n_2_349, \out_bs[2] [0]}), .in_size({
      in_data[19], in_data[18], in_data[17]}), .out_a(\out_as[3] ), .out_b({
      n_2_358, n_2_357, n_2_356, n_2_364, n_2_355, n_2_363, \out_bs[3] [0]}));
   range_extractor__3_357 ranges_4_range_extr_i (.in_a({n_2_358, n_2_357, 
      n_2_356, n_2_364, n_2_355, n_2_363, \out_bs[3] [0]}), .in_size({
      in_data[15], in_data[14], in_data[13]}), .out_a(\out_as[4] ), .out_b({
      n_2_359, \out_bs[4] [5], n_2_367, n_2_366, n_2_365, n_2_299, 
      \out_bs[4] [0]}));
   range_extractor__3_409 ranges_5_range_extr_i (.in_a({n_2_359, \out_bs[4] [5], 
      n_2_367, n_2_366, n_2_365, n_2_299, \out_bs[4] [0]}), .in_size({
      in_data[11], in_data[10], in_data[9]}), .out_a(\out_as[5] ), .out_b(
      \out_bs[5] ));
   OR3_X1 i_2_399_0 (.A1(n_2_399_0), .A2(n_130), .A3(n_131), .ZN(n_1213));
   INV_X1 i_2_399_1 (.A(n_952), .ZN(n_2_399_0));
   NAND2_X1 i_2_400_0 (.A1(n_2_400_3), .A2(n_2_400_0), .ZN(n_1214));
   INV_X1 i_2_400_1 (.A(n_2_400_1), .ZN(n_2_400_0));
   NAND2_X1 i_2_400_2 (.A1(n_952), .A2(n_2_400_2), .ZN(n_2_400_1));
   INV_X1 i_2_400_3 (.A(n_129), .ZN(n_2_400_2));
   INV_X1 i_2_400_4 (.A(n_834), .ZN(n_2_400_3));
   OAI21_X1 i_2_401_0 (.A(n_2_401_0), .B1(n_952), .B2(n_2_401_1), .ZN(n_1215));
   AOI21_X1 i_2_401_1 (.A(n_2_207), .B1(n_952), .B2(n_133), .ZN(n_2_401_0));
   INV_X1 i_2_401_2 (.A(n_134), .ZN(n_2_401_1));
   OAI21_X1 i_2_402_0 (.A(n_2_402_0), .B1(n_952), .B2(n_2_402_1), .ZN(n_1216));
   AOI21_X1 i_2_402_1 (.A(n_2_204), .B1(n_952), .B2(n_142), .ZN(n_2_402_0));
   INV_X1 i_2_402_2 (.A(n_143), .ZN(n_2_402_1));
   OAI21_X1 i_2_403_0 (.A(n_2_403_0), .B1(n_952), .B2(n_2_403_1), .ZN(n_1217));
   AOI21_X1 i_2_403_1 (.A(n_160), .B1(n_952), .B2(n_158), .ZN(n_2_403_0));
   INV_X1 i_2_403_2 (.A(n_159), .ZN(n_2_403_1));
   OAI21_X1 i_2_404_0 (.A(n_2_404_0), .B1(n_952), .B2(n_2_404_1), .ZN(n_1218));
   AOI21_X1 i_2_404_1 (.A(n_2_195), .B1(n_952), .B2(n_174), .ZN(n_2_404_0));
   INV_X1 i_2_404_2 (.A(n_175), .ZN(n_2_404_1));
   OAI21_X1 i_2_405_0 (.A(n_2_405_0), .B1(n_952), .B2(n_2_405_1), .ZN(n_1219));
   AOI21_X1 i_2_405_1 (.A(n_2_193), .B1(n_952), .B2(n_184), .ZN(n_2_405_0));
   INV_X1 i_2_405_2 (.A(n_185), .ZN(n_2_405_1));
   OAI21_X1 i_2_406_0 (.A(n_2_406_0), .B1(n_952), .B2(n_2_406_1), .ZN(n_1220));
   AOI21_X1 i_2_406_1 (.A(n_2_192), .B1(n_952), .B2(n_189), .ZN(n_2_406_0));
   INV_X1 i_2_406_2 (.A(n_190), .ZN(n_2_406_1));
   OAI21_X1 i_2_407_0 (.A(n_2_407_0), .B1(n_952), .B2(n_2_407_1), .ZN(n_1221));
   AOI21_X1 i_2_407_1 (.A(n_2_191), .B1(n_952), .B2(n_194), .ZN(n_2_407_0));
   INV_X1 i_2_407_2 (.A(n_195), .ZN(n_2_407_1));
   OAI21_X1 i_2_408_0 (.A(n_2_408_0), .B1(n_952), .B2(n_2_408_1), .ZN(n_1222));
   AOI21_X1 i_2_408_1 (.A(n_2_183), .B1(n_952), .B2(n_208), .ZN(n_2_408_0));
   INV_X1 i_2_408_2 (.A(n_209), .ZN(n_2_408_1));
   OAI21_X1 i_2_409_0 (.A(n_2_409_0), .B1(n_952), .B2(n_2_409_1), .ZN(n_1223));
   AOI21_X1 i_2_409_1 (.A(n_2_179), .B1(n_952), .B2(n_216), .ZN(n_2_409_0));
   INV_X1 i_2_409_2 (.A(n_217), .ZN(n_2_409_1));
   OAI21_X1 i_2_410_0 (.A(n_2_410_0), .B1(n_952), .B2(n_2_410_1), .ZN(n_1224));
   AOI21_X1 i_2_410_1 (.A(n_2_178), .B1(n_952), .B2(n_221), .ZN(n_2_410_0));
   INV_X1 i_2_410_2 (.A(n_222), .ZN(n_2_410_1));
   OAI21_X1 i_2_411_0 (.A(n_2_411_0), .B1(n_952), .B2(n_2_411_1), .ZN(n_1225));
   AOI21_X1 i_2_411_1 (.A(n_226), .B1(n_952), .B2(n_2_176), .ZN(n_2_411_0));
   INV_X1 i_2_411_2 (.A(n_2_177), .ZN(n_2_411_1));
   OAI21_X1 i_2_412_0 (.A(n_2_412_0), .B1(n_952), .B2(n_2_412_1), .ZN(n_1226));
   AOI21_X1 i_2_412_1 (.A(n_2_175), .B1(n_952), .B2(n_227), .ZN(n_2_412_0));
   INV_X1 i_2_412_2 (.A(n_228), .ZN(n_2_412_1));
   OAI21_X1 i_2_413_0 (.A(n_2_413_0), .B1(n_952), .B2(n_2_413_1), .ZN(n_1227));
   AOI21_X1 i_2_413_1 (.A(n_2_171), .B1(n_952), .B2(n_247), .ZN(n_2_413_0));
   INV_X1 i_2_413_2 (.A(n_248), .ZN(n_2_413_1));
   OAI21_X1 i_2_414_0 (.A(n_2_414_0), .B1(n_952), .B2(n_2_414_1), .ZN(n_1228));
   AOI21_X1 i_2_414_1 (.A(n_260), .B1(n_952), .B2(n_2_165), .ZN(n_2_414_0));
   INV_X1 i_2_414_2 (.A(n_2_166), .ZN(n_2_414_1));
   OAI21_X1 i_2_415_0 (.A(n_2_415_0), .B1(n_952), .B2(n_2_415_1), .ZN(n_1229));
   AOI21_X1 i_2_415_1 (.A(n_2_164), .B1(n_952), .B2(n_261), .ZN(n_2_415_0));
   INV_X1 i_2_415_2 (.A(n_262), .ZN(n_2_415_1));
   OAI21_X1 i_2_416_0 (.A(n_2_416_0), .B1(n_952), .B2(n_2_416_1), .ZN(n_1230));
   AOI21_X1 i_2_416_1 (.A(n_278), .B1(n_952), .B2(n_276), .ZN(n_2_416_0));
   INV_X1 i_2_416_2 (.A(n_277), .ZN(n_2_416_1));
   OAI21_X1 i_2_417_0 (.A(n_2_417_0), .B1(n_952), .B2(n_2_417_1), .ZN(n_1231));
   AOI21_X1 i_2_417_1 (.A(n_2_147), .B1(n_952), .B2(n_2_148), .ZN(n_2_417_0));
   INV_X1 i_2_417_2 (.A(n_2_149), .ZN(n_2_417_1));
   OAI21_X1 i_2_418_0 (.A(n_2_418_0), .B1(n_952), .B2(n_2_418_1), .ZN(n_1232));
   AOI21_X1 i_2_418_1 (.A(n_2_146), .B1(n_952), .B2(n_304), .ZN(n_2_418_0));
   INV_X1 i_2_418_2 (.A(n_305), .ZN(n_2_418_1));
   OAI21_X1 i_2_419_0 (.A(n_2_419_0), .B1(n_952), .B2(n_2_419_1), .ZN(n_1233));
   AOI21_X1 i_2_419_1 (.A(n_2_143), .B1(n_952), .B2(n_2_144), .ZN(n_2_419_0));
   INV_X1 i_2_419_2 (.A(n_2_145), .ZN(n_2_419_1));
   OAI21_X1 i_2_420_0 (.A(n_2_420_0), .B1(n_952), .B2(n_2_420_1), .ZN(n_1234));
   AOI21_X1 i_2_420_1 (.A(n_2_139), .B1(n_952), .B2(n_2_140), .ZN(n_2_420_0));
   INV_X1 i_2_420_2 (.A(n_2_141), .ZN(n_2_420_1));
   OAI21_X1 i_2_421_0 (.A(n_2_421_0), .B1(n_952), .B2(n_2_421_1), .ZN(n_1235));
   AOI21_X1 i_2_421_1 (.A(n_2_135), .B1(n_952), .B2(n_2_136), .ZN(n_2_421_0));
   INV_X1 i_2_421_2 (.A(n_2_137), .ZN(n_2_421_1));
   OAI21_X1 i_2_422_0 (.A(n_2_422_0), .B1(n_952), .B2(n_2_422_1), .ZN(n_1236));
   AOI21_X1 i_2_422_1 (.A(n_2_132), .B1(n_952), .B2(n_2_133), .ZN(n_2_422_0));
   INV_X1 i_2_422_2 (.A(n_2_134), .ZN(n_2_422_1));
   OAI21_X1 i_2_423_0 (.A(n_2_423_0), .B1(n_952), .B2(n_2_423_1), .ZN(n_1237));
   AOI21_X1 i_2_423_1 (.A(n_2_109), .B1(n_952), .B2(n_2_110), .ZN(n_2_423_0));
   INV_X1 i_2_423_2 (.A(n_2_111), .ZN(n_2_423_1));
   OAI21_X1 i_2_424_0 (.A(n_2_424_0), .B1(n_952), .B2(n_2_424_1), .ZN(n_1238));
   AOI21_X1 i_2_424_1 (.A(n_2_108), .B1(n_952), .B2(n_386), .ZN(n_2_424_0));
   INV_X1 i_2_424_2 (.A(n_387), .ZN(n_2_424_1));
   OAI21_X1 i_2_425_0 (.A(n_2_425_0), .B1(n_952), .B2(n_2_425_1), .ZN(n_1239));
   AOI21_X1 i_2_425_1 (.A(n_2_107), .B1(n_952), .B2(n_391), .ZN(n_2_425_0));
   INV_X1 i_2_425_2 (.A(n_392), .ZN(n_2_425_1));
   OAI21_X1 i_2_426_0 (.A(n_2_426_0), .B1(n_952), .B2(n_2_426_1), .ZN(n_1240));
   AOI21_X1 i_2_426_1 (.A(n_2_106), .B1(n_952), .B2(n_396), .ZN(n_2_426_0));
   INV_X1 i_2_426_2 (.A(n_397), .ZN(n_2_426_1));
   OAI21_X1 i_2_427_0 (.A(n_2_427_0), .B1(n_952), .B2(n_2_427_1), .ZN(n_1241));
   AOI21_X1 i_2_427_1 (.A(n_2_105), .B1(n_952), .B2(n_401), .ZN(n_2_427_0));
   INV_X1 i_2_427_2 (.A(n_402), .ZN(n_2_427_1));
   OAI21_X1 i_2_428_0 (.A(n_2_428_0), .B1(n_952), .B2(n_2_428_1), .ZN(n_1242));
   AOI21_X1 i_2_428_1 (.A(n_2_103), .B1(n_952), .B2(n_411), .ZN(n_2_428_0));
   INV_X1 i_2_428_2 (.A(n_412), .ZN(n_2_428_1));
   OAI21_X1 i_2_429_0 (.A(n_2_429_0), .B1(n_952), .B2(n_2_429_1), .ZN(n_1243));
   AOI21_X1 i_2_429_1 (.A(n_2_101), .B1(n_952), .B2(n_421), .ZN(n_2_429_0));
   INV_X1 i_2_429_2 (.A(n_422), .ZN(n_2_429_1));
   OAI21_X1 i_2_430_0 (.A(n_2_430_0), .B1(n_952), .B2(n_2_430_1), .ZN(n_1244));
   AOI21_X1 i_2_430_1 (.A(n_2_96), .B1(n_952), .B2(n_435), .ZN(n_2_430_0));
   INV_X1 i_2_430_2 (.A(n_436), .ZN(n_2_430_1));
   OAI21_X1 i_2_431_0 (.A(n_2_431_0), .B1(n_952), .B2(n_2_431_1), .ZN(n_1245));
   AOI21_X1 i_2_431_1 (.A(n_2_92), .B1(n_952), .B2(n_450), .ZN(n_2_431_0));
   INV_X1 i_2_431_2 (.A(n_451), .ZN(n_2_431_1));
   OAI21_X1 i_2_432_0 (.A(n_2_432_0), .B1(n_952), .B2(n_2_432_1), .ZN(n_1246));
   AOI21_X1 i_2_432_1 (.A(n_2_79), .B1(n_952), .B2(n_482), .ZN(n_2_432_0));
   INV_X1 i_2_432_2 (.A(n_483), .ZN(n_2_432_1));
   OAI21_X1 i_2_433_0 (.A(n_2_433_0), .B1(n_952), .B2(n_2_433_1), .ZN(n_1247));
   AOI21_X1 i_2_433_1 (.A(n_2_74), .B1(n_952), .B2(n_507), .ZN(n_2_433_0));
   INV_X1 i_2_433_2 (.A(n_508), .ZN(n_2_433_1));
   OAI21_X1 i_2_434_0 (.A(n_2_434_0), .B1(n_952), .B2(n_2_434_1), .ZN(n_1248));
   AOI21_X1 i_2_434_1 (.A(n_2_73), .B1(n_952), .B2(n_512), .ZN(n_2_434_0));
   INV_X1 i_2_434_2 (.A(n_513), .ZN(n_2_434_1));
   OAI21_X1 i_2_435_0 (.A(n_2_435_0), .B1(n_952), .B2(n_2_435_1), .ZN(n_1249));
   AOI21_X1 i_2_435_1 (.A(n_2_72), .B1(n_952), .B2(n_517), .ZN(n_2_435_0));
   INV_X1 i_2_435_2 (.A(n_518), .ZN(n_2_435_1));
   OAI21_X1 i_2_436_0 (.A(n_2_436_0), .B1(n_952), .B2(n_2_436_1), .ZN(n_1250));
   AOI21_X1 i_2_436_1 (.A(n_2_64), .B1(n_952), .B2(n_2_65), .ZN(n_2_436_0));
   INV_X1 i_2_436_2 (.A(n_2_66), .ZN(n_2_436_1));
   OAI21_X1 i_2_437_0 (.A(n_2_437_0), .B1(n_952), .B2(n_2_437_1), .ZN(n_1251));
   AOI21_X1 i_2_437_1 (.A(n_2_63), .B1(n_952), .B2(n_1291), .ZN(n_2_437_0));
   INV_X1 i_2_437_2 (.A(n_1292), .ZN(n_2_437_1));
   OAI21_X1 i_2_438_0 (.A(n_2_438_0), .B1(n_952), .B2(n_2_438_1), .ZN(n_1252));
   AOI21_X1 i_2_438_1 (.A(n_2_59), .B1(n_952), .B2(n_1293), .ZN(n_2_438_0));
   INV_X1 i_2_438_2 (.A(n_1294), .ZN(n_2_438_1));
   OAI21_X1 i_2_439_0 (.A(n_2_439_0), .B1(n_952), .B2(n_2_439_1), .ZN(n_1253));
   AOI21_X1 i_2_439_1 (.A(n_2_47), .B1(n_952), .B2(n_2_48), .ZN(n_2_439_0));
   INV_X1 i_2_439_2 (.A(n_2_49), .ZN(n_2_439_1));
   OAI21_X1 i_2_440_0 (.A(n_2_440_0), .B1(n_952), .B2(n_2_440_1), .ZN(n_1254));
   AOI21_X1 i_2_440_1 (.A(n_2_44), .B1(n_952), .B2(n_2_45), .ZN(n_2_440_0));
   INV_X1 i_2_440_2 (.A(n_2_46), .ZN(n_2_440_1));
   OAI21_X1 i_2_441_0 (.A(n_2_441_0), .B1(n_952), .B2(n_2_441_1), .ZN(n_1255));
   AOI21_X1 i_2_441_1 (.A(n_2_41), .B1(n_952), .B2(n_2_42), .ZN(n_2_441_0));
   INV_X1 i_2_441_2 (.A(n_2_43), .ZN(n_2_441_1));
   OAI21_X1 i_2_442_0 (.A(n_2_442_0), .B1(n_952), .B2(n_2_442_1), .ZN(n_1256));
   AOI21_X1 i_2_442_1 (.A(n_2_35), .B1(n_952), .B2(n_2_36), .ZN(n_2_442_0));
   INV_X1 i_2_442_2 (.A(n_2_37), .ZN(n_2_442_1));
   OAI21_X1 i_2_443_0 (.A(n_2_443_0), .B1(n_952), .B2(n_2_443_1), .ZN(n_1257));
   AOI21_X1 i_2_443_1 (.A(n_2_32), .B1(n_952), .B2(n_2_33), .ZN(n_2_443_0));
   INV_X1 i_2_443_2 (.A(n_2_34), .ZN(n_2_443_1));
   OAI21_X1 i_2_444_0 (.A(n_2_444_0), .B1(n_952), .B2(n_2_444_1), .ZN(n_1258));
   AOI21_X1 i_2_444_1 (.A(n_2_31), .B1(n_952), .B2(n_596), .ZN(n_2_444_0));
   INV_X1 i_2_444_2 (.A(n_597), .ZN(n_2_444_1));
   OAI21_X1 i_2_445_0 (.A(n_2_445_0), .B1(n_952), .B2(n_2_445_1), .ZN(n_1259));
   AOI21_X1 i_2_445_1 (.A(n_2_27), .B1(n_952), .B2(n_1295), .ZN(n_2_445_0));
   INV_X1 i_2_445_2 (.A(n_1296), .ZN(n_2_445_1));
   OAI21_X1 i_2_446_0 (.A(n_2_446_0), .B1(n_952), .B2(n_2_446_1), .ZN(n_1260));
   AOI21_X1 i_2_446_1 (.A(n_2_26), .B1(n_952), .B2(n_1297), .ZN(n_2_446_0));
   INV_X1 i_2_446_2 (.A(n_1298), .ZN(n_2_446_1));
   OAI21_X1 i_2_447_0 (.A(n_2_447_0), .B1(n_952), .B2(n_2_447_1), .ZN(n_1261));
   AOI21_X1 i_2_447_1 (.A(n_2_25), .B1(n_952), .B2(n_1299), .ZN(n_2_447_0));
   INV_X1 i_2_447_2 (.A(n_1300), .ZN(n_2_447_1));
   OAI21_X1 i_2_448_0 (.A(n_2_448_0), .B1(n_952), .B2(n_2_448_1), .ZN(n_1262));
   AOI21_X1 i_2_448_1 (.A(n_2_20), .B1(n_952), .B2(n_1301), .ZN(n_2_448_0));
   INV_X1 i_2_448_2 (.A(n_1302), .ZN(n_2_448_1));
   OAI21_X1 i_2_449_0 (.A(n_2_449_0), .B1(n_952), .B2(n_2_449_1), .ZN(n_1263));
   AOI21_X1 i_2_449_1 (.A(n_2_16), .B1(n_952), .B2(n_1303), .ZN(n_2_449_0));
   INV_X1 i_2_449_2 (.A(n_1304), .ZN(n_2_449_1));
   OAI21_X1 i_2_450_0 (.A(n_2_450_0), .B1(n_952), .B2(n_2_450_1), .ZN(n_1264));
   AOI21_X1 i_2_450_1 (.A(n_2_13), .B1(n_952), .B2(n_2_14), .ZN(n_2_450_0));
   INV_X1 i_2_450_2 (.A(n_2_15), .ZN(n_2_450_1));
   OAI21_X1 i_2_451_0 (.A(n_2_451_0), .B1(n_952), .B2(n_2_451_1), .ZN(n_1265));
   AOI21_X1 i_2_451_1 (.A(n_2_10), .B1(n_952), .B2(n_2_11), .ZN(n_2_451_0));
   INV_X1 i_2_451_2 (.A(n_2_12), .ZN(n_2_451_1));
   OAI21_X1 i_2_452_0 (.A(n_2_452_0), .B1(n_952), .B2(n_2_452_1), .ZN(n_1266));
   AOI21_X1 i_2_452_1 (.A(n_2_9), .B1(n_952), .B2(n_643), .ZN(n_2_452_0));
   INV_X1 i_2_452_2 (.A(n_644), .ZN(n_2_452_1));
   OAI21_X1 i_2_453_0 (.A(n_2_453_0), .B1(n_952), .B2(n_2_453_1), .ZN(n_1267));
   AOI21_X1 i_2_453_1 (.A(n_2_8), .B1(n_952), .B2(n_1307), .ZN(n_2_453_0));
   INV_X1 i_2_453_2 (.A(n_1308), .ZN(n_2_453_1));
   AND2_X1 i_2_454_0 (.A1(n_740), .A2(n_2_234), .ZN(n_2_11));
   OR2_X1 i_2_455_0 (.A1(n_2_234), .A2(n_740), .ZN(n_2_12));
   AND2_X1 i_2_456_0 (.A1(n_636), .A2(n_2_235), .ZN(n_2_14));
   OR2_X1 i_2_457_0 (.A1(n_2_235), .A2(n_636), .ZN(n_2_15));
   AND2_X1 i_2_458_0 (.A1(n_592), .A2(n_2_250), .ZN(n_2_33));
   OR2_X1 i_2_459_0 (.A1(n_2_250), .A2(n_592), .ZN(n_2_34));
   AND2_X1 i_2_460_0 (.A1(n_588), .A2(n_2_251), .ZN(n_2_36));
   OR2_X1 i_2_461_0 (.A1(n_2_251), .A2(n_588), .ZN(n_2_37));
   AND2_X1 i_2_462_0 (.A1(n_582), .A2(n_2_253), .ZN(n_2_42));
   OR2_X1 i_2_463_0 (.A1(n_2_253), .A2(n_582), .ZN(n_2_43));
   AND2_X1 i_2_464_0 (.A1(n_578), .A2(n_2_254), .ZN(n_2_45));
   OR2_X1 i_2_465_0 (.A1(n_2_254), .A2(n_578), .ZN(n_2_46));
   AND2_X1 i_2_466_0 (.A1(n_742), .A2(n_2_263), .ZN(n_2_65));
   OR2_X1 i_2_467_0 (.A1(n_2_263), .A2(n_742), .ZN(n_2_66));
   AND2_X1 i_2_468_0 (.A1(n_770), .A2(n_2_268), .ZN(n_2_110));
   OR2_X1 i_2_469_0 (.A1(n_2_268), .A2(n_770), .ZN(n_2_111));
   AND2_X1 i_2_470_0 (.A1(n_765), .A2(n_2_273), .ZN(n_2_133));
   OR2_X1 i_2_471_0 (.A1(n_2_273), .A2(n_765), .ZN(n_2_134));
   AND2_X1 i_2_472_0 (.A1(n_764), .A2(n_2_274), .ZN(n_2_136));
   OR2_X1 i_2_473_0 (.A1(n_2_274), .A2(n_764), .ZN(n_2_137));
   AND2_X1 i_2_474_0 (.A1(n_763), .A2(n_2_275), .ZN(n_2_140));
   OR2_X1 i_2_475_0 (.A1(n_2_275), .A2(n_763), .ZN(n_2_141));
   AND2_X1 i_2_476_0 (.A1(n_762), .A2(n_2_276), .ZN(n_2_144));
   OR2_X1 i_2_477_0 (.A1(n_2_276), .A2(n_762), .ZN(n_2_145));
   AND2_X1 i_2_478_0 (.A1(n_761), .A2(n_2_277), .ZN(n_2_148));
   OR2_X1 i_2_479_0 (.A1(n_2_277), .A2(n_761), .ZN(n_2_149));
   INV_X1 i_2_480_0 (.A(n_132), .ZN(n_2_480_0));
   AOI22_X1 i_2_480_1 (.A1(n_2_480_0), .A2(n_2_0), .B1(in_data[0]), .B2(n_132), 
      .ZN(n_2_480_1));
   INV_X1 i_2_480_2 (.A(n_2_480_1), .ZN(n_1268));
   AND2_X1 i_2_481_0 (.A1(n_754), .A2(n_2_284), .ZN(n_2_176));
   OR2_X1 i_2_482_0 (.A1(n_2_284), .A2(n_754), .ZN(n_2_177));
   AND2_X1 i_2_483_0 (.A1(n_756), .A2(n_2_282), .ZN(n_2_165));
   OR2_X1 i_2_484_0 (.A1(n_2_282), .A2(n_756), .ZN(n_2_166));
   INV_X1 i_2_485_0 (.A(n_2_485_0), .ZN(n_1269));
   OAI21_X1 i_2_485_1 (.A(n_2_485_1), .B1(n_1188), .B2(n_1309), .ZN(n_2_485_0));
   NAND2_X1 i_2_485_2 (.A1(n_1309), .A2(n_2_485_2), .ZN(n_2_485_1));
   INV_X1 i_2_485_3 (.A(in_data[0]), .ZN(n_2_485_2));
   AND2_X1 i_2_486_0 (.A1(n_574), .A2(n_2_255), .ZN(n_2_48));
   OR2_X1 i_2_487_0 (.A1(n_2_255), .A2(n_574), .ZN(n_2_49));
   datapath__1_14044 i_2_488 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, 1'b0}), .p_0(n_2_229));
   datapath__1_14076 i_2_489 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_2_230));
   datapath__1_14108 i_2_490 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, 1'b0, 1'b0}), .p_0(n_2_231));
   datapath__1_14300 i_2_491 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, 1'b0}), .p_0(n_2_238));
   datapath__1_14364 i_2_492 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, 1'b0, 1'b0}), .p_0(n_2_242));
   datapath__1_14396 i_2_493 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_2_243));
   datapath__1_14524 i_2_494 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_2_249));
   datapath__1_14652 i_2_495 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_2_252));
   datapath__1_14780 i_2_496 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_2_256));
   datapath__1_14812 i_2_497 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, 1'b0}), .p_0(n_2_257));
   datapath__1_14844 i_2_498 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_2_258));
   datapath__1_14908 i_2_499 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_2_260));
   datapath__1_15420 i_2_500 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_2_264));
   datapath__1_15452 i_2_501 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, 1'b0}), .p_0(n_2_265));
   datapath__1_15484 i_2_502 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_2_266));
   datapath__1_15516 i_2_503 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      1'b0, 1'b0, 1'b0, 1'b0}), .p_0(n_1270));
   datapath__1_15676 i_2_504 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_1271));
   datapath__1_15740 i_2_505 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_2_267));
   datapath__1_16117 i_2_506 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_2_269));
   datapath__1_16149 i_2_507 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, 1'b0, 1'b0}), .p_0(n_2_270));
   datapath__1_16309 i_2_508 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_2_271));
   datapath__1_16437 i_2_509 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_2_272));
   datapath__1_16725 i_2_510 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, 1'b0}), .p_0(n_2_278));
   datapath__1_16757 i_2_511 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_2_279));
   datapath__1_16821 i_2_512 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_2_280));
   datapath__1_16885 i_2_513 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_2_281));
   datapath__1_17109 i_2_514 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, 1'b0}), .p_0(n_2_283));
   datapath__1_17397 i_2_515 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_2_285));
   datapath__1_17461 i_2_516 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_2_286));
   datapath__1_17493 i_2_517 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, 1'b0}), .p_0(n_2_287));
   datapath__1_17525 i_2_518 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_2_288));
   datapath__1_17781 i_2_519 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_2_289));
   datapath__1_17877 i_2_520 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, 1'b0}), .p_0(n_2_290));
   datapath__1_17909 i_2_521 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_2_291));
   datapath__1_17973 i_2_522 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_1272));
   NAND2_X1 i_2_523_0 (.A1(n_2_523_0), .A2(n_2_523_1), .ZN(n_1273));
   INV_X1 i_2_523_1 (.A(n_2_232), .ZN(n_2_523_0));
   INV_X1 i_2_523_2 (.A(n_1267), .ZN(n_2_523_1));
   OR2_X1 i_2_524_0 (.A1(n_2_292), .A2(n_733), .ZN(n_2_232));
   OAI21_X1 i_2_525_0 (.A(n_2_525_0), .B1(n_2_525_1), .B2(n_2_232), .ZN(n_1274));
   NAND2_X1 i_2_525_1 (.A1(n_2_232), .A2(in_data[0]), .ZN(n_2_525_0));
   INV_X1 i_2_525_2 (.A(n_971), .ZN(n_2_525_1));
   datapath__1_13530 i_2_526 (.to_int6126({uc_193, \out_bs[7] [6], 
      \out_bs[7] [5], \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], 
      \out_bs[7] [1], \out_bs[7] [0]}), .p_0(n_2_292));
   AND2_X1 i_2_527_0 (.A1(n_2_292), .A2(n_733), .ZN(n_1275));
   NAND2_X1 i_2_528_0 (.A1(n_2_528_0), .A2(n_2_528_1), .ZN(n_1276));
   INV_X1 i_2_528_1 (.A(n_2_236), .ZN(n_2_528_0));
   INV_X1 i_2_528_2 (.A(n_1263), .ZN(n_2_528_1));
   OR2_X1 i_2_529_0 (.A1(n_2_293), .A2(n_730), .ZN(n_2_236));
   OAI21_X1 i_2_530_0 (.A(n_2_530_0), .B1(n_2_530_1), .B2(n_2_236), .ZN(n_1277));
   NAND2_X1 i_2_530_1 (.A1(n_2_236), .A2(in_data[0]), .ZN(n_2_530_0));
   INV_X1 i_2_530_2 (.A(n_972), .ZN(n_2_530_1));
   datapath__1_13546 i_2_531 (.to_int6126({uc_194, \out_bs[7] [6], 
      \out_bs[7] [5], \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], 
      \out_bs[7] [1], \out_bs[7] [0]}), .p_0(n_2_293));
   AND2_X1 i_2_532_0 (.A1(n_2_293), .A2(n_730), .ZN(n_1278));
   NAND2_X1 i_2_533_0 (.A1(n_2_533_0), .A2(n_2_533_1), .ZN(n_1279));
   INV_X1 i_2_533_1 (.A(n_2_239), .ZN(n_2_533_0));
   INV_X1 i_2_533_2 (.A(n_1262), .ZN(n_2_533_1));
   OR2_X1 i_2_534_0 (.A1(n_2_294), .A2(n_728), .ZN(n_2_239));
   OAI21_X1 i_2_535_0 (.A(n_2_535_0), .B1(n_2_535_1), .B2(n_2_239), .ZN(n_1280));
   NAND2_X1 i_2_535_1 (.A1(n_2_239), .A2(in_data[0]), .ZN(n_2_535_0));
   INV_X1 i_2_535_2 (.A(n_973), .ZN(n_2_535_1));
   datapath__1_13554 i_2_536 (.to_int6126({uc_195, \out_bs[7] [6], 
      \out_bs[7] [5], \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], 
      \out_bs[7] [1], \out_bs[7] [0]}), .p_0(n_2_294));
   AND2_X1 i_2_537_0 (.A1(n_2_294), .A2(n_728), .ZN(n_1281));
   OAI21_X1 i_2_538_0 (.A(n_2_538_0), .B1(n_2_538_1), .B2(n_2_245), .ZN(n_1282));
   NAND2_X1 i_2_538_1 (.A1(n_2_245), .A2(in_data[0]), .ZN(n_2_538_0));
   INV_X1 i_2_538_2 (.A(n_975), .ZN(n_2_538_1));
   NAND2_X1 i_2_539_0 (.A1(n_2_539_0), .A2(n_2_539_1), .ZN(n_1283));
   INV_X1 i_2_539_1 (.A(n_2_247), .ZN(n_2_539_0));
   INV_X1 i_2_539_2 (.A(n_1259), .ZN(n_2_539_1));
   OR2_X1 i_2_540_0 (.A1(n_2_296), .A2(n_724), .ZN(n_2_247));
   OAI21_X1 i_2_541_0 (.A(n_2_541_0), .B1(n_2_541_1), .B2(n_2_247), .ZN(n_1284));
   NAND2_X1 i_2_541_1 (.A1(n_2_247), .A2(in_data[0]), .ZN(n_2_541_0));
   INV_X1 i_2_541_2 (.A(n_977), .ZN(n_2_541_1));
   NAND2_X1 i_2_544_0 (.A1(n_2_544_0), .A2(n_2_544_1), .ZN(n_1285));
   INV_X1 i_2_544_1 (.A(n_2_261), .ZN(n_2_544_0));
   INV_X1 i_2_544_2 (.A(n_1251), .ZN(n_2_544_1));
   OR2_X1 i_2_545_0 (.A1(n_2_297), .A2(n_710), .ZN(n_2_261));
   OAI21_X1 i_2_546_0 (.A(n_2_546_0), .B1(n_2_546_1), .B2(n_2_261), .ZN(n_1286));
   NAND2_X1 i_2_546_1 (.A1(n_2_261), .A2(in_data[0]), .ZN(n_2_546_0));
   INV_X1 i_2_546_2 (.A(n_976), .ZN(n_2_546_1));
   datapath__1_13630 i_2_547 (.to_int6126({uc_196, \out_bs[7] [6], 
      \out_bs[7] [5], \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], 
      \out_bs[7] [1], uc_197}), .p_0(n_2_297));
   AND2_X1 i_2_548_0 (.A1(n_2_297), .A2(n_710), .ZN(n_1287));
   DFFS_X1 buf_is_empty_reg (.D(1'b0), .SN(n_2_373), .CK(n_2_298), .Q(
      buf_is_empty), .QN());
   NOR3_X1 i_2_549_0 (.A1(buf_is_empty), .A2(rst), .A3(n_2_549_68), .ZN(n_2_300));
   NOR2_X1 i_2_549_1 (.A1(n_2_549_1), .A2(n_2_549_0), .ZN(n_2_301));
   OAI22_X1 i_2_549_2 (.A1(n_904), .A2(n_2_549_64), .B1(n_2_549_63), .B2(n_983), 
      .ZN(n_2_549_0));
   OAI22_X1 i_2_549_3 (.A1(n_2_549_66), .A2(n_923), .B1(n_2_549_69), .B2(n_857), 
      .ZN(n_2_549_1));
   NOR2_X1 i_2_549_4 (.A1(n_2_549_3), .A2(n_2_549_2), .ZN(n_2_302));
   OAI22_X1 i_2_549_5 (.A1(n_905), .A2(n_2_549_64), .B1(n_2_549_63), .B2(n_882), 
      .ZN(n_2_549_2));
   OAI22_X1 i_2_549_6 (.A1(n_2_549_66), .A2(n_924), .B1(n_2_549_69), .B2(n_858), 
      .ZN(n_2_549_3));
   NOR2_X1 i_2_549_7 (.A1(n_2_549_5), .A2(n_2_549_4), .ZN(n_2_303));
   OAI22_X1 i_2_549_8 (.A1(n_906), .A2(n_2_549_64), .B1(n_2_549_63), .B2(n_883), 
      .ZN(n_2_549_4));
   OAI22_X1 i_2_549_9 (.A1(n_2_549_66), .A2(n_925), .B1(n_2_549_69), .B2(n_859), 
      .ZN(n_2_549_5));
   NOR2_X1 i_2_549_10 (.A1(n_2_549_7), .A2(n_2_549_6), .ZN(n_2_304));
   OAI22_X1 i_2_549_11 (.A1(n_907), .A2(n_2_549_64), .B1(n_2_549_63), .B2(n_884), 
      .ZN(n_2_549_6));
   OAI22_X1 i_2_549_12 (.A1(n_2_549_66), .A2(n_979), .B1(n_2_549_69), .B2(n_860), 
      .ZN(n_2_549_7));
   NOR2_X1 i_2_549_13 (.A1(n_2_549_9), .A2(n_2_549_8), .ZN(n_2_305));
   OAI22_X1 i_2_549_14 (.A1(n_908), .A2(n_2_549_64), .B1(n_2_549_63), .B2(n_982), 
      .ZN(n_2_549_8));
   OAI22_X1 i_2_549_15 (.A1(n_2_549_66), .A2(n_926), .B1(n_2_549_69), .B2(n_986), 
      .ZN(n_2_549_9));
   NOR2_X1 i_2_549_16 (.A1(n_2_549_11), .A2(n_2_549_10), .ZN(n_2_306));
   OAI22_X1 i_2_549_17 (.A1(n_998), .A2(n_2_549_64), .B1(n_2_549_63), .B2(n_885), 
      .ZN(n_2_549_10));
   OAI22_X1 i_2_549_18 (.A1(n_2_549_66), .A2(n_927), .B1(n_2_549_69), .B2(n_985), 
      .ZN(n_2_549_11));
   NOR2_X1 i_2_549_19 (.A1(n_2_549_13), .A2(n_2_549_12), .ZN(n_2_307));
   OAI22_X1 i_2_549_20 (.A1(n_909), .A2(n_2_549_64), .B1(n_2_549_63), .B2(n_886), 
      .ZN(n_2_549_12));
   OAI22_X1 i_2_549_21 (.A1(n_2_549_66), .A2(n_928), .B1(n_2_549_69), .B2(n_861), 
      .ZN(n_2_549_13));
   NOR2_X1 i_2_549_22 (.A1(n_2_549_15), .A2(n_2_549_14), .ZN(n_2_308));
   OAI22_X1 i_2_549_23 (.A1(n_1009), .A2(n_2_549_64), .B1(n_2_549_63), .B2(n_991), 
      .ZN(n_2_549_14));
   OAI22_X1 i_2_549_24 (.A1(n_2_549_66), .A2(n_929), .B1(n_2_549_69), .B2(n_862), 
      .ZN(n_2_549_15));
   NOR2_X1 i_2_549_25 (.A1(n_2_549_17), .A2(n_2_549_16), .ZN(n_2_309));
   OAI22_X1 i_2_549_26 (.A1(n_999), .A2(n_2_549_64), .B1(n_2_549_63), .B2(n_887), 
      .ZN(n_2_549_16));
   OAI22_X1 i_2_549_27 (.A1(n_2_549_66), .A2(n_930), .B1(n_2_549_69), .B2(n_863), 
      .ZN(n_2_549_17));
   NOR2_X1 i_2_549_28 (.A1(n_2_549_19), .A2(n_2_549_18), .ZN(n_2_310));
   OAI22_X1 i_2_549_29 (.A1(n_910), .A2(n_2_549_64), .B1(n_2_549_63), .B2(n_992), 
      .ZN(n_2_549_18));
   OAI22_X1 i_2_549_30 (.A1(n_2_549_66), .A2(n_931), .B1(n_2_549_69), .B2(n_987), 
      .ZN(n_2_549_19));
   NOR2_X1 i_2_549_31 (.A1(n_2_549_21), .A2(n_2_549_20), .ZN(n_2_311));
   OAI22_X1 i_2_549_32 (.A1(n_1000), .A2(n_2_549_64), .B1(n_2_549_63), .B2(n_888), 
      .ZN(n_2_549_20));
   OAI22_X1 i_2_549_33 (.A1(n_2_549_66), .A2(n_932), .B1(n_2_549_69), .B2(n_864), 
      .ZN(n_2_549_21));
   NOR2_X1 i_2_549_34 (.A1(n_2_549_23), .A2(n_2_549_22), .ZN(n_2_312));
   OAI22_X1 i_2_549_35 (.A1(n_1001), .A2(n_2_549_64), .B1(n_2_549_63), .B2(n_889), 
      .ZN(n_2_549_22));
   OAI22_X1 i_2_549_36 (.A1(n_2_549_66), .A2(n_933), .B1(n_2_549_69), .B2(n_865), 
      .ZN(n_2_549_23));
   NOR2_X1 i_2_549_37 (.A1(n_2_549_25), .A2(n_2_549_24), .ZN(n_2_313));
   OAI22_X1 i_2_549_38 (.A1(n_911), .A2(n_2_549_64), .B1(n_2_549_63), .B2(n_890), 
      .ZN(n_2_549_24));
   OAI22_X1 i_2_549_39 (.A1(n_2_549_66), .A2(n_934), .B1(n_2_549_69), .B2(n_988), 
      .ZN(n_2_549_25));
   NOR2_X1 i_2_549_40 (.A1(n_2_549_27), .A2(n_2_549_26), .ZN(n_2_314));
   OAI22_X1 i_2_549_41 (.A1(n_912), .A2(n_2_549_64), .B1(n_2_549_63), .B2(n_993), 
      .ZN(n_2_549_26));
   OAI22_X1 i_2_549_42 (.A1(n_2_549_66), .A2(n_935), .B1(n_2_549_69), .B2(n_866), 
      .ZN(n_2_549_27));
   NOR2_X1 i_2_549_43 (.A1(n_2_549_29), .A2(n_2_549_28), .ZN(n_2_315));
   OAI22_X1 i_2_549_44 (.A1(n_913), .A2(n_2_549_64), .B1(n_2_549_63), .B2(n_891), 
      .ZN(n_2_549_28));
   OAI22_X1 i_2_549_45 (.A1(n_2_549_66), .A2(n_936), .B1(n_2_549_69), .B2(n_867), 
      .ZN(n_2_549_29));
   NOR2_X1 i_2_549_46 (.A1(n_2_549_31), .A2(n_2_549_30), .ZN(n_2_316));
   OAI22_X1 i_2_549_47 (.A1(n_914), .A2(n_2_549_64), .B1(n_2_549_63), .B2(n_892), 
      .ZN(n_2_549_30));
   OAI22_X1 i_2_549_48 (.A1(n_2_549_66), .A2(n_937), .B1(n_2_549_69), .B2(n_868), 
      .ZN(n_2_549_31));
   NOR2_X1 i_2_549_49 (.A1(n_2_549_33), .A2(n_2_549_32), .ZN(n_2_317));
   OAI22_X1 i_2_549_50 (.A1(n_1002), .A2(n_2_549_64), .B1(n_2_549_63), .B2(n_893), 
      .ZN(n_2_549_32));
   OAI22_X1 i_2_549_51 (.A1(n_2_549_66), .A2(n_951), .B1(n_2_549_69), .B2(n_869), 
      .ZN(n_2_549_33));
   NOR2_X1 i_2_549_52 (.A1(n_2_549_35), .A2(n_2_549_34), .ZN(n_2_318));
   OAI22_X1 i_2_549_53 (.A1(n_1003), .A2(n_2_549_64), .B1(n_2_549_63), .B2(n_894), 
      .ZN(n_2_549_34));
   OAI22_X1 i_2_549_54 (.A1(n_2_549_66), .A2(n_978), .B1(n_2_549_69), .B2(n_870), 
      .ZN(n_2_549_35));
   NOR2_X1 i_2_549_55 (.A1(n_2_549_37), .A2(n_2_549_36), .ZN(n_2_319));
   OAI22_X1 i_2_549_56 (.A1(n_1004), .A2(n_2_549_64), .B1(n_2_549_63), .B2(n_895), 
      .ZN(n_2_549_36));
   OAI22_X1 i_2_549_57 (.A1(n_2_549_66), .A2(n_938), .B1(n_2_549_69), .B2(n_984), 
      .ZN(n_2_549_37));
   NOR2_X1 i_2_549_58 (.A1(n_2_549_39), .A2(n_2_549_38), .ZN(n_2_320));
   OAI22_X1 i_2_549_59 (.A1(n_915), .A2(n_2_549_64), .B1(n_2_549_63), .B2(n_896), 
      .ZN(n_2_549_38));
   OAI22_X1 i_2_549_60 (.A1(n_2_549_66), .A2(n_939), .B1(n_2_549_69), .B2(n_871), 
      .ZN(n_2_549_39));
   NOR2_X1 i_2_549_61 (.A1(n_2_549_41), .A2(n_2_549_40), .ZN(n_2_321));
   OAI22_X1 i_2_549_62 (.A1(n_1005), .A2(n_2_549_64), .B1(n_2_549_63), .B2(n_994), 
      .ZN(n_2_549_40));
   OAI22_X1 i_2_549_63 (.A1(n_2_549_66), .A2(n_940), .B1(n_2_549_69), .B2(n_872), 
      .ZN(n_2_549_41));
   NOR2_X1 i_2_549_64 (.A1(n_2_549_43), .A2(n_2_549_42), .ZN(n_2_322));
   OAI22_X1 i_2_549_65 (.A1(n_1006), .A2(n_2_549_64), .B1(n_2_549_63), .B2(n_995), 
      .ZN(n_2_549_42));
   OAI22_X1 i_2_549_66 (.A1(n_2_549_66), .A2(n_941), .B1(n_2_549_69), .B2(n_873), 
      .ZN(n_2_549_43));
   NOR2_X1 i_2_549_67 (.A1(n_2_549_45), .A2(n_2_549_44), .ZN(n_2_323));
   OAI22_X1 i_2_549_68 (.A1(n_1007), .A2(n_2_549_64), .B1(n_2_549_63), .B2(n_996), 
      .ZN(n_2_549_44));
   OAI22_X1 i_2_549_69 (.A1(n_2_549_66), .A2(n_942), .B1(n_2_549_69), .B2(n_874), 
      .ZN(n_2_549_45));
   NOR2_X1 i_2_549_70 (.A1(n_2_549_47), .A2(n_2_549_46), .ZN(n_2_324));
   OAI22_X1 i_2_549_71 (.A1(n_1008), .A2(n_2_549_64), .B1(n_2_549_63), .B2(n_997), 
      .ZN(n_2_549_46));
   OAI22_X1 i_2_549_72 (.A1(n_2_549_66), .A2(n_943), .B1(n_2_549_69), .B2(n_875), 
      .ZN(n_2_549_47));
   NOR2_X1 i_2_549_73 (.A1(n_2_549_49), .A2(n_2_549_48), .ZN(n_2_325));
   OAI22_X1 i_2_549_74 (.A1(n_980), .A2(n_2_549_64), .B1(n_2_549_63), .B2(n_897), 
      .ZN(n_2_549_48));
   OAI22_X1 i_2_549_75 (.A1(n_2_549_66), .A2(n_944), .B1(n_2_549_69), .B2(n_876), 
      .ZN(n_2_549_49));
   NOR2_X1 i_2_549_76 (.A1(n_2_549_51), .A2(n_2_549_50), .ZN(n_2_326));
   OAI22_X1 i_2_549_77 (.A1(n_916), .A2(n_2_549_64), .B1(n_2_549_63), .B2(n_898), 
      .ZN(n_2_549_50));
   OAI22_X1 i_2_549_78 (.A1(n_2_549_66), .A2(n_945), .B1(n_2_549_69), .B2(n_989), 
      .ZN(n_2_549_51));
   NOR2_X1 i_2_549_79 (.A1(n_2_549_53), .A2(n_2_549_52), .ZN(n_2_327));
   OAI22_X1 i_2_549_80 (.A1(n_917), .A2(n_2_549_64), .B1(n_2_549_63), .B2(n_899), 
      .ZN(n_2_549_52));
   OAI22_X1 i_2_549_81 (.A1(n_2_549_66), .A2(n_946), .B1(n_2_549_69), .B2(n_877), 
      .ZN(n_2_549_53));
   NOR2_X1 i_2_549_82 (.A1(n_2_549_55), .A2(n_2_549_54), .ZN(n_2_328));
   OAI22_X1 i_2_549_83 (.A1(n_918), .A2(n_2_549_64), .B1(n_2_549_63), .B2(n_900), 
      .ZN(n_2_549_54));
   OAI22_X1 i_2_549_84 (.A1(n_2_549_66), .A2(n_947), .B1(n_2_549_69), .B2(n_878), 
      .ZN(n_2_549_55));
   NOR2_X1 i_2_549_85 (.A1(n_2_549_57), .A2(n_2_549_56), .ZN(n_2_329));
   OAI22_X1 i_2_549_86 (.A1(n_919), .A2(n_2_549_64), .B1(n_2_549_63), .B2(n_901), 
      .ZN(n_2_549_56));
   OAI22_X1 i_2_549_87 (.A1(n_2_549_66), .A2(n_1010), .B1(n_2_549_69), .B2(n_879), 
      .ZN(n_2_549_57));
   NOR2_X1 i_2_549_88 (.A1(n_2_549_59), .A2(n_2_549_58), .ZN(n_2_330));
   OAI22_X1 i_2_549_89 (.A1(n_920), .A2(n_2_549_64), .B1(n_2_549_63), .B2(n_902), 
      .ZN(n_2_549_58));
   OAI22_X1 i_2_549_90 (.A1(n_2_549_66), .A2(n_948), .B1(n_2_549_69), .B2(n_880), 
      .ZN(n_2_549_59));
   NOR2_X1 i_2_549_91 (.A1(n_2_549_61), .A2(n_2_549_60), .ZN(n_2_331));
   OAI22_X1 i_2_549_92 (.A1(n_921), .A2(n_2_549_64), .B1(n_2_549_63), .B2(n_903), 
      .ZN(n_2_549_60));
   OAI22_X1 i_2_549_93 (.A1(n_2_549_66), .A2(n_949), .B1(n_2_549_69), .B2(n_881), 
      .ZN(n_2_549_61));
   NOR2_X1 i_2_549_94 (.A1(n_2_549_65), .A2(n_2_549_62), .ZN(n_2_332));
   OAI22_X1 i_2_549_95 (.A1(n_922), .A2(n_2_549_64), .B1(n_2_549_63), .B2(n_981), 
      .ZN(n_2_549_62));
   NAND2_X1 i_2_549_96 (.A1(n_2_549_78), .A2(buf_flush_i[6]), .ZN(n_2_549_63));
   NAND2_X1 i_2_549_97 (.A1(n_2_549_79), .A2(buf_flush_i[5]), .ZN(n_2_549_64));
   OAI22_X1 i_2_549_98 (.A1(n_2_549_66), .A2(n_950), .B1(n_2_549_69), .B2(n_990), 
      .ZN(n_2_549_65));
   NAND2_X1 i_2_549_99 (.A1(n_2_549_79), .A2(n_2_549_78), .ZN(n_2_549_66));
   NOR2_X1 i_2_549_100 (.A1(n_2_334), .A2(n_2_549_67), .ZN(n_2_333));
   OAI21_X1 i_2_549_101 (.A(state_wait), .B1(n_2_549_74), .B2(n_2_549_70), 
      .ZN(n_2_549_67));
   NOR2_X1 i_2_549_102 (.A1(buf_is_empty), .A2(n_2_549_68), .ZN(n_2_334));
   AOI22_X1 i_2_549_103 (.A1(n_2_549_74), .A2(n_2_549_71), .B1(n_2_549_70), 
      .B2(n_2_549_76), .ZN(n_2_549_68));
   NAND2_X1 i_2_549_104 (.A1(buf_flush_i[6]), .A2(buf_flush_i[5]), .ZN(
      n_2_549_69));
   OAI22_X1 i_2_549_105 (.A1(n_2_549_79), .A2(\out_as[0] [6]), .B1(n_2_549_78), 
      .B2(\out_as[0] [5]), .ZN(n_2_549_70));
   INV_X1 i_2_549_106 (.A(n_2_549_72), .ZN(n_2_549_71));
   AOI211_X1 i_2_549_107 (.A(buf_fill_flush_diff[6]), .B(buf_fill_flush_diff[5]), 
      .C1(\out_as[0] [1]), .C2(n_2_549_73), .ZN(n_2_549_72));
   AND4_X1 i_2_549_108 (.A1(\out_as[0] [4]), .A2(\out_as[0] [3]), .A3(
      \out_as[0] [2]), .A4(\out_as[0] [0]), .ZN(n_2_549_73));
   NAND3_X1 i_2_549_109 (.A1(n_2_549_77), .A2(n_2_549_75), .A3(n_2_549_76), 
      .ZN(n_2_549_74));
   AOI211_X1 i_2_549_110 (.A(\out_as[0] [4]), .B(\out_as[0] [3]), .C1(n_2_549_78), 
      .C2(\out_as[0] [5]), .ZN(n_2_549_75));
   NAND2_X1 i_2_549_111 (.A1(n_2_549_79), .A2(\out_as[0] [6]), .ZN(n_2_549_76));
   NOR3_X1 i_2_549_112 (.A1(\out_as[0] [2]), .A2(\out_as[0] [1]), .A3(
      \out_as[0] [0]), .ZN(n_2_549_77));
   INV_X1 i_2_549_113 (.A(rst), .ZN(n_2_373));
   INV_X1 i_2_549_114 (.A(buf_flush_i[5]), .ZN(n_2_549_78));
   INV_X1 i_2_549_115 (.A(buf_flush_i[6]), .ZN(n_2_549_79));
   DFFR_X1 out_ready_reg (.D(n_2_334), .RN(n_2_373), .CK(clk), .Q(out_ready), 
      .QN());
   DFFS_X1 error_success_reg (.D(n_2_335), .SN(n_2_373), .CK(clk), .Q(
      error_success), .QN());
   int_adder__parameterized1 fill_flush_diff_subtractor (.a({\out_as[0] [6], 
      \out_as[0] [5], uc_198, uc_199, uc_200, uc_201, uc_202}), .b({
      buf_flush_i_inv[6], buf_flush_i_inc[5], uc_203, uc_204, uc_205, uc_206, 
      uc_207}), .cin(), .enbl(), .c({buf_fill_flush_diff[6], 
      buf_fill_flush_diff[5], uc_208, uc_209, uc_210, uc_211, uc_212}), .cout());
   OR2_X1 i_2_550_0 (.A1(n_1260), .A2(n_2_245), .ZN(n_1288));
   OR2_X1 i_2_551_0 (.A1(n_2_295), .A2(n_737), .ZN(n_2_245));
   datapath__1_13570 i_2_552 (.to_int6126({uc_213, \out_bs[7] [6], 
      \out_bs[7] [5], \out_bs[7] [4], \out_bs[7] [3], \out_bs[7] [2], 
      \out_bs[7] [1], \out_bs[7] [0]}), .p_0(n_2_295));
   AND2_X1 i_2_553_0 (.A1(n_737), .A2(n_2_295), .ZN(n_1289));
   OR2_X1 i_2_554_0 (.A1(n_1240), .A2(n_855), .ZN(n_1290));
   AND2_X1 i_2_555_0 (.A1(n_550), .A2(n_2_262), .ZN(n_1291));
   OR2_X1 i_2_556_0 (.A1(n_2_262), .A2(n_550), .ZN(n_1292));
   AND2_X1 i_2_557_0 (.A1(n_558), .A2(n_2_259), .ZN(n_1293));
   OR2_X1 i_2_558_0 (.A1(n_2_259), .A2(n_558), .ZN(n_1294));
   AND2_X1 i_2_559_0 (.A1(n_605), .A2(n_2_248), .ZN(n_1295));
   OR2_X1 i_2_560_0 (.A1(n_2_248), .A2(n_605), .ZN(n_1296));
   AND2_X1 i_2_561_0 (.A1(n_741), .A2(n_2_246), .ZN(n_1297));
   OR2_X1 i_2_562_0 (.A1(n_2_246), .A2(n_741), .ZN(n_1298));
   AND2_X1 i_2_563_0 (.A1(n_612), .A2(n_2_244), .ZN(n_1299));
   OR2_X1 i_2_564_0 (.A1(n_2_244), .A2(n_612), .ZN(n_1300));
   AND2_X1 i_2_565_0 (.A1(n_624), .A2(n_2_240), .ZN(n_1301));
   OR2_X1 i_2_566_0 (.A1(n_2_240), .A2(n_624), .ZN(n_1302));
   AND2_X1 i_2_567_0 (.A1(n_632), .A2(n_2_237), .ZN(n_1303));
   OR2_X1 i_2_568_0 (.A1(n_2_237), .A2(n_632), .ZN(n_1304));
   OR2_X1 i_2_569_0 (.A1(n_1264), .A2(n_856), .ZN(n_1305));
   OR2_X1 i_2_570_0 (.A1(n_1265), .A2(n_854), .ZN(n_1306));
   AND2_X1 i_2_571_0 (.A1(n_648), .A2(n_2_233), .ZN(n_1307));
   OR2_X1 i_2_572_0 (.A1(n_2_233), .A2(n_648), .ZN(n_1308));
   datapath__1_14204 i_2_573 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_2_234));
   datapath__1_14236 i_2_574 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, 1'b0, 1'b0, 1'b0}), .p_0(n_2_235));
   datapath__1_14588 i_2_575 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_2_250));
   datapath__1_14620 i_2_576 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, 1'b0, 1'b0}), .p_0(n_2_251));
   datapath__1_14684 i_2_577 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, 1'b0}), .p_0(n_2_253));
   datapath__1_14716 i_2_578 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_2_254));
   datapath__1_14972 i_2_579 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_2_263));
   datapath__1_16053 i_2_580 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_2_268));
   datapath__1_16469 i_2_581 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, 1'b0}), .p_0(n_2_273));
   datapath__1_16501 i_2_582 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_2_274));
   datapath__1_16565 i_2_583 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_2_275));
   datapath__1_16629 i_2_584 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_2_276));
   datapath__1_16693 i_2_585 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_2_277));
   datapath__1_17301 i_2_586 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, 1'b0, 1'b0, 1'b0}), .p_0(n_2_284));
   datapath__1_17045 i_2_587 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0}), .p_0(n_2_282));
   AND2_X1 i_2_588_0 (.A1(n_716), .A2(n_853), .ZN(n_1309));
   datapath__1_14748 i_2_589 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, 1'b0, 1'b0, 1'b0}), .p_0(n_2_255));
   datapath__1_14940 i_2_590 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, 1'b0}), .p_0(n_2_262));
   datapath__1_14460 i_2_591 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_2_246));
   datapath__1_14428 i_2_592 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, 1'b0}), .p_0(n_2_244));
   datapath__1_14332 i_2_593 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_2_240));
   datapath__1_14268 i_2_594 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_2_237));
   datapath__1_14140 i_2_595 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, n_1311, \out_bs[6] [0]}), .p_0(n_2_233));
   datapath__1_14876 i_2_596 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      n_847, n_851, 1'b0, 1'b0}), .p_0(n_2_259));
   datapath__1_14492 i_2_597 (.to_int5359({1'b0, \out_bs[6] [6], n_1312, n_850, 
      1'b0, 1'b0, 1'b0, 1'b0}), .p_0(n_2_248));
   INV_X1 error_success_reg_enable_mux_0 (.A(error_success), .ZN(
      error_success_reg_enable_mux_n_0));
   NOR2_X1 error_success_reg_enable_mux_1 (.A1(error_success_reg_enable_mux_n_0), 
      .A2(n_2_333), .ZN(n_2_335));
   int_adder__parameterized0 buf_flush_i_adder (.a({buf_flush_i[6], 
      buf_flush_i[5], uc_214, uc_215, uc_216, uc_217, uc_218}), .b(), .cin(), 
      .enbl(), .c({buf_flush_i_inc[6], buf_flush_i_inc[5], uc_219, uc_220, 
      uc_221, uc_222, uc_223}), .cout());
   INV_X1 i_2_598_6 (.A(buf_flush_i[6]), .ZN(buf_flush_i_inv[6]));
   DFFS_X1 \buf_fill_i_reg[6]  (.D(\out_bs[7] [6]), .SN(n_2_373), .CK(n_2_298), 
      .Q(buf_fill_i[6]), .QN());
   DFFS_X2 \buf_fill_i_reg[5]  (.D(\out_bs[7] [5]), .SN(n_2_373), .CK(n_2_298), 
      .Q(buf_fill_i[5]), .QN());
   DFFS_X2 \buf_fill_i_reg[4]  (.D(\out_bs[7] [4]), .SN(n_2_373), .CK(n_2_298), 
      .Q(buf_fill_i[4]), .QN());
   DFFS_X1 \buf_fill_i_reg[3]  (.D(\out_bs[7] [3]), .SN(n_2_373), .CK(n_2_298), 
      .Q(buf_fill_i[3]), .QN());
   DFFS_X1 \buf_fill_i_reg[2]  (.D(\out_bs[7] [2]), .SN(n_2_373), .CK(n_2_298), 
      .Q(buf_fill_i[2]), .QN());
   DFFS_X1 \buf_fill_i_reg[1]  (.D(\out_bs[7] [1]), .SN(n_2_373), .CK(n_2_298), 
      .Q(buf_fill_i[1]), .QN());
   DFFS_X2 \buf_fill_i_reg[0]  (.D(\out_bs[7] [0]), .SN(n_2_373), .CK(n_2_298), 
      .Q(buf_fill_i[0]), .QN());
   CLKGATETST_X1 clk_gate_out_data_reg (.CK(clk), .E(n_2_300), .SE(1'b0), 
      .GCK(n_2_336));
   DFF_X1 \out_data_reg[31]  (.D(n_2_332), .CK(n_2_336), .Q(out_data[31]), .QN());
   DFF_X1 \out_data_reg[30]  (.D(n_2_331), .CK(n_2_336), .Q(out_data[30]), .QN());
   DFF_X1 \out_data_reg[29]  (.D(n_2_330), .CK(n_2_336), .Q(out_data[29]), .QN());
   DFF_X1 \out_data_reg[28]  (.D(n_2_329), .CK(n_2_336), .Q(out_data[28]), .QN());
   DFF_X1 \out_data_reg[27]  (.D(n_2_328), .CK(n_2_336), .Q(out_data[27]), .QN());
   DFF_X1 \out_data_reg[26]  (.D(n_2_327), .CK(n_2_336), .Q(out_data[26]), .QN());
   DFF_X1 \out_data_reg[25]  (.D(n_2_326), .CK(n_2_336), .Q(out_data[25]), .QN());
   DFF_X1 \out_data_reg[24]  (.D(n_2_325), .CK(n_2_336), .Q(out_data[24]), .QN());
   DFF_X1 \out_data_reg[23]  (.D(n_2_324), .CK(n_2_336), .Q(out_data[23]), .QN());
   DFF_X1 \out_data_reg[22]  (.D(n_2_323), .CK(n_2_336), .Q(out_data[22]), .QN());
   DFF_X1 \out_data_reg[21]  (.D(n_2_322), .CK(n_2_336), .Q(out_data[21]), .QN());
   DFF_X1 \out_data_reg[20]  (.D(n_2_321), .CK(n_2_336), .Q(out_data[20]), .QN());
   DFF_X1 \out_data_reg[19]  (.D(n_2_320), .CK(n_2_336), .Q(out_data[19]), .QN());
   DFF_X1 \out_data_reg[18]  (.D(n_2_319), .CK(n_2_336), .Q(out_data[18]), .QN());
   DFF_X1 \out_data_reg[17]  (.D(n_2_318), .CK(n_2_336), .Q(out_data[17]), .QN());
   DFF_X1 \out_data_reg[16]  (.D(n_2_317), .CK(n_2_336), .Q(out_data[16]), .QN());
   DFF_X1 \out_data_reg[15]  (.D(n_2_316), .CK(n_2_336), .Q(out_data[15]), .QN());
   DFF_X1 \out_data_reg[14]  (.D(n_2_315), .CK(n_2_336), .Q(out_data[14]), .QN());
   DFF_X1 \out_data_reg[13]  (.D(n_2_314), .CK(n_2_336), .Q(out_data[13]), .QN());
   DFF_X1 \out_data_reg[12]  (.D(n_2_313), .CK(n_2_336), .Q(out_data[12]), .QN());
   DFF_X1 \out_data_reg[11]  (.D(n_2_312), .CK(n_2_336), .Q(out_data[11]), .QN());
   DFF_X1 \out_data_reg[10]  (.D(n_2_311), .CK(n_2_336), .Q(out_data[10]), .QN());
   DFF_X1 \out_data_reg[9]  (.D(n_2_310), .CK(n_2_336), .Q(out_data[9]), .QN());
   DFF_X1 \out_data_reg[8]  (.D(n_2_309), .CK(n_2_336), .Q(out_data[8]), .QN());
   DFF_X1 \out_data_reg[7]  (.D(n_2_308), .CK(n_2_336), .Q(out_data[7]), .QN());
   DFF_X1 \out_data_reg[6]  (.D(n_2_307), .CK(n_2_336), .Q(out_data[6]), .QN());
   DFF_X1 \out_data_reg[5]  (.D(n_2_306), .CK(n_2_336), .Q(out_data[5]), .QN());
   DFF_X1 \out_data_reg[4]  (.D(n_2_305), .CK(n_2_336), .Q(out_data[4]), .QN());
   DFF_X1 \out_data_reg[3]  (.D(n_2_304), .CK(n_2_336), .Q(out_data[3]), .QN());
   DFF_X1 \out_data_reg[2]  (.D(n_2_303), .CK(n_2_336), .Q(out_data[2]), .QN());
   DFF_X1 \out_data_reg[1]  (.D(n_2_302), .CK(n_2_336), .Q(out_data[1]), .QN());
   DFF_X1 \out_data_reg[0]  (.D(n_2_301), .CK(n_2_336), .Q(out_data[0]), .QN());
   DFFR_X1 \buf_flush_i_reg[5]  (.D(n_2_337), .RN(n_2_373), .CK(clk), .Q(
      buf_flush_i[5]), .QN());
   MUX2_X1 \buf_flush_i_reg[5]_enable_mux_0  (.A(buf_flush_i[5]), .B(
      buf_flush_i_inc[5]), .S(n_2_334), .Z(n_2_337));
   DFFR_X1 \buf_flush_i_reg[6]  (.D(n_2_338), .RN(n_2_373), .CK(clk), .Q(
      buf_flush_i[6]), .QN());
   MUX2_X1 \buf_flush_i_reg[6]_enable_mux_0  (.A(buf_flush_i[6]), .B(
      buf_flush_i_inc[6]), .S(n_2_334), .Z(n_2_338));
   BUF_X1 rt_shieldBuf__15 (.A(n_2_345), .Z(\out_bs[0] [6]));
   BUF_X1 rt_shieldBuf__15__15__0 (.A(n_2_344), .Z(\out_bs[0] [5]));
   BUF_X1 rt_shieldBuf__15__15__1 (.A(n_2_343), .Z(\out_bs[0] [4]));
   BUF_X1 rt_shieldBuf__15__15__2 (.A(n_2_342), .Z(\out_bs[0] [3]));
   BUF_X1 rt_shieldBuf__15__15__3 (.A(n_2_341), .Z(\out_bs[0] [2]));
   BUF_X1 rt_shieldBuf__15__15__4 (.A(n_2_340), .Z(\out_bs[0] [1]));
   BUF_X1 rt_shieldBuf__15__15__5 (.A(n_2_348), .Z(\out_bs[1] [6]));
   BUF_X1 rt_shieldBuf__15__15__6 (.A(n_2_347), .Z(\out_bs[1] [2]));
   BUF_X1 rt_shieldBuf__15__15__7 (.A(n_2_346), .Z(\out_bs[1] [1]));
   BUF_X1 rt_shieldBuf__15__15__8 (.A(n_2_354), .Z(\out_bs[2] [6]));
   BUF_X1 rt_shieldBuf__15__15__9 (.A(n_2_353), .Z(\out_bs[2] [5]));
   BUF_X1 rt_shieldBuf__15__15__10 (.A(n_2_352), .Z(\out_bs[2] [4]));
   BUF_X1 rt_shieldBuf__15__15__11 (.A(n_2_351), .Z(\out_bs[2] [3]));
   BUF_X1 rt_shieldBuf__15__15__12 (.A(n_2_350), .Z(\out_bs[2] [2]));
   BUF_X1 rt_shieldBuf__15__15__13 (.A(n_2_349), .Z(\out_bs[2] [1]));
   BUF_X1 rt_shieldBuf__15__15__14 (.A(n_2_358), .Z(\out_bs[3] [6]));
   BUF_X1 rt_shieldBuf__15__15__15 (.A(n_2_357), .Z(\out_bs[3] [5]));
   BUF_X1 rt_shieldBuf__15__15__16 (.A(n_2_356), .Z(\out_bs[3] [4]));
   BUF_X1 rt_shieldBuf__15__15__17 (.A(n_2_355), .Z(\out_bs[3] [2]));
   BUF_X1 rt_shieldBuf__15__15__18 (.A(n_2_359), .Z(\out_bs[4] [6]));
   BUF_X1 rt_shieldBuf__15__15__19 (.A(\out_bs[5] [5]), .Z(n_2_368));
   BUF_X1 rt_shieldBuf__15__15__20 (.A(n_2_360), .Z(\out_bs[0] [0]));
   BUF_X1 rt_shieldBuf__15__15__21 (.A(n_2_362), .Z(\out_bs[1] [5]));
   BUF_X1 rt_shieldBuf__15__15__22 (.A(n_2_361), .Z(\out_bs[1] [0]));
   BUF_X1 rt_shieldBuf__15__15__23 (.A(n_2_364), .Z(\out_bs[3] [3]));
   BUF_X1 rt_shieldBuf__15__15__24 (.A(n_2_363), .Z(\out_bs[3] [1]));
   BUF_X1 rt_shieldBuf__15__15__25 (.A(n_2_367), .Z(\out_bs[4] [4]));
   BUF_X1 rt_shieldBuf__15__15__26 (.A(n_2_365), .Z(\out_bs[4] [2]));
   BUF_X1 rt_shieldBuf__15__15__27 (.A(n_1089), .Z(n_2_369));
   BUF_X1 rt_shieldBuf__15__15__28 (.A(n_2_366), .Z(\out_bs[4] [3]));
   BUF_X1 rt_shieldBuf__15__15__29 (.A(\out_bs[5] [1]), .Z(n_2_371));
   BUF_X1 rt_shieldBuf__15__15__30 (.A(n_2_299), .Z(\out_bs[4] [1]));
   BUF_X1 rt_shieldBuf__15__15__31 (.A(n_2_372), .Z(\out_bs[1] [4]));
   BUF_X1 rt_shieldBuf__15__15__32 (.A(n_2_370), .Z(\out_bs[1] [3]));
   NOR2_X1 i_2_542_2 (.A1(\out_bs[7] [5]), .A2(\out_bs[7] [4]), .ZN(n_2_542_0));
   INV_X1 i_2_542_0 (.A(\out_bs[7] [6]), .ZN(n_2_542_1));
   NAND2_X1 i_2_542_1 (.A1(n_2_542_1), .A2(n_2_542_0), .ZN(n_2_296));
   INV_X1 i_2_542_3 (.A(n_2_542_0), .ZN(n_2_542_2));
   NAND2_X1 i_2_542_4 (.A1(n_724), .A2(n_2_542_2), .ZN(n_2_542_3));
   INV_X1 i_2_542_5 (.A(n_724), .ZN(n_2_542_4));
   OAI21_X1 i_2_542_6 (.A(n_2_542_3), .B1(n_2_542_1), .B2(n_2_542_4), .ZN(n_1310));
   BUF_X1 rt_shieldBuf__9 (.A(\out_bs[6] [1]), .Z(n_1311));
   BUF_X1 rt_shieldBuf__10 (.A(\out_bs[6] [5]), .Z(n_1312));
   BUF_X1 rt_shieldBuf__11 (.A(\out_bs[5] [1]), .Z(n_1313));
endmodule

module full_adder__4_196(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(f));
   AND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(cout));
endmodule

module full_adder__4_200(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(f));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(cin), .B1(a), .B2(b), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module full_adder__4_204(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__4_208(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__4_212(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__4_216(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__4_220(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__4_224(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__4_228(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__4_232(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__4_236(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__4_240(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__4_244(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__4_248(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__4_252(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__4_0(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
endmodule

module int_adder__parameterized2(a, b, cin, enbl, c, cout);
   input [15:0]a;
   input [1:0]b;
   input cin;
   input enbl;
   output [15:0]c;
   output cout;

   full_adder__4_196 full_adder_0_0_full_adder_0_i (.a(a[0]), .b(b[0]), .cin(), 
      .f(c[0]), .cout(n_0));
   full_adder__4_200 full_adder_0_1_full_adder_0_i (.a(a[1]), .b(b[1]), .cin(n_0), 
      .f(c[1]), .cout(n_1));
   full_adder__4_204 full_adder_0_2_full_adder_0_i (.a(a[2]), .b(), .cin(n_1), 
      .f(c[2]), .cout(n_2));
   full_adder__4_208 full_adder_0_3_full_adder_0_i (.a(a[3]), .b(), .cin(n_2), 
      .f(c[3]), .cout(n_3));
   full_adder__4_212 full_adder_0_4_full_adder_0_i (.a(a[4]), .b(), .cin(n_3), 
      .f(c[4]), .cout(n_4));
   full_adder__4_216 full_adder_0_5_full_adder_0_i (.a(a[5]), .b(), .cin(n_4), 
      .f(c[5]), .cout(n_5));
   full_adder__4_220 full_adder_0_6_full_adder_0_i (.a(a[6]), .b(), .cin(n_5), 
      .f(c[6]), .cout(n_6));
   full_adder__4_224 full_adder_0_7_full_adder_0_i (.a(a[7]), .b(), .cin(n_6), 
      .f(c[7]), .cout(n_7));
   full_adder__4_228 full_adder_0_8_full_adder_0_i (.a(a[8]), .b(), .cin(n_7), 
      .f(c[8]), .cout(n_8));
   full_adder__4_232 full_adder_0_9_full_adder_0_i (.a(a[9]), .b(), .cin(n_8), 
      .f(c[9]), .cout(n_9));
   full_adder__4_236 full_adder_0_10_full_adder_0_i (.a(a[10]), .b(), .cin(n_9), 
      .f(c[10]), .cout(n_10));
   full_adder__4_240 full_adder_0_11_full_adder_0_i (.a(a[11]), .b(), .cin(n_10), 
      .f(c[11]), .cout(n_11));
   full_adder__4_244 full_adder_0_12_full_adder_0_i (.a(a[12]), .b(), .cin(n_11), 
      .f(c[12]), .cout(n_12));
   full_adder__4_248 full_adder_0_13_full_adder_0_i (.a(a[13]), .b(), .cin(n_12), 
      .f(c[13]), .cout(n_13));
   full_adder__4_252 full_adder_0_14_full_adder_0_i (.a(a[14]), .b(), .cin(n_13), 
      .f(c[14]), .cout(n_14));
   full_adder__4_0 full_adder_0_15_full_adder_0_i (.a(a[15]), .b(), .cin(n_14), 
      .f(c[15]), .cout());
endmodule

module datapath__0_5921(b, a, i);
   input [2:0]b;
   input [15:0]a;
   output [15:0]i;

   FA_X1 i_147 (.A(n_8), .B(n_7), .CI(n_30), .CO(n_0), .S(i[3]));
   FA_X1 i_148 (.A(n_6), .B(n_5), .CI(n_0), .CO(n_1), .S(i[4]));
   FA_X1 i_149 (.A(n_4), .B(n_11), .CI(n_1), .CO(n_2), .S(i[5]));
   FA_X1 i_150 (.A(n_12), .B(n_23), .CI(n_2), .CO(n_3), .S(i[6]));
   FA_X1 i_151 (.A(n_24), .B(n_25), .CI(n_3), .CO(i[8]), .S(i[7]));
   NOR2_X1 i_0 (.A1(n_9), .A2(n_24), .ZN(n_23));
   AND2_X1 i_1 (.A1(n_21), .A2(n_25), .ZN(n_24));
   AND2_X1 i_2 (.A1(b[2]), .A2(a[5]), .ZN(n_25));
   AOI22_X1 i_3 (.A1(b[1]), .A2(a[5]), .B1(b[2]), .B2(a[4]), .ZN(n_9));
   OAI21_X1 i_4 (.A(n_13), .B1(n_16), .B2(n_15), .ZN(n_12));
   XOR2_X1 i_5 (.A(n_16), .B(n_10), .Z(n_11));
   NAND2_X1 i_6 (.A1(n_14), .A2(n_13), .ZN(n_10));
   NAND3_X1 i_7 (.A1(b[0]), .A2(a[5]), .A3(n_21), .ZN(n_13));
   INV_X1 i_8 (.A(n_15), .ZN(n_14));
   AOI21_X1 i_9 (.A(n_21), .B1(b[0]), .B2(a[5]), .ZN(n_15));
   NAND2_X1 i_10 (.A1(b[2]), .A2(a[3]), .ZN(n_16));
   OAI21_X1 i_11 (.A(n_20), .B1(n_22), .B2(n_19), .ZN(n_4));
   XOR2_X1 i_12 (.A(n_22), .B(n_17), .Z(n_5));
   NAND2_X1 i_13 (.A1(n_20), .A2(n_18), .ZN(n_17));
   INV_X1 i_14 (.A(n_19), .ZN(n_18));
   AOI22_X1 i_15 (.A1(b[1]), .A2(a[3]), .B1(b[0]), .B2(a[4]), .ZN(n_19));
   NAND3_X1 i_16 (.A1(b[0]), .A2(a[3]), .A3(n_21), .ZN(n_20));
   AND2_X1 i_17 (.A1(b[1]), .A2(a[4]), .ZN(n_21));
   NAND2_X1 i_18 (.A1(b[2]), .A2(a[2]), .ZN(n_22));
   OAI21_X1 i_19 (.A(n_29), .B1(n_37), .B2(n_31), .ZN(n_6));
   INV_X1 i_20 (.A(n_26), .ZN(n_30));
   AOI22_X1 i_21 (.A1(n_38), .A2(n_34), .B1(n_39), .B2(n_33), .ZN(n_26));
   XOR2_X1 i_22 (.A(n_36), .B(n_27), .Z(n_7));
   NOR2_X1 i_23 (.A1(n_31), .A2(n_28), .ZN(n_27));
   INV_X1 i_24 (.A(n_29), .ZN(n_28));
   NAND3_X1 i_25 (.A1(b[1]), .A2(a[3]), .A3(n_38), .ZN(n_29));
   AOI22_X1 i_26 (.A1(b[0]), .A2(a[3]), .B1(b[1]), .B2(a[2]), .ZN(n_31));
   NOR2_X1 i_27 (.A1(n_39), .A2(n_32), .ZN(i[1]));
   AOI22_X1 i_28 (.A1(b[1]), .A2(a[0]), .B1(b[0]), .B2(a[1]), .ZN(n_32));
   XNOR2_X1 i_29 (.A(n_40), .B(n_33), .ZN(i[2]));
   XOR2_X1 i_30 (.A(n_38), .B(n_34), .Z(n_33));
   NOR2_X1 i_31 (.A1(n_8), .A2(n_35), .ZN(n_34));
   AOI22_X1 i_32 (.A1(b[1]), .A2(a[1]), .B1(b[2]), .B2(a[0]), .ZN(n_35));
   AND3_X1 i_33 (.A1(b[1]), .A2(a[0]), .A3(n_36), .ZN(n_8));
   INV_X1 i_34 (.A(n_37), .ZN(n_36));
   NAND2_X1 i_35 (.A1(b[2]), .A2(a[1]), .ZN(n_37));
   AND2_X1 i_36 (.A1(b[0]), .A2(a[2]), .ZN(n_38));
   INV_X1 i_37 (.A(n_40), .ZN(n_39));
   NAND3_X1 i_38 (.A1(b[1]), .A2(a[1]), .A3(i[0]), .ZN(n_40));
   AND2_X1 i_39 (.A1(b[0]), .A2(a[0]), .ZN(i[0]));
endmodule

module int_multiplier__parameterized0(a, b, enbl, c);
   input [15:0]a;
   input [2:0]b;
   input enbl;
   output [15:0]c;

   datapath__0_5921 i_0 (.b(b), .a({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      uc_0, uc_1, uc_2, a[5], a[4], a[3], a[2], a[1], a[0]}), .i({uc_3, uc_4, 
      uc_5, uc_6, uc_7, uc_8, uc_9, c[8], c[7], c[6], c[5], c[4], c[3], c[2], 
      c[1], c[0]}));
endmodule

module full_adder__4_312(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   INV_X1 i_3 (.A(b), .ZN(f));
endmodule

module full_adder__4_308(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(b), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(b), .ZN(cout));
endmodule

module full_adder__4_304(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XNOR2_X1 i_0_0 (.A(b), .B(cin), .ZN(f));
   OR2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(cout));
endmodule

module full_adder__4_300(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XNOR2_X1 i_0_0 (.A(b), .B(cin), .ZN(f));
   OR2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(cout));
endmodule

module full_adder__4_296(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(b), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(b), .ZN(cout));
endmodule

module full_adder__4_292(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XNOR2_X1 i_0_0 (.A(b), .B(cin), .ZN(f));
   OR2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(cout));
endmodule

module full_adder__4_288(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XNOR2_X1 i_0_0 (.A(b), .B(cin), .ZN(f));
   OR2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(cout));
endmodule

module full_adder__4_284(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XNOR2_X1 i_0_0 (.A(b), .B(cin), .ZN(f));
   OR2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(cout));
endmodule

module full_adder__4_280(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(b), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(b), .ZN(cout));
endmodule

module int_adder__parameterized3__4_317(a, b, cin, enbl, c, cout);
   input [15:0]a;
   input [15:0]b;
   input cin;
   input enbl;
   output [15:0]c;
   output cout;

   full_adder__4_312 full_adder_0_1_full_adder_0_i (.a(), .b(b[1]), .cin(), 
      .f(c[1]), .cout());
   full_adder__4_308 full_adder_0_2_full_adder_0_i (.a(), .b(b[2]), .cin(b[1]), 
      .f(c[2]), .cout(n_2));
   full_adder__4_304 full_adder_0_3_full_adder_0_i (.a(), .b(b[3]), .cin(n_2), 
      .f(c[3]), .cout(n_3));
   full_adder__4_300 full_adder_0_4_full_adder_0_i (.a(), .b(b[4]), .cin(n_3), 
      .f(c[4]), .cout(n_4));
   full_adder__4_296 full_adder_0_5_full_adder_0_i (.a(), .b(b[5]), .cin(n_4), 
      .f(c[5]), .cout(n_5));
   full_adder__4_292 full_adder_0_6_full_adder_0_i (.a(), .b(b[6]), .cin(n_5), 
      .f(c[6]), .cout(n_6));
   full_adder__4_288 full_adder_0_7_full_adder_0_i (.a(), .b(b[7]), .cin(n_6), 
      .f(c[7]), .cout(n_0));
   full_adder__4_284 full_adder_0_8_full_adder_0_i (.a(), .b(b[8]), .cin(n_0), 
      .f(c[8]), .cout(n_1));
   full_adder__4_280 full_adder_0_9_full_adder_0_i (.a(), .b(b[9]), .cin(n_1), 
      .f(c[9]), .cout(c[10]));
endmodule

module full_adder__4_440(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   INV_X1 i_3 (.A(b), .ZN(f));
endmodule

module full_adder__4_436(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XNOR2_X1 i_0_0 (.A(b), .B(cin), .ZN(f));
   OR2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(cout));
endmodule

module full_adder__4_432(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(b), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(b), .ZN(cout));
endmodule

module full_adder__4_428(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XNOR2_X1 i_0_0 (.A(b), .B(cin), .ZN(f));
   OR2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(cout));
endmodule

module full_adder__4_424(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   INV_X1 i_3 (.A(cin), .ZN(f));
endmodule

module int_adder__parameterized4__4_449(a, b, cin, enbl, c, cout);
   input [15:0]a;
   input [5:0]b;
   input cin;
   input enbl;
   output [15:0]c;
   output cout;

   full_adder__4_440 full_adder_0_2_full_adder_0_i (.a(), .b(b[2]), .cin(), 
      .f(c[2]), .cout());
   full_adder__4_436 full_adder_0_3_full_adder_0_i (.a(), .b(b[3]), .cin(b[2]), 
      .f(c[3]), .cout(n_0));
   full_adder__4_432 full_adder_0_4_full_adder_0_i (.a(), .b(b[4]), .cin(n_0), 
      .f(c[4]), .cout(n_1));
   full_adder__4_428 full_adder_0_5_full_adder_0_i (.a(), .b(b[5]), .cin(n_1), 
      .f(c[5]), .cout(c[7]));
   full_adder__4_424 full_adder_0_6_full_adder_0_i (.a(), .b(), .cin(c[7]), 
      .f(c[6]), .cout());
endmodule

module full_adder__4_76(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   INV_X1 i_3 (.A(b), .ZN(f));
endmodule

module full_adder__4_80(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(b), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(b), .ZN(cout));
endmodule

module full_adder__4_84(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XNOR2_X1 i_0_0 (.A(b), .B(cin), .ZN(f));
   OR2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(cout));
endmodule

module full_adder__4_88(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(b), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(b), .ZN(cout));
endmodule

module int_adder__parameterized4(a, b, cin, enbl, c, cout);
   input [15:0]a;
   input [5:0]b;
   input cin;
   input enbl;
   output [15:0]c;
   output cout;

   full_adder__4_76 full_adder_0_2_full_adder_0_i (.a(), .b(b[2]), .cin(), 
      .f(c[2]), .cout());
   full_adder__4_80 full_adder_0_3_full_adder_0_i (.a(), .b(b[3]), .cin(b[2]), 
      .f(c[3]), .cout(n_0));
   full_adder__4_84 full_adder_0_4_full_adder_0_i (.a(), .b(b[4]), .cin(n_0), 
      .f(c[4]), .cout(n_1));
   full_adder__4_88 full_adder_0_5_full_adder_0_i (.a(), .b(b[5]), .cin(n_1), 
      .f(c[5]), .cout(c[6]));
endmodule

module datapath__4_383(to_int6153, to_int, i);
   input [16:0]to_int6153;
   input [16:0]to_int;
   output [31:0]i;

   HA_X1 i_164 (.A(n_20), .B(n_19), .CO(n_12), .S(n_11));
   FA_X1 i_179 (.A(n_18), .B(n_17), .CI(n_28), .CO(n_40), .S(n_39));
   HA_X1 i_180 (.A(n_16), .B(n_12), .CO(n_42), .S(n_41));
   FA_X1 i_203 (.A(n_54), .B(n_44), .CI(n_66), .CO(n_69), .S(n_68));
   HA_X1 i_204 (.A(n_42), .B(n_40), .CO(n_77), .S(n_76));
   FA_X1 i_227 (.A(n_51), .B(n_15), .CI(n_55), .CO(n_87), .S(n_86));
   FA_X1 i_228 (.A(n_81), .B(n_78), .CI(n_77), .CO(n_89), .S(n_88));
   HA_X1 i_229 (.A(n_86), .B(n_69), .CO(n_91), .S(n_90));
   FA_X1 i_253 (.A(n_82), .B(n_87), .CI(n_91), .CO(n_100), .S(n_99));
   HA_X1 i_254 (.A(n_89), .B(n_94), .CO(n_102), .S(n_101));
   FA_X1 i_286 (.A(1'b0), .B(n_104), .CI(n_95), .CO(n_107), .S(n_106));
   HA_X1 i_287 (.A(n_102), .B(n_100), .CO(n_109), .S(n_108));
   FA_X1 i_320 (.A(1'b0), .B(n_110), .CI(n_105), .CO(n_112), .S(n_111));
   HA_X1 i_321 (.A(n_109), .B(n_107), .CO(n_114), .S(n_113));
   HA_X1 i_355 (.A(n_114), .B(n_112), .CO(n_116), .S(n_115));
   FA_X1 i_522 (.A(n_14), .B(n_13), .CI(n_10), .CO(n_0), .S(i[3]));
   FA_X1 i_523 (.A(n_9), .B(n_11), .CI(n_0), .CO(n_1), .S(i[4]));
   FA_X1 i_524 (.A(n_41), .B(n_39), .CI(n_1), .CO(n_2), .S(i[5]));
   FA_X1 i_525 (.A(n_76), .B(n_68), .CI(n_2), .CO(n_3), .S(i[6]));
   FA_X1 i_526 (.A(n_88), .B(n_90), .CI(n_3), .CO(n_4), .S(i[7]));
   FA_X1 i_527 (.A(n_99), .B(n_101), .CI(n_4), .CO(n_5), .S(i[8]));
   FA_X1 i_528 (.A(n_108), .B(n_106), .CI(n_5), .CO(n_6), .S(i[9]));
   FA_X1 i_529 (.A(n_113), .B(n_111), .CI(n_6), .CO(n_7), .S(i[10]));
   FA_X1 i_530 (.A(1'b0), .B(n_115), .CI(n_7), .CO(n_8), .S(i[11]));
   XNOR2_X1 i_0 (.A(n_73), .B(n_21), .ZN(n_9));
   NOR2_X1 i_1 (.A1(n_65), .A2(n_63), .ZN(n_21));
   OAI21_X1 i_2 (.A(n_92), .B1(n_79), .B2(to_int6153[2]), .ZN(n_10));
   XNOR2_X1 i_3 (.A(n_71), .B(n_22), .ZN(n_13));
   NOR2_X1 i_4 (.A1(n_74), .A2(n_72), .ZN(n_22));
   XOR2_X1 i_5 (.A(n_84), .B(n_61), .Z(n_14));
   OAI22_X1 i_6 (.A1(n_25), .A2(n_29), .B1(n_33), .B2(n_27), .ZN(n_95));
   NOR2_X1 i_7 (.A1(n_23), .A2(n_105), .ZN(n_104));
   AND3_X1 i_8 (.A1(to_int6153[4]), .A2(to_int[4]), .A3(n_110), .ZN(n_105));
   AND2_X1 i_9 (.A1(to_int6153[5]), .A2(to_int[5]), .ZN(n_110));
   AOI22_X1 i_10 (.A1(to_int6153[4]), .A2(to_int[5]), .B1(to_int[4]), .B2(
      to_int6153[5]), .ZN(n_23));
   XNOR2_X1 i_11 (.A(n_29), .B(n_24), .ZN(n_94));
   NOR2_X1 i_12 (.A1(n_26), .A2(n_25), .ZN(n_24));
   AOI22_X1 i_13 (.A1(to_int6153[3]), .A2(to_int[5]), .B1(to_int[4]), .B2(
      to_int6153[4]), .ZN(n_25));
   NOR2_X1 i_14 (.A1(n_33), .A2(n_27), .ZN(n_26));
   NAND2_X1 i_15 (.A1(to_int6153[4]), .A2(to_int[5]), .ZN(n_27));
   NAND2_X1 i_16 (.A1(to_int6153[5]), .A2(to_int[3]), .ZN(n_29));
   AND2_X1 i_17 (.A1(n_32), .A2(n_30), .ZN(n_82));
   OAI21_X1 i_18 (.A(n_34), .B1(n_33), .B2(n_47), .ZN(n_30));
   XNOR2_X1 i_19 (.A(n_34), .B(n_31), .ZN(n_81));
   XOR2_X1 i_20 (.A(n_47), .B(n_33), .Z(n_31));
   NAND2_X1 i_21 (.A1(n_47), .A2(n_33), .ZN(n_32));
   NAND2_X1 i_22 (.A1(to_int6153[3]), .A2(to_int[4]), .ZN(n_33));
   NAND2_X1 i_23 (.A1(to_int6153[4]), .A2(to_int[3]), .ZN(n_34));
   OAI22_X1 i_24 (.A1(n_45), .A2(n_48), .B1(n_60), .B2(n_47), .ZN(n_55));
   NOR2_X1 i_25 (.A1(n_15), .A2(n_35), .ZN(n_66));
   NOR2_X1 i_26 (.A1(n_37), .A2(n_36), .ZN(n_35));
   AND2_X1 i_27 (.A1(n_37), .A2(n_36), .ZN(n_15));
   OAI22_X1 i_28 (.A1(n_57), .A2(n_62), .B1(n_70), .B2(n_59), .ZN(n_36));
   OAI22_X1 i_29 (.A1(n_50), .A2(n_53), .B1(n_64), .B2(n_73), .ZN(n_37));
   XOR2_X1 i_30 (.A(n_64), .B(n_38), .Z(n_44));
   NOR2_X1 i_31 (.A1(n_64), .A2(n_38), .ZN(n_51));
   AND2_X1 i_32 (.A1(to_int6153[5]), .A2(to_int[2]), .ZN(n_78));
   NAND2_X1 i_33 (.A1(to_int6153[5]), .A2(to_int[1]), .ZN(n_38));
   XNOR2_X1 i_34 (.A(n_48), .B(n_43), .ZN(n_54));
   NOR2_X1 i_35 (.A1(n_46), .A2(n_45), .ZN(n_43));
   AOI22_X1 i_36 (.A1(to_int6153[1]), .A2(to_int[5]), .B1(to_int[4]), .B2(
      to_int6153[2]), .ZN(n_45));
   NOR2_X1 i_37 (.A1(n_60), .A2(n_47), .ZN(n_46));
   NAND2_X1 i_38 (.A1(to_int6153[2]), .A2(to_int[5]), .ZN(n_47));
   NAND2_X1 i_39 (.A1(to_int6153[3]), .A2(to_int[3]), .ZN(n_48));
   XNOR2_X1 i_40 (.A(n_53), .B(n_49), .ZN(n_16));
   NOR2_X1 i_41 (.A1(n_52), .A2(n_50), .ZN(n_49));
   AOI22_X1 i_42 (.A1(to_int6153[3]), .A2(to_int[2]), .B1(to_int[1]), .B2(
      to_int6153[4]), .ZN(n_50));
   NOR2_X1 i_43 (.A1(n_73), .A2(n_64), .ZN(n_52));
   NAND2_X1 i_44 (.A1(to_int6153[5]), .A2(to_int[0]), .ZN(n_53));
   XNOR2_X1 i_45 (.A(n_62), .B(n_56), .ZN(n_28));
   NOR2_X1 i_46 (.A1(n_58), .A2(n_57), .ZN(n_56));
   AOI22_X1 i_47 (.A1(to_int6153[0]), .A2(to_int[5]), .B1(to_int[4]), .B2(
      to_int6153[1]), .ZN(n_57));
   NOR2_X1 i_48 (.A1(n_70), .A2(n_59), .ZN(n_58));
   NAND2_X1 i_49 (.A1(to_int6153[1]), .A2(to_int[5]), .ZN(n_59));
   AOI21_X1 i_50 (.A(n_61), .B1(n_60), .B2(n_84), .ZN(n_17));
   NAND2_X1 i_51 (.A1(to_int6153[1]), .A2(to_int[4]), .ZN(n_60));
   NAND2_X1 i_52 (.A1(to_int6153[0]), .A2(to_int[3]), .ZN(n_61));
   NAND2_X1 i_53 (.A1(to_int6153[2]), .A2(to_int[3]), .ZN(n_62));
   OAI22_X1 i_54 (.A1(n_65), .A2(n_73), .B1(n_96), .B2(n_64), .ZN(n_18));
   NOR2_X1 i_55 (.A1(n_96), .A2(n_64), .ZN(n_63));
   NAND2_X1 i_56 (.A1(to_int6153[4]), .A2(to_int[2]), .ZN(n_64));
   AOI22_X1 i_57 (.A1(to_int6153[2]), .A2(to_int[2]), .B1(to_int[0]), .B2(
      to_int6153[4]), .ZN(n_65));
   XOR2_X1 i_58 (.A(n_70), .B(n_67), .Z(n_19));
   OAI211_X1 i_59 (.A(to_int6153[1]), .B(to_int[3]), .C1(n_79), .C2(n_119), 
      .ZN(n_67));
   NAND2_X1 i_60 (.A1(to_int6153[0]), .A2(to_int[4]), .ZN(n_70));
   OAI22_X1 i_61 (.A1(n_74), .A2(n_71), .B1(n_73), .B2(n_96), .ZN(n_20));
   NAND2_X1 i_62 (.A1(to_int6153[1]), .A2(to_int[2]), .ZN(n_71));
   NOR2_X1 i_63 (.A1(n_96), .A2(n_73), .ZN(n_72));
   NAND2_X1 i_64 (.A1(to_int6153[3]), .A2(to_int[1]), .ZN(n_73));
   AOI22_X1 i_65 (.A1(to_int6153[2]), .A2(to_int[1]), .B1(to_int[0]), .B2(
      to_int6153[3]), .ZN(n_74));
   NOR2_X1 i_66 (.A1(n_80), .A2(n_75), .ZN(i[1]));
   INV_X1 i_67 (.A(n_79), .ZN(n_75));
   NAND4_X1 i_68 (.A1(to_int6153[1]), .A2(to_int6153[0]), .A3(to_int[1]), 
      .A4(to_int[0]), .ZN(n_79));
   AOI22_X1 i_69 (.A1(to_int6153[0]), .A2(to_int[1]), .B1(to_int[0]), .B2(
      to_int6153[1]), .ZN(n_80));
   NOR3_X1 i_70 (.A1(n_97), .A2(n_85), .A3(n_83), .ZN(i[2]));
   AOI21_X1 i_71 (.A(to_int6153[0]), .B1(n_93), .B2(n_84), .ZN(n_83));
   OR2_X1 i_72 (.A1(n_117), .A2(n_96), .ZN(n_84));
   AOI21_X1 i_73 (.A(n_92), .B1(to_int[0]), .B2(n_119), .ZN(n_85));
   NAND3_X1 i_74 (.A1(n_93), .A2(to_int[2]), .A3(to_int6153[0]), .ZN(n_92));
   NAND2_X1 i_75 (.A1(n_117), .A2(n_96), .ZN(n_93));
   NAND2_X1 i_76 (.A1(to_int6153[2]), .A2(to_int[0]), .ZN(n_96));
   AOI21_X1 i_77 (.A(to_int[2]), .B1(n_103), .B2(n_98), .ZN(n_97));
   NAND2_X1 i_78 (.A1(i[0]), .A2(n_119), .ZN(n_98));
   AND2_X1 i_79 (.A1(to_int6153[0]), .A2(to_int[0]), .ZN(i[0]));
   NAND2_X1 i_80 (.A1(n_118), .A2(n_117), .ZN(n_103));
   NAND2_X1 i_81 (.A1(to_int6153[1]), .A2(to_int[1]), .ZN(n_117));
   INV_X1 i_82 (.A(to_int[0]), .ZN(n_118));
   INV_X1 i_83 (.A(to_int6153[2]), .ZN(n_119));
endmodule

module int_multiplier__4_384(a, b, enbl, c);
   input [15:0]a;
   input [15:0]b;
   input enbl;
   output [15:0]c;

   datapath__4_383 i_0 (.to_int6153({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, uc_0, uc_1, 
      uc_2, uc_3, uc_4, uc_5, b[5], b[4], b[3], b[2], b[1], b[0]}), .to_int({
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, uc_6, uc_7, uc_8, uc_9, uc_10, uc_11, a[5], 
      a[4], a[3], a[2], a[1], a[0]}), .i({uc_12, uc_13, uc_14, uc_15, uc_16, 
      uc_17, uc_18, uc_19, uc_20, uc_21, uc_22, uc_23, uc_24, uc_25, uc_26, 
      uc_27, uc_28, uc_29, uc_30, uc_31, c[11], c[10], c[9], c[8], c[7], c[6], 
      c[5], c[4], c[3], c[2], c[1], c[0]}));
endmodule

module full_adder__4_373(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   INV_X1 i_3 (.A(b), .ZN(f));
endmodule

module full_adder__4_369(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XNOR2_X1 i_0_0 (.A(b), .B(cin), .ZN(f));
   OR2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(cout));
endmodule

module full_adder__4_365(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(b), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(b), .ZN(cout));
endmodule

module full_adder__4_361(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(b), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(b), .ZN(cout));
endmodule

module full_adder__4_357(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(b), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(b), .ZN(cout));
endmodule

module full_adder__4_353(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XNOR2_X1 i_0_0 (.A(b), .B(cin), .ZN(f));
   OR2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(cout));
endmodule

module full_adder__4_349(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XNOR2_X1 i_0_0 (.A(b), .B(cin), .ZN(f));
   OR2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(cout));
endmodule

module full_adder__4_345(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XNOR2_X1 i_0_0 (.A(b), .B(cin), .ZN(f));
   OR2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(cout));
endmodule

module full_adder__4_341(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(b), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(b), .ZN(cout));
endmodule

module full_adder__4_337(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(b), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(b), .ZN(cout));
endmodule

module full_adder__4_333(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XNOR2_X1 i_0_0 (.A(b), .B(cin), .ZN(f));
   OR2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(cout));
endmodule

module int_adder__parameterized3__4_382(a, b, cin, enbl, c, cout);
   input [15:0]a;
   input [15:0]b;
   input cin;
   input enbl;
   output [15:0]c;
   output cout;

   full_adder__4_373 full_adder_0_2_full_adder_0_i (.a(), .b(b[2]), .cin(), 
      .f(c[2]), .cout());
   full_adder__4_369 full_adder_0_3_full_adder_0_i (.a(), .b(b[3]), .cin(b[2]), 
      .f(c[3]), .cout(n_3));
   full_adder__4_365 full_adder_0_4_full_adder_0_i (.a(), .b(b[4]), .cin(n_3), 
      .f(c[4]), .cout(n_4));
   full_adder__4_361 full_adder_0_5_full_adder_0_i (.a(), .b(b[5]), .cin(n_4), 
      .f(c[5]), .cout(n_5));
   full_adder__4_357 full_adder_0_6_full_adder_0_i (.a(), .b(b[6]), .cin(n_5), 
      .f(c[6]), .cout(n_6));
   full_adder__4_353 full_adder_0_7_full_adder_0_i (.a(), .b(b[7]), .cin(n_6), 
      .f(c[7]), .cout(n_7));
   full_adder__4_349 full_adder_0_8_full_adder_0_i (.a(), .b(b[8]), .cin(n_7), 
      .f(c[8]), .cout(n_8));
   full_adder__4_345 full_adder_0_9_full_adder_0_i (.a(), .b(b[9]), .cin(n_8), 
      .f(c[9]), .cout(n_0));
   full_adder__4_341 full_adder_0_10_full_adder_0_i (.a(), .b(b[10]), .cin(n_0), 
      .f(c[10]), .cout(n_1));
   full_adder__4_337 full_adder_0_11_full_adder_0_i (.a(), .b(b[11]), .cin(n_1), 
      .f(c[11]), .cout(n_2));
   full_adder__4_333 full_adder_0_12_full_adder_0_i (.a(), .b(b[12]), .cin(n_2), 
      .f(c[12]), .cout(c[13]));
endmodule

module datapath__0_5915(to_int6153, to_int, i);
   input [16:0]to_int6153;
   input [16:0]to_int;
   output [31:0]i;

   HA_X1 i_164 (.A(n_44), .B(n_38), .CO(n_15), .S(n_14));
   FA_X1 i_179 (.A(n_37), .B(n_36), .CI(n_35), .CO(n_41), .S(n_40));
   HA_X1 i_180 (.A(n_35), .B(n_15), .CO(n_43), .S(n_42));
   FA_X1 i_203 (.A(n_54), .B(n_48), .CI(1'b0), .CO(n_1), .S(n_0));
   HA_X1 i_204 (.A(n_43), .B(n_41), .CO(n_3), .S(n_2));
   FA_X1 i_227 (.A(n_51), .B(n_32), .CI(n_55), .CO(n_5), .S(n_4));
   HA_X1 i_229 (.A(n_4), .B(n_1), .CO(n_7), .S(n_6));
   FA_X1 i_253 (.A(n_31), .B(n_5), .CI(n_7), .CO(n_9), .S(n_8));
   HA_X1 i_254 (.A(n_33), .B(to_int6153[4]), .CO(n_11), .S(n_10));
   HA_X1 i_287 (.A(n_11), .B(n_9), .CO(n_13), .S(n_12));
   FA_X1 i_320 (.A(1'b0), .B(to_int6153[5]), .CI(n_34), .CO(n_17), .S(n_16));
   FA_X1 i_522 (.A(n_29), .B(n_39), .CI(n_28), .CO(n_18), .S(i[3]));
   FA_X1 i_523 (.A(n_27), .B(n_14), .CI(n_18), .CO(n_19), .S(i[4]));
   FA_X1 i_524 (.A(n_42), .B(n_40), .CI(n_19), .CO(n_20), .S(i[5]));
   FA_X1 i_525 (.A(n_2), .B(n_0), .CI(n_20), .CO(n_21), .S(i[6]));
   FA_X1 i_526 (.A(n_3), .B(n_6), .CI(n_21), .CO(n_22), .S(i[7]));
   FA_X1 i_527 (.A(n_8), .B(n_10), .CI(n_22), .CO(n_23), .S(i[8]));
   FA_X1 i_528 (.A(n_12), .B(n_30), .CI(n_23), .CO(n_24), .S(i[9]));
   FA_X1 i_529 (.A(n_13), .B(n_16), .CI(n_24), .CO(n_25), .S(i[10]));
   FA_X1 i_530 (.A(1'b0), .B(n_17), .CI(n_25), .CO(n_26), .S(i[11]));
   XNOR2_X1 i_0 (.A(n_62), .B(n_57), .ZN(n_27));
   AOI21_X1 i_1 (.A(n_64), .B1(n_65), .B2(n_62), .ZN(n_28));
   OAI33_X1 i_2 (.A1(n_64), .A2(n_63), .A3(n_44), .B1(n_64), .B2(n_61), .B3(n_39), 
      .ZN(n_29));
   AND2_X1 i_3 (.A1(to_int6153[5]), .A2(to_int[3]), .ZN(n_30));
   AND2_X1 i_4 (.A1(to_int6153[4]), .A2(to_int[3]), .ZN(n_31));
   OAI21_X1 i_5 (.A(n_46), .B1(n_63), .B2(n_45), .ZN(n_55));
   OAI21_X1 i_6 (.A(n_49), .B1(n_53), .B2(n_52), .ZN(n_32));
   XNOR2_X1 i_7 (.A(n_63), .B(n_48), .ZN(n_54));
   NOR2_X1 i_8 (.A1(n_51), .A2(n_45), .ZN(n_48));
   AOI22_X1 i_9 (.A1(to_int6153[5]), .A2(to_int6153[1]), .B1(to_int6153[4]), 
      .B2(to_int[2]), .ZN(n_45));
   INV_X1 i_10 (.A(n_46), .ZN(n_51));
   NAND2_X1 i_11 (.A1(n_44), .A2(n_34), .ZN(n_46));
   AND2_X1 i_12 (.A1(to_int6153[5]), .A2(to_int[2]), .ZN(n_33));
   AND2_X1 i_13 (.A1(to_int6153[5]), .A2(to_int6153[4]), .ZN(n_34));
   XOR2_X1 i_14 (.A(n_53), .B(n_47), .Z(n_35));
   NAND2_X1 i_15 (.A1(n_50), .A2(n_49), .ZN(n_47));
   NAND3_X1 i_16 (.A1(to_int6153[5]), .A2(to_int6153[0]), .A3(n_59), .ZN(n_49));
   INV_X1 i_17 (.A(n_52), .ZN(n_50));
   AOI21_X1 i_18 (.A(n_59), .B1(to_int6153[5]), .B2(to_int6153[0]), .ZN(n_52));
   NAND2_X1 i_19 (.A1(to_int[3]), .A2(to_int[2]), .ZN(n_53));
   NAND2_X1 i_20 (.A1(n_58), .A2(n_56), .ZN(n_36));
   AOI21_X1 i_21 (.A(n_60), .B1(n_62), .B2(n_58), .ZN(n_37));
   XNOR2_X1 i_22 (.A(n_57), .B(n_56), .ZN(n_38));
   NAND2_X1 i_23 (.A1(n_44), .A2(n_39), .ZN(n_56));
   AOI21_X1 i_24 (.A(n_60), .B1(n_59), .B2(n_39), .ZN(n_57));
   NAND2_X1 i_25 (.A1(n_59), .A2(n_39), .ZN(n_58));
   NOR2_X1 i_26 (.A1(n_64), .A2(n_63), .ZN(n_39));
   AND2_X1 i_27 (.A1(to_int6153[4]), .A2(to_int6153[1]), .ZN(n_59));
   AOI22_X1 i_28 (.A1(to_int6153[4]), .A2(to_int6153[0]), .B1(to_int6153[1]), 
      .B2(to_int[3]), .ZN(n_60));
   INV_X1 i_29 (.A(n_61), .ZN(n_44));
   NAND2_X1 i_30 (.A1(to_int6153[1]), .A2(to_int[2]), .ZN(n_61));
   NOR2_X1 i_31 (.A1(n_65), .A2(to_int6153[0]), .ZN(i[2]));
   INV_X1 i_32 (.A(to_int[2]), .ZN(n_62));
   INV_X1 i_33 (.A(to_int[3]), .ZN(n_63));
   INV_X1 i_34 (.A(to_int6153[0]), .ZN(n_64));
   INV_X1 i_35 (.A(to_int6153[1]), .ZN(n_65));
endmodule

module int_multiplier(a, b, enbl, c);
   input [15:0]a;
   input [15:0]b;
   input enbl;
   output [15:0]c;

   datapath__0_5915 i_0 (.to_int6153({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, uc_0, uc_1, 
      uc_2, uc_3, uc_4, uc_5, a[5], a[4], uc_6, uc_7, a[1], a[0]}), .to_int({
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, 
      uc_14, uc_15, a[3], a[2], uc_16, uc_17}), .i({uc_18, uc_19, uc_20, uc_21, 
      uc_22, uc_23, uc_24, uc_25, uc_26, uc_27, uc_28, uc_29, uc_30, uc_31, 
      uc_32, uc_33, uc_34, uc_35, uc_36, uc_37, c[11], c[10], c[9], c[8], c[7], 
      c[6], c[5], c[4], c[3], c[2], uc_38, uc_39}));
endmodule

module next_adr(in_data, enbl, clk, rst, out_adr, done, state_test);
   input [31:0]in_data;
   input enbl;
   input clk;
   input rst;
   output [15:0]out_adr;
   output done;
   output [3:0]state_test;

   wire [15:0]new_adr;
   wire [15:0]hdr_tsize_m;
   wire [15:0]max_us_adr;
   wire [15:0]max_u0_adr;
   wire [15:0]max_x_adr;
   wire [15:0]hdr_n_m;
   wire [15:0]max_b_adr;
   wire [15:0]hdr_n_square;
   wire [25:20]i;
   wire [18:17]fpu_mode;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_166;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_180;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_190;
   wire n_0_191;
   wire n_0_192;
   wire n_0_193;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_200;
   wire n_0_201;
   wire n_0_202;
   wire n_0_203;
   wire n_0_204;

   int_adder__parameterized2 iterator (.a(out_adr), .b({n_69, fpu_mode[17]}), 
      .cin(), .enbl(), .c(new_adr), .cout());
   int_multiplier__parameterized0 max_us_adr_mul (.a({uc_0, uc_1, uc_2, uc_3, 
      uc_4, uc_5, uc_6, uc_7, uc_8, uc_9, i[25], i[24], i[23], i[22], i[21], 
      i[20]}), .b({n_27, n_28, n_29}), .enbl(), .c({uc_10, uc_11, uc_12, uc_13, 
      uc_14, uc_15, uc_16, hdr_tsize_m[8], hdr_tsize_m[7], hdr_tsize_m[6], 
      hdr_tsize_m[5], hdr_tsize_m[4], hdr_tsize_m[3], hdr_tsize_m[2], 
      hdr_tsize_m[1], hdr_tsize_m[0]}));
   int_adder__parameterized3__4_317 max_us_adr_add (.a(), .b({uc_17, uc_18, 
      uc_19, uc_20, uc_21, uc_22, hdr_tsize_m[8], hdr_tsize_m[7], hdr_tsize_m[6], 
      hdr_tsize_m[5], hdr_tsize_m[4], hdr_tsize_m[3], hdr_tsize_m[2], 
      hdr_tsize_m[1], hdr_tsize_m[0], uc_23}), .cin(), .enbl(), .c({uc_24, uc_25, 
      uc_26, uc_27, uc_28, max_us_adr[10], max_us_adr[9], max_us_adr[8], 
      max_us_adr[7], max_us_adr[6], max_us_adr[5], max_us_adr[4], max_us_adr[3], 
      max_us_adr[2], max_us_adr[1], uc_29}), .cout());
   int_adder__parameterized4__4_449 max_u0_adr_add (.a(), .b({i[24], i[23], 
      i[22], i[21], uc_30, uc_31}), .cin(), .enbl(), .c({uc_32, uc_33, uc_34, 
      uc_35, uc_36, uc_37, uc_38, uc_39, max_u0_adr[7], max_u0_adr[6], 
      max_u0_adr[5], max_u0_adr[4], max_u0_adr[3], max_u0_adr[2], uc_40, uc_41}), 
      .cout());
   int_adder__parameterized4 max_x_adr_add (.a(), .b({n_22, n_23, n_24, n_25, 
      uc_42, uc_43}), .cin(), .enbl(), .c({uc_44, uc_45, uc_46, uc_47, uc_48, 
      uc_49, uc_50, uc_51, uc_52, max_x_adr[6], max_x_adr[5], max_x_adr[4], 
      max_x_adr[3], max_x_adr[2], uc_53, uc_54}), .cout());
   int_multiplier__4_384 max_b_adr_mul (.a({uc_55, uc_56, uc_57, uc_58, uc_59, 
      uc_60, uc_61, uc_62, uc_63, uc_64, n_21, n_22, n_23, n_24, n_25, n_26}), 
      .b({uc_65, uc_66, uc_67, uc_68, uc_69, uc_70, uc_71, uc_72, uc_73, uc_74, 
      i[25], i[24], i[23], i[22], i[21], i[20]}), .enbl(), .c({uc_75, uc_76, 
      uc_77, uc_78, hdr_n_m[11], hdr_n_m[10], hdr_n_m[9], hdr_n_m[8], hdr_n_m[7], 
      hdr_n_m[6], hdr_n_m[5], hdr_n_m[4], hdr_n_m[3], hdr_n_m[2], hdr_n_m[1], 
      hdr_n_m[0]}));
   int_adder__parameterized3__4_382 max_b_adr_add (.a(), .b({uc_79, uc_80, uc_81, 
      hdr_n_m[11], hdr_n_m[10], hdr_n_m[9], hdr_n_m[8], hdr_n_m[7], hdr_n_m[6], 
      hdr_n_m[5], hdr_n_m[4], hdr_n_m[3], hdr_n_m[2], hdr_n_m[1], uc_82, uc_83}), 
      .cin(), .enbl(), .c({uc_84, uc_85, max_b_adr[13], max_b_adr[12], 
      max_b_adr[11], max_b_adr[10], max_b_adr[9], max_b_adr[8], max_b_adr[7], 
      max_b_adr[6], max_b_adr[5], max_b_adr[4], max_b_adr[3], max_b_adr[2], 
      uc_86, uc_87}), .cout());
   int_multiplier max_a_adr_mul (.a({uc_88, uc_89, uc_90, uc_91, uc_92, uc_93, 
      uc_94, uc_95, uc_96, uc_97, n_21, n_22, n_23, n_24, n_25, n_26}), .b(), 
      .enbl(), .c({uc_98, uc_99, uc_100, uc_101, hdr_n_square[11], 
      hdr_n_square[10], hdr_n_square[9], hdr_n_square[8], hdr_n_square[7], 
      hdr_n_square[6], hdr_n_square[5], hdr_n_square[4], hdr_n_square[3], 
      hdr_n_square[2], uc_102, uc_103}));
   DFFR_X1 done_reg (.D(n_68), .RN(n_71), .CK(n_70), .Q(done), .QN());
   DFFS_X1 \cur_adr_reg[15]  (.D(n_67), .SN(n_71), .CK(n_70), .Q(n_0), .QN());
   DFFS_X1 \cur_adr_reg[14]  (.D(n_66), .SN(n_71), .CK(n_70), .Q(n_1), .QN());
   DFFS_X1 \cur_adr_reg[13]  (.D(n_65), .SN(n_71), .CK(n_70), .Q(n_2), .QN());
   DFFS_X1 \cur_adr_reg[12]  (.D(n_64), .SN(n_71), .CK(n_70), .Q(n_3), .QN());
   DFFS_X1 \cur_adr_reg[11]  (.D(n_63), .SN(n_71), .CK(n_70), .Q(n_4), .QN());
   DFFS_X1 \cur_adr_reg[10]  (.D(n_62), .SN(n_71), .CK(n_70), .Q(n_5), .QN());
   DFFS_X1 \cur_adr_reg[9]  (.D(n_61), .SN(n_71), .CK(n_70), .Q(n_6), .QN());
   DFFS_X1 \cur_adr_reg[8]  (.D(n_60), .SN(n_71), .CK(n_70), .Q(n_7), .QN());
   DFFS_X1 \cur_adr_reg[7]  (.D(n_59), .SN(n_71), .CK(n_70), .Q(n_8), .QN());
   DFFS_X1 \cur_adr_reg[6]  (.D(n_58), .SN(n_71), .CK(n_70), .Q(n_9), .QN());
   DFFS_X1 \cur_adr_reg[5]  (.D(n_57), .SN(n_71), .CK(n_70), .Q(n_10), .QN());
   DFFS_X1 \cur_adr_reg[4]  (.D(n_56), .SN(n_71), .CK(n_70), .Q(n_11), .QN());
   DFFS_X1 \cur_adr_reg[3]  (.D(n_55), .SN(n_71), .CK(n_70), .Q(n_12), .QN());
   DFFS_X1 \cur_adr_reg[2]  (.D(n_54), .SN(n_71), .CK(n_70), .Q(n_13), .QN());
   DFFS_X1 \cur_adr_reg[1]  (.D(n_52), .SN(n_71), .CK(n_70), .Q(n_14), .QN());
   DFFS_X1 \cur_adr_reg[0]  (.D(n_51), .SN(n_71), .CK(n_70), .Q(n_15), .QN());
   TBUF_X1 i_5 (.A(n_15), .EN(n_53), .Z(out_adr[0]));
   TBUF_X1 i_7 (.A(n_14), .EN(n_53), .Z(out_adr[1]));
   TBUF_X1 i_9 (.A(n_13), .EN(n_53), .Z(out_adr[2]));
   TBUF_X1 i_11 (.A(n_12), .EN(n_53), .Z(out_adr[3]));
   TBUF_X1 i_13 (.A(n_11), .EN(n_53), .Z(out_adr[4]));
   TBUF_X1 i_15 (.A(n_10), .EN(n_53), .Z(out_adr[5]));
   TBUF_X1 i_17 (.A(n_9), .EN(n_53), .Z(out_adr[6]));
   TBUF_X1 i_19 (.A(n_8), .EN(n_53), .Z(out_adr[7]));
   TBUF_X1 i_21 (.A(n_7), .EN(n_53), .Z(out_adr[8]));
   TBUF_X1 i_23 (.A(n_6), .EN(n_53), .Z(out_adr[9]));
   TBUF_X1 i_25 (.A(n_5), .EN(n_53), .Z(out_adr[10]));
   TBUF_X1 i_27 (.A(n_4), .EN(n_53), .Z(out_adr[11]));
   TBUF_X1 i_29 (.A(n_3), .EN(n_53), .Z(out_adr[12]));
   TBUF_X1 i_31 (.A(n_2), .EN(n_53), .Z(out_adr[13]));
   TBUF_X1 i_33 (.A(n_1), .EN(n_53), .Z(out_adr[14]));
   TBUF_X1 i_35 (.A(n_0), .EN(n_53), .Z(out_adr[15]));
   INV_X1 i_36 (.A(n_16), .ZN(n_53));
   DFFS_X1 i_39 (.D(n_50), .SN(n_71), .CK(n_70), .Q(n_16), .QN());
   DFFR_X1 \state_reg[3]  (.D(n_49), .RN(n_71), .CK(n_70), .Q(n_17), .QN());
   DFFR_X1 \state_reg[2]  (.D(n_48), .RN(n_71), .CK(n_70), .Q(n_18), .QN());
   DFFR_X1 \state_reg[1]  (.D(n_47), .RN(n_71), .CK(n_70), .Q(n_19), .QN());
   DFFR_X1 \state_reg[0]  (.D(n_46), .RN(n_71), .CK(n_70), .Q(n_20), .QN());
   DFF_X1 \header_reg[31]  (.D(n_45), .CK(n_70), .Q(n_21), .QN());
   DFF_X1 \header_reg[30]  (.D(n_44), .CK(n_70), .Q(n_22), .QN());
   DFF_X1 \header_reg[29]  (.D(n_43), .CK(n_70), .Q(n_23), .QN());
   DFF_X1 \header_reg[28]  (.D(n_42), .CK(n_70), .Q(n_24), .QN());
   DFF_X1 \header_reg[27]  (.D(n_41), .CK(n_70), .Q(n_25), .QN());
   DFF_X1 \header_reg[26]  (.D(n_40), .CK(n_70), .Q(n_26), .QN());
   DFF_X1 \header_reg[25]  (.D(n_39), .CK(n_70), .Q(i[25]), .QN());
   DFF_X1 \header_reg[24]  (.D(n_38), .CK(n_70), .Q(i[24]), .QN());
   DFF_X1 \header_reg[23]  (.D(n_37), .CK(n_70), .Q(i[23]), .QN());
   DFF_X1 \header_reg[22]  (.D(n_36), .CK(n_70), .Q(i[22]), .QN());
   DFF_X1 \header_reg[21]  (.D(n_35), .CK(n_70), .Q(i[21]), .QN());
   DFF_X1 \header_reg[20]  (.D(n_34), .CK(n_70), .Q(i[20]), .QN());
   DFF_X1 \header_reg[17]  (.D(n_33), .CK(n_70), .Q(fpu_mode[17]), .QN());
   DFF_X1 \header_reg[16]  (.D(n_32), .CK(n_70), .Q(n_27), .QN());
   DFF_X1 \header_reg[15]  (.D(n_31), .CK(n_70), .Q(n_28), .QN());
   DFF_X1 \header_reg[14]  (.D(n_30), .CK(n_70), .Q(n_29), .QN());
   MUX2_X1 i_0_0 (.A(n_29), .B(in_data[14]), .S(n_0_1), .Z(n_30));
   MUX2_X1 i_0_1 (.A(n_28), .B(in_data[15]), .S(n_0_1), .Z(n_31));
   MUX2_X1 i_0_2 (.A(n_27), .B(in_data[16]), .S(n_0_1), .Z(n_32));
   OAI21_X1 i_0_3 (.A(n_0_0), .B1(n_0_1), .B2(n_69), .ZN(n_33));
   NAND2_X1 i_0_4 (.A1(in_data[17]), .A2(n_0_1), .ZN(n_0_0));
   MUX2_X1 i_0_5 (.A(i[20]), .B(in_data[20]), .S(n_0_1), .Z(n_34));
   MUX2_X1 i_0_6 (.A(i[21]), .B(in_data[21]), .S(n_0_1), .Z(n_35));
   MUX2_X1 i_0_7 (.A(i[22]), .B(in_data[22]), .S(n_0_1), .Z(n_36));
   MUX2_X1 i_0_8 (.A(i[23]), .B(in_data[23]), .S(n_0_1), .Z(n_37));
   MUX2_X1 i_0_9 (.A(i[24]), .B(in_data[24]), .S(n_0_1), .Z(n_38));
   MUX2_X1 i_0_10 (.A(i[25]), .B(in_data[25]), .S(n_0_1), .Z(n_39));
   MUX2_X1 i_0_11 (.A(n_26), .B(in_data[26]), .S(n_0_1), .Z(n_40));
   MUX2_X1 i_0_12 (.A(n_25), .B(in_data[27]), .S(n_0_1), .Z(n_41));
   MUX2_X1 i_0_13 (.A(n_24), .B(in_data[28]), .S(n_0_1), .Z(n_42));
   MUX2_X1 i_0_14 (.A(n_23), .B(in_data[29]), .S(n_0_1), .Z(n_43));
   MUX2_X1 i_0_15 (.A(n_22), .B(in_data[30]), .S(n_0_1), .Z(n_44));
   MUX2_X1 i_0_16 (.A(n_21), .B(in_data[31]), .S(n_0_1), .Z(n_45));
   NOR4_X1 i_0_17 (.A1(n_0_175), .A2(n_0_173), .A3(n_20), .A4(rst), .ZN(n_0_1));
   OAI211_X1 i_0_18 (.A(n_0_10), .B(n_0_8), .C1(n_0_2), .C2(n_20), .ZN(n_46));
   OAI21_X1 i_0_19 (.A(n_0_202), .B1(n_0_75), .B2(n_0_3), .ZN(n_0_2));
   NOR3_X1 i_0_20 (.A1(n_0_5), .A2(n_0_4), .A3(new_adr[13]), .ZN(n_0_3));
   NAND3_X1 i_0_21 (.A1(new_adr[2]), .A2(n_0_164), .A3(n_0_155), .ZN(n_0_4));
   NAND4_X1 i_0_22 (.A1(new_adr[0]), .A2(n_0_196), .A3(n_0_7), .A4(n_0_6), 
      .ZN(n_0_5));
   NOR4_X1 i_0_23 (.A1(new_adr[12]), .A2(new_adr[10]), .A3(new_adr[9]), .A4(
      new_adr[1]), .ZN(n_0_6));
   NOR4_X1 i_0_24 (.A1(new_adr[8]), .A2(new_adr[6]), .A3(new_adr[4]), .A4(n_18), 
      .ZN(n_0_7));
   AOI22_X1 i_0_25 (.A1(n_0_176), .A2(n_0_9), .B1(n_0_76), .B2(n_0_78), .ZN(
      n_0_8));
   OAI22_X1 i_0_26 (.A1(n_0_179), .A2(n_0_174), .B1(n_0_173), .B2(n_20), 
      .ZN(n_0_9));
   OAI21_X1 i_0_27 (.A(n_20), .B1(n_0_11), .B2(n_0_173), .ZN(n_0_10));
   OAI21_X1 i_0_28 (.A(n_0_12), .B1(n_0_143), .B2(n_0_199), .ZN(n_0_11));
   NAND2_X1 i_0_29 (.A1(n_0_24), .A2(n_0_199), .ZN(n_0_12));
   AOI21_X1 i_0_30 (.A(n_0_13), .B1(n_0_16), .B2(n_0_121), .ZN(n_47));
   OAI22_X1 i_0_31 (.A1(n_0_14), .A2(n_0_199), .B1(n_19), .B2(n_0_170), .ZN(
      n_0_13));
   INV_X1 i_0_32 (.A(n_0_15), .ZN(n_0_14));
   OAI21_X1 i_0_33 (.A(n_0_70), .B1(n_0_147), .B2(n_0_203), .ZN(n_0_15));
   NOR3_X1 i_0_34 (.A1(n_0_203), .A2(n_18), .A3(n_0_198), .ZN(n_0_16));
   NAND2_X1 i_0_35 (.A1(n_0_67), .A2(n_0_17), .ZN(n_48));
   OAI21_X1 i_0_36 (.A(n_18), .B1(n_0_148), .B2(n_0_72), .ZN(n_0_17));
   OAI21_X1 i_0_37 (.A(n_0_200), .B1(n_0_147), .B2(n_0_18), .ZN(n_49));
   NAND3_X1 i_0_38 (.A1(n_18), .A2(n_20), .A3(enbl), .ZN(n_0_18));
   AOI21_X1 i_0_39 (.A(n_0_172), .B1(n_0_85), .B2(n_0_197), .ZN(n_50));
   INV_X1 i_0_40 (.A(n_0_19), .ZN(n_51));
   AOI222_X1 i_0_41 (.A1(n_0_23), .A2(n_0_170), .B1(n_15), .B2(n_0_85), .C1(
      n_0_52), .C2(new_adr[0]), .ZN(n_0_19));
   OAI21_X1 i_0_42 (.A(n_0_20), .B1(n_0_147), .B2(n_0_169), .ZN(n_52));
   AOI22_X1 i_0_43 (.A1(n_0_21), .A2(new_adr[1]), .B1(n_14), .B2(n_0_85), 
      .ZN(n_0_20));
   OAI211_X1 i_0_44 (.A(n_0_87), .B(n_0_22), .C1(n_0_23), .C2(n_0_203), .ZN(
      n_0_21));
   AOI21_X1 i_0_45 (.A(n_0_204), .B1(n_0_141), .B2(n_0_131), .ZN(n_0_22));
   OAI21_X1 i_0_46 (.A(n_0_144), .B1(n_0_24), .B2(n_18), .ZN(n_0_23));
   NOR2_X1 i_0_47 (.A1(n_0_121), .A2(n_0_198), .ZN(n_0_24));
   NAND3_X1 i_0_48 (.A1(n_0_53), .A2(n_0_26), .A3(n_0_25), .ZN(n_54));
   AOI21_X1 i_0_49 (.A(n_0_38), .B1(n_0_85), .B2(n_13), .ZN(n_0_25));
   OAI21_X1 i_0_50 (.A(new_adr[2]), .B1(n_0_139), .B2(n_0_27), .ZN(n_0_26));
   OAI211_X1 i_0_51 (.A(n_0_59), .B(n_0_28), .C1(n_19), .C2(n_0_171), .ZN(n_0_27));
   NAND2_X1 i_0_52 (.A1(n_0_90), .A2(n_0_78), .ZN(n_0_28));
   NAND3_X1 i_0_53 (.A1(n_0_50), .A2(n_0_30), .A3(n_0_29), .ZN(n_55));
   NAND2_X1 i_0_54 (.A1(n_12), .A2(n_0_85), .ZN(n_0_29));
   NAND2_X1 i_0_55 (.A1(n_0_31), .A2(new_adr[3]), .ZN(n_0_30));
   NAND3_X1 i_0_56 (.A1(n_0_169), .A2(n_0_88), .A3(n_0_138), .ZN(n_0_31));
   NAND3_X1 i_0_57 (.A1(n_0_74), .A2(n_0_33), .A3(n_0_32), .ZN(n_56));
   AOI21_X1 i_0_58 (.A(n_0_45), .B1(n_0_85), .B2(n_11), .ZN(n_0_32));
   NAND2_X1 i_0_59 (.A1(n_0_34), .A2(new_adr[4]), .ZN(n_0_33));
   NAND3_X1 i_0_60 (.A1(n_0_142), .A2(n_0_36), .A3(n_0_35), .ZN(n_0_34));
   OAI211_X1 i_0_61 (.A(n_19), .B(n_0_202), .C1(n_0_122), .C2(n_18), .ZN(n_0_35));
   NAND3_X1 i_0_62 (.A1(n_0_175), .A2(n_0_37), .A3(n_0_202), .ZN(n_0_36));
   NAND2_X1 i_0_63 (.A1(n_0_49), .A2(n_20), .ZN(n_0_37));
   OAI21_X1 i_0_64 (.A(n_0_39), .B1(n_0_144), .B2(n_0_169), .ZN(n_57));
   NOR2_X1 i_0_65 (.A1(n_0_169), .A2(n_0_144), .ZN(n_0_38));
   AOI22_X1 i_0_66 (.A1(n_0_40), .A2(new_adr[5]), .B1(n_10), .B2(n_0_85), 
      .ZN(n_0_39));
   NAND4_X1 i_0_67 (.A1(n_0_119), .A2(n_0_59), .A3(n_0_42), .A4(n_0_41), 
      .ZN(n_0_40));
   NAND3_X1 i_0_68 (.A1(n_0_90), .A2(n_0_131), .A3(n_19), .ZN(n_0_41));
   OR2_X1 i_0_69 (.A1(n_0_64), .A2(n_19), .ZN(n_0_42));
   NAND3_X1 i_0_70 (.A1(n_0_43), .A2(n_0_62), .A3(n_0_73), .ZN(n_58));
   AOI22_X1 i_0_71 (.A1(n_9), .A2(n_0_85), .B1(n_0_63), .B2(new_adr[6]), 
      .ZN(n_0_43));
   NAND4_X1 i_0_72 (.A1(n_0_67), .A2(n_0_62), .A3(n_0_46), .A4(n_0_44), .ZN(n_59));
   AOI21_X1 i_0_73 (.A(n_0_45), .B1(n_0_85), .B2(n_8), .ZN(n_0_44));
   NOR2_X1 i_0_74 (.A1(n_0_169), .A2(n_0_147), .ZN(n_0_45));
   OAI21_X1 i_0_75 (.A(new_adr[7]), .B1(n_0_47), .B2(n_0_204), .ZN(n_0_46));
   OAI211_X1 i_0_76 (.A(n_0_140), .B(n_0_48), .C1(n_0_49), .C2(n_0_203), 
      .ZN(n_0_47));
   NAND2_X1 i_0_77 (.A1(n_0_94), .A2(n_0_78), .ZN(n_0_48));
   NAND2_X1 i_0_78 (.A1(n_0_151), .A2(n_18), .ZN(n_0_49));
   NAND3_X1 i_0_79 (.A1(n_0_50), .A2(n_0_74), .A3(n_0_51), .ZN(n_60));
   AND2_X1 i_0_80 (.A1(n_0_73), .A2(n_0_67), .ZN(n_0_50));
   AOI22_X1 i_0_81 (.A1(n_0_52), .A2(new_adr[8]), .B1(n_7), .B2(n_0_85), 
      .ZN(n_0_51));
   OAI21_X1 i_0_82 (.A(n_0_142), .B1(n_0_173), .B2(n_0_176), .ZN(n_0_52));
   NAND3_X1 i_0_83 (.A1(n_0_53), .A2(n_0_54), .A3(n_0_55), .ZN(n_61));
   AOI21_X1 i_0_84 (.A(n_0_66), .B1(n_0_75), .B2(n_0_78), .ZN(n_0_53));
   NAND2_X1 i_0_85 (.A1(n_6), .A2(n_0_85), .ZN(n_0_54));
   OAI21_X1 i_0_86 (.A(new_adr[9]), .B1(n_0_71), .B2(n_0_60), .ZN(n_0_55));
   NAND2_X1 i_0_87 (.A1(n_0_57), .A2(n_0_56), .ZN(n_62));
   AOI22_X1 i_0_88 (.A1(n_5), .A2(n_0_85), .B1(n_0_78), .B2(n_0_75), .ZN(n_0_56));
   OAI21_X1 i_0_89 (.A(new_adr[10]), .B1(n_0_60), .B2(n_0_58), .ZN(n_0_57));
   OAI21_X1 i_0_90 (.A(n_0_119), .B1(n_0_59), .B2(n_0_198), .ZN(n_0_58));
   NAND3_X1 i_0_91 (.A1(n_0_148), .A2(n_0_170), .A3(n_18), .ZN(n_0_59));
   OAI22_X1 i_0_92 (.A1(n_0_76), .A2(n_0_77), .B1(n_0_171), .B2(n_0_70), 
      .ZN(n_0_60));
   NAND3_X1 i_0_93 (.A1(n_0_61), .A2(n_0_62), .A3(n_0_73), .ZN(n_63));
   AOI22_X1 i_0_94 (.A1(n_4), .A2(n_0_85), .B1(n_0_63), .B2(new_adr[11]), 
      .ZN(n_0_61));
   NAND2_X1 i_0_95 (.A1(n_0_78), .A2(n_0_76), .ZN(n_0_62));
   NAND3_X1 i_0_96 (.A1(n_0_142), .A2(n_0_82), .A3(n_0_64), .ZN(n_0_63));
   OAI211_X1 i_0_97 (.A(n_18), .B(n_0_202), .C1(n_0_94), .C2(n_20), .ZN(n_0_64));
   NAND2_X1 i_0_98 (.A1(n_0_68), .A2(n_0_65), .ZN(n_64));
   AOI21_X1 i_0_99 (.A(n_0_66), .B1(n_0_85), .B2(n_3), .ZN(n_0_65));
   INV_X1 i_0_100 (.A(n_0_67), .ZN(n_0_66));
   NAND4_X1 i_0_101 (.A1(n_19), .A2(n_0_170), .A3(n_0_121), .A4(n_0_199), 
      .ZN(n_0_67));
   OAI21_X1 i_0_102 (.A(new_adr[12]), .B1(n_0_71), .B2(n_0_69), .ZN(n_0_68));
   OAI21_X1 i_0_103 (.A(n_0_87), .B1(n_0_70), .B2(n_0_169), .ZN(n_0_69));
   NAND2_X1 i_0_104 (.A1(n_0_198), .A2(n_0_151), .ZN(n_0_70));
   OAI21_X1 i_0_105 (.A(n_0_138), .B1(n_0_149), .B2(n_0_72), .ZN(n_0_71));
   NAND2_X1 i_0_106 (.A1(n_19), .A2(n_0_170), .ZN(n_0_72));
   NAND4_X1 i_0_107 (.A1(n_0_80), .A2(n_0_79), .A3(n_0_74), .A4(n_0_73), 
      .ZN(n_65));
   NAND3_X1 i_0_108 (.A1(n_0_143), .A2(n_0_170), .A3(n_18), .ZN(n_0_73));
   OAI21_X1 i_0_109 (.A(n_0_78), .B1(n_0_76), .B2(n_0_75), .ZN(n_0_74));
   NOR2_X1 i_0_110 (.A1(n_0_94), .A2(n_19), .ZN(n_0_75));
   NOR2_X1 i_0_111 (.A1(n_0_198), .A2(n_0_90), .ZN(n_0_76));
   INV_X1 i_0_112 (.A(n_0_78), .ZN(n_0_77));
   NOR2_X1 i_0_113 (.A1(n_0_171), .A2(n_20), .ZN(n_0_78));
   NAND2_X1 i_0_114 (.A1(n_2), .A2(n_0_85), .ZN(n_0_79));
   NAND2_X1 i_0_115 (.A1(n_0_81), .A2(new_adr[13]), .ZN(n_0_80));
   NAND3_X1 i_0_116 (.A1(n_0_171), .A2(n_0_142), .A3(n_0_82), .ZN(n_0_81));
   NAND2_X1 i_0_117 (.A1(n_0_120), .A2(n_19), .ZN(n_0_82));
   INV_X1 i_0_118 (.A(n_0_83), .ZN(n_66));
   AOI22_X1 i_0_119 (.A1(n_0_86), .A2(new_adr[14]), .B1(n_1), .B2(n_0_85), 
      .ZN(n_0_83));
   INV_X1 i_0_120 (.A(n_0_84), .ZN(n_67));
   AOI22_X1 i_0_121 (.A1(n_0_86), .A2(new_adr[15]), .B1(n_0), .B2(n_0_85), 
      .ZN(n_0_84));
   OAI21_X1 i_0_122 (.A(enbl), .B1(n_0_176), .B2(n_0_200), .ZN(n_0_85));
   OAI211_X1 i_0_123 (.A(n_0_119), .B(n_0_87), .C1(n_0_169), .C2(n_0_143), 
      .ZN(n_0_86));
   OR2_X1 i_0_124 (.A1(n_0_88), .A2(n_20), .ZN(n_0_87));
   OR2_X1 i_0_125 (.A1(n_0_173), .A2(n_0_89), .ZN(n_0_88));
   AOI22_X1 i_0_126 (.A1(n_0_94), .A2(n_0_93), .B1(n_0_90), .B2(n_19), .ZN(
      n_0_89));
   NAND4_X1 i_0_127 (.A1(n_0_115), .A2(n_0_92), .A3(n_0_91), .A4(n_0_117), 
      .ZN(n_0_90));
   NOR4_X1 i_0_128 (.A1(n_0_165), .A2(n_0_118), .A3(n_0_116), .A4(n_0_112), 
      .ZN(n_0_91));
   NOR2_X1 i_0_129 (.A1(n_0_114), .A2(n_0_113), .ZN(n_0_92));
   NOR2_X1 i_0_130 (.A1(n_0_199), .A2(n_19), .ZN(n_0_93));
   NAND3_X1 i_0_131 (.A1(n_0_97), .A2(n_0_96), .A3(n_0_95), .ZN(n_0_94));
   NOR4_X1 i_0_132 (.A1(n_0_110), .A2(n_0_108), .A3(n_0_106), .A4(n_0_101), 
      .ZN(n_0_95));
   NOR4_X1 i_0_133 (.A1(n_0_111), .A2(n_0_107), .A3(n_0_103), .A4(n_0_99), 
      .ZN(n_0_96));
   NOR3_X1 i_0_134 (.A1(n_0_195), .A2(n_0_105), .A3(n_0_98), .ZN(n_0_97));
   NAND4_X1 i_0_135 (.A1(n_0_109), .A2(n_0_104), .A3(n_0_102), .A4(n_0_100), 
      .ZN(n_0_98));
   XOR2_X1 i_0_136 (.A(new_adr[4]), .B(max_b_adr[4]), .Z(n_0_99));
   XNOR2_X1 i_0_137 (.A(new_adr[13]), .B(max_b_adr[13]), .ZN(n_0_100));
   XOR2_X1 i_0_138 (.A(new_adr[1]), .B(hdr_n_m[0]), .Z(n_0_101));
   XNOR2_X1 i_0_139 (.A(new_adr[10]), .B(max_b_adr[10]), .ZN(n_0_102));
   XOR2_X1 i_0_140 (.A(new_adr[5]), .B(max_b_adr[5]), .Z(n_0_103));
   XNOR2_X1 i_0_141 (.A(new_adr[8]), .B(max_b_adr[8]), .ZN(n_0_104));
   XOR2_X1 i_0_142 (.A(new_adr[2]), .B(max_b_adr[2]), .Z(n_0_105));
   XOR2_X1 i_0_143 (.A(new_adr[7]), .B(max_b_adr[7]), .Z(n_0_106));
   XOR2_X1 i_0_144 (.A(new_adr[11]), .B(max_b_adr[11]), .Z(n_0_107));
   XOR2_X1 i_0_145 (.A(new_adr[6]), .B(max_b_adr[6]), .Z(n_0_108));
   XNOR2_X1 i_0_146 (.A(new_adr[3]), .B(max_b_adr[3]), .ZN(n_0_109));
   XOR2_X1 i_0_147 (.A(new_adr[9]), .B(max_b_adr[9]), .Z(n_0_110));
   XOR2_X1 i_0_148 (.A(new_adr[12]), .B(max_b_adr[12]), .Z(n_0_111));
   XOR2_X1 i_0_149 (.A(new_adr[2]), .B(max_u0_adr[2]), .Z(n_0_112));
   XOR2_X1 i_0_150 (.A(new_adr[7]), .B(max_u0_adr[7]), .Z(n_0_113));
   XOR2_X1 i_0_151 (.A(new_adr[3]), .B(max_u0_adr[3]), .Z(n_0_114));
   XNOR2_X1 i_0_152 (.A(new_adr[4]), .B(max_u0_adr[4]), .ZN(n_0_115));
   XOR2_X1 i_0_153 (.A(new_adr[6]), .B(max_u0_adr[6]), .Z(n_0_116));
   XNOR2_X1 i_0_154 (.A(new_adr[1]), .B(i[20]), .ZN(n_0_117));
   XOR2_X1 i_0_155 (.A(new_adr[5]), .B(max_u0_adr[5]), .Z(n_0_118));
   AOI21_X1 i_0_156 (.A(n_0_204), .B1(n_0_120), .B2(n_0_141), .ZN(n_0_119));
   AOI21_X1 i_0_157 (.A(n_0_173), .B1(n_0_121), .B2(n_20), .ZN(n_0_120));
   INV_X1 i_0_158 (.A(n_0_122), .ZN(n_0_121));
   NAND3_X1 i_0_159 (.A1(n_0_133), .A2(n_0_129), .A3(n_0_123), .ZN(n_0_122));
   NOR3_X1 i_0_160 (.A1(n_0_157), .A2(n_0_127), .A3(n_0_124), .ZN(n_0_123));
   NAND4_X1 i_0_161 (.A1(n_0_135), .A2(n_0_132), .A3(n_0_126), .A4(n_0_125), 
      .ZN(n_0_124));
   NOR4_X1 i_0_162 (.A1(n_0_136), .A2(n_0_134), .A3(n_0_130), .A4(n_0_128), 
      .ZN(n_0_125));
   XNOR2_X1 i_0_163 (.A(new_adr[9]), .B(hdr_n_square[8]), .ZN(n_0_126));
   NAND4_X1 i_0_164 (.A1(new_adr[2]), .A2(n_0_196), .A3(n_0_137), .A4(n_0_201), 
      .ZN(n_0_127));
   XOR2_X1 i_0_165 (.A(new_adr[11]), .B(hdr_n_square[10]), .Z(n_0_128));
   XNOR2_X1 i_0_166 (.A(new_adr[10]), .B(hdr_n_square[9]), .ZN(n_0_129));
   XOR2_X1 i_0_167 (.A(new_adr[12]), .B(hdr_n_square[11]), .Z(n_0_130));
   NOR2_X1 i_0_168 (.A1(n_0_173), .A2(n_20), .ZN(n_0_131));
   XNOR2_X1 i_0_169 (.A(new_adr[8]), .B(hdr_n_square[7]), .ZN(n_0_132));
   XNOR2_X1 i_0_170 (.A(new_adr[5]), .B(hdr_n_square[4]), .ZN(n_0_133));
   XOR2_X1 i_0_171 (.A(new_adr[6]), .B(hdr_n_square[5]), .Z(n_0_134));
   XNOR2_X1 i_0_172 (.A(new_adr[4]), .B(hdr_n_square[3]), .ZN(n_0_135));
   XOR2_X1 i_0_173 (.A(new_adr[3]), .B(hdr_n_square[2]), .Z(n_0_136));
   XNOR2_X1 i_0_174 (.A(new_adr[7]), .B(hdr_n_square[6]), .ZN(n_0_137));
   INV_X1 i_0_175 (.A(n_0_139), .ZN(n_0_138));
   OAI21_X1 i_0_176 (.A(n_0_142), .B1(n_0_140), .B2(n_18), .ZN(n_0_139));
   NAND2_X1 i_0_177 (.A1(n_19), .A2(n_0_202), .ZN(n_0_140));
   NOR2_X1 i_0_178 (.A1(n_0_198), .A2(n_18), .ZN(n_0_141));
   OR3_X1 i_0_179 (.A1(n_0_175), .A2(n_0_174), .A3(n_20), .ZN(n_0_142));
   NAND2_X1 i_0_180 (.A1(n_0_147), .A2(n_0_144), .ZN(n_0_143));
   OR4_X1 i_0_181 (.A1(n_0_157), .A2(n_0_153), .A3(n_0_145), .A4(n_19), .ZN(
      n_0_144));
   NAND2_X1 i_0_182 (.A1(new_adr[8]), .A2(n_0_146), .ZN(n_0_145));
   NOR2_X1 i_0_183 (.A1(n_0_168), .A2(n_0_152), .ZN(n_0_146));
   NAND2_X1 i_0_184 (.A1(n_19), .A2(n_0_149), .ZN(n_0_147));
   INV_X1 i_0_185 (.A(n_0_149), .ZN(n_0_148));
   NOR4_X1 i_0_186 (.A1(n_0_165), .A2(n_0_163), .A3(n_0_154), .A4(n_0_150), 
      .ZN(n_0_149));
   NAND4_X1 i_0_187 (.A1(new_adr[7]), .A2(new_adr[6]), .A3(new_adr[4]), .A4(
      n_0_164), .ZN(n_0_150));
   OR4_X1 i_0_188 (.A1(n_0_167), .A2(n_0_157), .A3(n_0_153), .A4(n_0_152), 
      .ZN(n_0_151));
   NAND4_X1 i_0_189 (.A1(n_0_159), .A2(n_0_155), .A3(new_adr[10]), .A4(
      new_adr[9]), .ZN(n_0_152));
   NAND4_X1 i_0_190 (.A1(n_0_162), .A2(n_0_161), .A3(n_0_160), .A4(n_0_156), 
      .ZN(n_0_153));
   XOR2_X1 i_0_191 (.A(new_adr[1]), .B(n_29), .Z(n_0_154));
   NOR2_X1 i_0_192 (.A1(new_adr[11]), .A2(new_adr[7]), .ZN(n_0_155));
   XNOR2_X1 i_0_193 (.A(new_adr[4]), .B(max_x_adr[4]), .ZN(n_0_156));
   NAND2_X1 i_0_194 (.A1(n_0_158), .A2(new_adr[0]), .ZN(n_0_157));
   XNOR2_X1 i_0_195 (.A(new_adr[1]), .B(n_26), .ZN(n_0_158));
   XNOR2_X1 i_0_196 (.A(new_adr[6]), .B(max_x_adr[6]), .ZN(n_0_159));
   XNOR2_X1 i_0_197 (.A(new_adr[2]), .B(max_x_adr[2]), .ZN(n_0_160));
   XNOR2_X1 i_0_198 (.A(new_adr[3]), .B(max_x_adr[3]), .ZN(n_0_161));
   XNOR2_X1 i_0_199 (.A(new_adr[5]), .B(max_x_adr[5]), .ZN(n_0_162));
   XOR2_X1 i_0_200 (.A(new_adr[2]), .B(n_28), .Z(n_0_163));
   NOR2_X1 i_0_201 (.A1(new_adr[5]), .A2(new_adr[3]), .ZN(n_0_164));
   OR4_X1 i_0_202 (.A1(n_0_167), .A2(n_0_166), .A3(new_adr[10]), .A4(new_adr[9]), 
      .ZN(n_0_165));
   NAND2_X1 i_0_203 (.A1(new_adr[11]), .A2(new_adr[0]), .ZN(n_0_166));
   NAND3_X1 i_0_204 (.A1(new_adr[8]), .A2(n_0_196), .A3(n_0_190), .ZN(n_0_167));
   NAND2_X1 i_0_205 (.A1(n_0_196), .A2(n_0_190), .ZN(n_0_168));
   NAND2_X1 i_0_206 (.A1(n_18), .A2(n_0_170), .ZN(n_0_169));
   AND2_X1 i_0_207 (.A1(n_20), .A2(n_0_202), .ZN(n_0_170));
   NAND2_X1 i_0_208 (.A1(n_18), .A2(n_0_202), .ZN(n_0_171));
   OR2_X1 i_0_209 (.A1(done), .A2(n_0_172), .ZN(n_68));
   NOR3_X1 i_0_210 (.A1(n_0_177), .A2(n_0_175), .A3(n_0_174), .ZN(n_0_172));
   NAND2_X1 i_0_211 (.A1(n_0_200), .A2(enbl), .ZN(n_0_173));
   NAND2_X1 i_0_212 (.A1(n_17), .A2(enbl), .ZN(n_0_174));
   NAND2_X1 i_0_213 (.A1(n_0_199), .A2(n_0_198), .ZN(n_0_175));
   NOR2_X1 i_0_214 (.A1(n_18), .A2(n_19), .ZN(n_0_176));
   NOR2_X1 i_0_215 (.A1(n_20), .A2(n_0_178), .ZN(n_0_177));
   INV_X1 i_0_216 (.A(n_0_179), .ZN(n_0_178));
   NAND3_X1 i_0_217 (.A1(n_0_186), .A2(n_0_182), .A3(n_0_180), .ZN(n_0_179));
   NOR3_X1 i_0_218 (.A1(n_0_181), .A2(n_0_193), .A3(n_0_191), .ZN(n_0_180));
   NAND3_X1 i_0_219 (.A1(new_adr[11]), .A2(n_0_190), .A3(n_0_189), .ZN(n_0_181));
   NOR4_X1 i_0_220 (.A1(n_0_195), .A2(n_0_185), .A3(n_0_184), .A4(n_0_183), 
      .ZN(n_0_182));
   XOR2_X1 i_0_221 (.A(max_us_adr[6]), .B(new_adr[6]), .Z(n_0_183));
   XOR2_X1 i_0_222 (.A(max_us_adr[2]), .B(new_adr[2]), .Z(n_0_184));
   XOR2_X1 i_0_223 (.A(max_us_adr[10]), .B(new_adr[10]), .Z(n_0_185));
   NOR4_X1 i_0_224 (.A1(n_0_194), .A2(n_0_192), .A3(n_0_188), .A4(n_0_187), 
      .ZN(n_0_186));
   XOR2_X1 i_0_225 (.A(max_us_adr[5]), .B(new_adr[5]), .Z(n_0_187));
   XOR2_X1 i_0_226 (.A(max_us_adr[8]), .B(new_adr[8]), .Z(n_0_188));
   XNOR2_X1 i_0_227 (.A(max_us_adr[1]), .B(new_adr[1]), .ZN(n_0_189));
   NOR2_X1 i_0_228 (.A1(n_0_201), .A2(new_adr[12]), .ZN(n_0_190));
   XOR2_X1 i_0_229 (.A(max_us_adr[4]), .B(new_adr[4]), .Z(n_0_191));
   XOR2_X1 i_0_230 (.A(max_us_adr[7]), .B(new_adr[7]), .Z(n_0_192));
   XOR2_X1 i_0_231 (.A(max_us_adr[9]), .B(new_adr[9]), .Z(n_0_193));
   XOR2_X1 i_0_232 (.A(max_us_adr[3]), .B(new_adr[3]), .Z(n_0_194));
   NAND2_X1 i_0_233 (.A1(new_adr[0]), .A2(n_0_196), .ZN(n_0_195));
   NOR2_X1 i_0_234 (.A1(new_adr[15]), .A2(new_adr[14]), .ZN(n_0_196));
   INV_X1 i_0_235 (.A(fpu_mode[17]), .ZN(n_69));
   INV_X1 i_0_236 (.A(n_16), .ZN(n_0_197));
   INV_X1 i_0_237 (.A(clk), .ZN(n_70));
   INV_X1 i_0_238 (.A(rst), .ZN(n_71));
   INV_X1 i_0_239 (.A(n_19), .ZN(n_0_198));
   INV_X1 i_0_240 (.A(n_18), .ZN(n_0_199));
   INV_X1 i_0_241 (.A(n_17), .ZN(n_0_200));
   INV_X1 i_0_242 (.A(new_adr[13]), .ZN(n_0_201));
   INV_X1 i_0_243 (.A(n_0_173), .ZN(n_0_202));
   INV_X1 i_0_244 (.A(n_0_170), .ZN(n_0_203));
   INV_X1 i_0_245 (.A(n_0_142), .ZN(n_0_204));
endmodule

module io(in_state, clk, rst, cpu_data, in_data, adr, interrupt, error_success);
   input [1:0]in_state;
   input clk;
   input rst;
   inout [31:0]cpu_data;
   inout [31:0]in_data;
   output [15:0]adr;
   output interrupt;
   output error_success;

   wire dcm_error_success;
   wire [31:0]dcm_out_data;
   wire dcm_out_ready;
   wire nau_done;
   wire [15:0]nau_out_adr;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_0_7;
   wire to_std_logic;
   wire n_0_0_13;
   wire n_0_0;
   wire n_0_0_15;
   wire n_0_21;
   wire n_0_0_8;
   wire n_0_1;
   wire n_0_0_9;
   wire n_0_88;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_0_12;
   wire n_0_56;
   wire n_0_0_14;
   wire n_0_57;
   wire n_0_0_17;
   wire n_0_58;
   wire n_0_0_18;
   wire n_0_59;
   wire n_0_0_19;
   wire n_0_60;
   wire n_0_0_20;
   wire n_0_61;
   wire n_0_0_21;
   wire n_0_62;
   wire n_0_0_22;
   wire n_0_63;
   wire n_0_0_23;
   wire n_0_64;
   wire n_0_0_24;
   wire n_0_65;
   wire n_0_0_25;
   wire n_0_66;
   wire n_0_0_26;
   wire n_0_67;
   wire n_0_0_27;
   wire n_0_68;
   wire n_0_0_28;
   wire n_0_69;
   wire n_0_0_29;
   wire n_0_70;
   wire n_0_0_30;
   wire n_0_71;
   wire n_0_0_31;
   wire n_0_72;
   wire n_0_0_32;
   wire n_0_73;
   wire n_0_0_33;
   wire n_0_74;
   wire n_0_0_34;
   wire n_0_75;
   wire n_0_0_35;
   wire n_0_76;
   wire n_0_0_36;
   wire n_0_77;
   wire n_0_0_37;
   wire n_0_78;
   wire n_0_0_38;
   wire n_0_79;
   wire n_0_0_39;
   wire n_0_80;
   wire n_0_0_40;
   wire n_0_81;
   wire n_0_0_41;
   wire n_0_82;
   wire n_0_0_42;
   wire n_0_83;
   wire n_0_0_43;
   wire n_0_84;
   wire n_0_0_44;
   wire n_0_85;
   wire n_0_0_45;
   wire n_0_86;
   wire n_0_0_46;
   wire n_0_87;
   wire n_0_0_47;
   wire n_0_20;
   wire n_0_0_48;
   wire n_0_0_49;
   wire n_0_0_50;
   wire n_0_0_16;
   wire n_0_0_51;

   decompressor decompressor (.in_data(cpu_data), .rst(rst), .enbl_in(
      to_std_logic), .clk(clk), .state_wait(n_0), .out_ready(dcm_out_ready), 
      .out_data(dcm_out_data), .error_success(dcm_error_success), .buf_test());
   next_adr nau (.in_data({dcm_out_data[31], dcm_out_data[30], dcm_out_data[29], 
      dcm_out_data[28], dcm_out_data[27], dcm_out_data[26], dcm_out_data[25], 
      dcm_out_data[24], dcm_out_data[23], dcm_out_data[22], dcm_out_data[21], 
      dcm_out_data[20], uc_0, uc_1, dcm_out_data[17], dcm_out_data[16], 
      dcm_out_data[15], dcm_out_data[14], uc_2, uc_3, uc_4, uc_5, uc_6, uc_7, 
      uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, uc_15}), .enbl(
      dcm_out_ready), .clk(clk), .rst(rst), .out_adr(nau_out_adr), .done(
      nau_done), .state_test());
   DLH_X1 \adr_reg[15]  (.D(nau_out_adr[15]), .G(n_0_20), .Q(n_0_2));
   DLH_X1 \adr_reg[14]  (.D(nau_out_adr[14]), .G(n_0_20), .Q(n_0_3));
   DLH_X1 \adr_reg[13]  (.D(nau_out_adr[13]), .G(n_0_20), .Q(n_0_4));
   DLH_X1 \adr_reg[12]  (.D(nau_out_adr[12]), .G(n_0_20), .Q(n_0_5));
   DLH_X1 \adr_reg[11]  (.D(nau_out_adr[11]), .G(n_0_20), .Q(n_0_6));
   DLH_X1 \adr_reg[10]  (.D(nau_out_adr[10]), .G(n_0_20), .Q(n_0_7));
   DLH_X1 \adr_reg[9]  (.D(nau_out_adr[9]), .G(n_0_20), .Q(n_0_8));
   DLH_X1 \adr_reg[8]  (.D(nau_out_adr[8]), .G(n_0_20), .Q(n_0_9));
   DLH_X1 \adr_reg[7]  (.D(nau_out_adr[7]), .G(n_0_20), .Q(n_0_10));
   DLH_X1 \adr_reg[6]  (.D(nau_out_adr[6]), .G(n_0_20), .Q(n_0_11));
   DLH_X1 \adr_reg[5]  (.D(nau_out_adr[5]), .G(n_0_20), .Q(n_0_12));
   DLH_X1 \adr_reg[4]  (.D(nau_out_adr[4]), .G(n_0_20), .Q(n_0_13));
   DLH_X1 \adr_reg[3]  (.D(nau_out_adr[3]), .G(n_0_20), .Q(n_0_14));
   DLH_X1 \adr_reg[2]  (.D(nau_out_adr[2]), .G(n_0_20), .Q(n_0_15));
   DLH_X1 \adr_reg[1]  (.D(nau_out_adr[1]), .G(n_0_20), .Q(n_0_16));
   DLH_X1 \adr_reg[0]  (.D(nau_out_adr[0]), .G(n_0_20), .Q(n_0_17));
   TBUF_X1 i_0_5 (.A(n_0_17), .EN(n_0_18), .Z(adr[0]));
   TBUF_X1 i_0_7 (.A(n_0_16), .EN(n_0_18), .Z(adr[1]));
   TBUF_X1 i_0_9 (.A(n_0_15), .EN(n_0_18), .Z(adr[2]));
   TBUF_X1 i_0_11 (.A(n_0_14), .EN(n_0_18), .Z(adr[3]));
   TBUF_X1 i_0_13 (.A(n_0_13), .EN(n_0_18), .Z(adr[4]));
   TBUF_X1 i_0_15 (.A(n_0_12), .EN(n_0_18), .Z(adr[5]));
   TBUF_X1 i_0_17 (.A(n_0_11), .EN(n_0_18), .Z(adr[6]));
   TBUF_X1 i_0_19 (.A(n_0_10), .EN(n_0_18), .Z(adr[7]));
   TBUF_X1 i_0_21 (.A(n_0_9), .EN(n_0_18), .Z(adr[8]));
   TBUF_X1 i_0_23 (.A(n_0_8), .EN(n_0_18), .Z(adr[9]));
   TBUF_X1 i_0_25 (.A(n_0_7), .EN(n_0_18), .Z(adr[10]));
   TBUF_X1 i_0_27 (.A(n_0_6), .EN(n_0_18), .Z(adr[11]));
   TBUF_X1 i_0_29 (.A(n_0_5), .EN(n_0_18), .Z(adr[12]));
   TBUF_X1 i_0_31 (.A(n_0_4), .EN(n_0_18), .Z(adr[13]));
   TBUF_X1 i_0_33 (.A(n_0_3), .EN(n_0_18), .Z(adr[14]));
   TBUF_X1 i_0_35 (.A(n_0_2), .EN(n_0_18), .Z(adr[15]));
   INV_X1 i_0_36 (.A(n_0_19), .ZN(n_0_18));
   DLH_X1 i_0_37 (.D(n_0_21), .G(n_0_20), .Q(n_0_19));
   DLH_X1 \cpu_data_reg[31]  (.D(n_0_87), .G(n_0_88), .Q(n_0_22));
   DLH_X1 \cpu_data_reg[30]  (.D(n_0_86), .G(n_0_88), .Q(n_0_23));
   DLH_X1 \cpu_data_reg[29]  (.D(n_0_85), .G(n_0_88), .Q(n_0_24));
   DLH_X1 \cpu_data_reg[28]  (.D(n_0_84), .G(n_0_88), .Q(n_0_25));
   DLH_X1 \cpu_data_reg[27]  (.D(n_0_83), .G(n_0_88), .Q(n_0_26));
   DLH_X1 \cpu_data_reg[26]  (.D(n_0_82), .G(n_0_88), .Q(n_0_27));
   DLH_X1 \cpu_data_reg[25]  (.D(n_0_81), .G(n_0_88), .Q(n_0_28));
   DLH_X1 \cpu_data_reg[24]  (.D(n_0_80), .G(n_0_88), .Q(n_0_29));
   DLH_X1 \cpu_data_reg[23]  (.D(n_0_79), .G(n_0_88), .Q(n_0_30));
   DLH_X1 \cpu_data_reg[22]  (.D(n_0_78), .G(n_0_88), .Q(n_0_31));
   DLH_X1 \cpu_data_reg[21]  (.D(n_0_77), .G(n_0_88), .Q(n_0_32));
   DLH_X1 \cpu_data_reg[20]  (.D(n_0_76), .G(n_0_88), .Q(n_0_33));
   DLH_X1 \cpu_data_reg[19]  (.D(n_0_75), .G(n_0_88), .Q(n_0_34));
   DLH_X1 \cpu_data_reg[18]  (.D(n_0_74), .G(n_0_88), .Q(n_0_35));
   DLH_X1 \cpu_data_reg[17]  (.D(n_0_73), .G(n_0_88), .Q(n_0_36));
   DLH_X1 \cpu_data_reg[16]  (.D(n_0_72), .G(n_0_88), .Q(n_0_37));
   DLH_X1 \cpu_data_reg[15]  (.D(n_0_71), .G(n_0_88), .Q(n_0_38));
   DLH_X1 \cpu_data_reg[14]  (.D(n_0_70), .G(n_0_88), .Q(n_0_39));
   DLH_X1 \cpu_data_reg[13]  (.D(n_0_69), .G(n_0_88), .Q(n_0_40));
   DLH_X1 \cpu_data_reg[12]  (.D(n_0_68), .G(n_0_88), .Q(n_0_41));
   DLH_X1 \cpu_data_reg[11]  (.D(n_0_67), .G(n_0_88), .Q(n_0_42));
   DLH_X1 \cpu_data_reg[10]  (.D(n_0_66), .G(n_0_88), .Q(n_0_43));
   DLH_X1 \cpu_data_reg[9]  (.D(n_0_65), .G(n_0_88), .Q(n_0_44));
   DLH_X1 \cpu_data_reg[8]  (.D(n_0_64), .G(n_0_88), .Q(n_0_45));
   DLH_X1 \cpu_data_reg[7]  (.D(n_0_63), .G(n_0_88), .Q(n_0_46));
   DLH_X1 \cpu_data_reg[6]  (.D(n_0_62), .G(n_0_88), .Q(n_0_47));
   DLH_X1 \cpu_data_reg[5]  (.D(n_0_61), .G(n_0_88), .Q(n_0_48));
   DLH_X1 \cpu_data_reg[4]  (.D(n_0_60), .G(n_0_88), .Q(n_0_49));
   DLH_X1 \cpu_data_reg[3]  (.D(n_0_59), .G(n_0_88), .Q(n_0_50));
   DLH_X1 \cpu_data_reg[2]  (.D(n_0_58), .G(n_0_88), .Q(n_0_51));
   DLH_X1 \cpu_data_reg[1]  (.D(n_0_57), .G(n_0_88), .Q(n_0_52));
   DLH_X1 \cpu_data_reg[0]  (.D(n_0_56), .G(n_0_88), .Q(n_0_53));
   TBUF_X1 i_0_55 (.A(n_0_53), .EN(n_0_54), .Z(cpu_data[0]));
   TBUF_X1 i_0_57 (.A(n_0_52), .EN(n_0_54), .Z(cpu_data[1]));
   TBUF_X1 i_0_59 (.A(n_0_51), .EN(n_0_54), .Z(cpu_data[2]));
   TBUF_X1 i_0_61 (.A(n_0_50), .EN(n_0_54), .Z(cpu_data[3]));
   TBUF_X1 i_0_63 (.A(n_0_49), .EN(n_0_54), .Z(cpu_data[4]));
   TBUF_X1 i_0_65 (.A(n_0_48), .EN(n_0_54), .Z(cpu_data[5]));
   TBUF_X1 i_0_67 (.A(n_0_47), .EN(n_0_54), .Z(cpu_data[6]));
   TBUF_X1 i_0_69 (.A(n_0_46), .EN(n_0_54), .Z(cpu_data[7]));
   TBUF_X1 i_0_71 (.A(n_0_45), .EN(n_0_54), .Z(cpu_data[8]));
   TBUF_X1 i_0_73 (.A(n_0_44), .EN(n_0_54), .Z(cpu_data[9]));
   TBUF_X1 i_0_75 (.A(n_0_43), .EN(n_0_54), .Z(cpu_data[10]));
   TBUF_X1 i_0_77 (.A(n_0_42), .EN(n_0_54), .Z(cpu_data[11]));
   TBUF_X1 i_0_79 (.A(n_0_41), .EN(n_0_54), .Z(cpu_data[12]));
   TBUF_X1 i_0_81 (.A(n_0_40), .EN(n_0_54), .Z(cpu_data[13]));
   TBUF_X1 i_0_83 (.A(n_0_39), .EN(n_0_54), .Z(cpu_data[14]));
   TBUF_X1 i_0_85 (.A(n_0_38), .EN(n_0_54), .Z(cpu_data[15]));
   TBUF_X1 i_0_87 (.A(n_0_37), .EN(n_0_54), .Z(cpu_data[16]));
   TBUF_X1 i_0_89 (.A(n_0_36), .EN(n_0_54), .Z(cpu_data[17]));
   TBUF_X1 i_0_91 (.A(n_0_35), .EN(n_0_54), .Z(cpu_data[18]));
   TBUF_X1 i_0_93 (.A(n_0_34), .EN(n_0_54), .Z(cpu_data[19]));
   TBUF_X1 i_0_95 (.A(n_0_33), .EN(n_0_54), .Z(cpu_data[20]));
   TBUF_X1 i_0_97 (.A(n_0_32), .EN(n_0_54), .Z(cpu_data[21]));
   TBUF_X1 i_0_99 (.A(n_0_31), .EN(n_0_54), .Z(cpu_data[22]));
   TBUF_X1 i_0_101 (.A(n_0_30), .EN(n_0_54), .Z(cpu_data[23]));
   TBUF_X1 i_0_103 (.A(n_0_29), .EN(n_0_54), .Z(cpu_data[24]));
   TBUF_X1 i_0_105 (.A(n_0_28), .EN(n_0_54), .Z(cpu_data[25]));
   TBUF_X1 i_0_107 (.A(n_0_27), .EN(n_0_54), .Z(cpu_data[26]));
   TBUF_X1 i_0_109 (.A(n_0_26), .EN(n_0_54), .Z(cpu_data[27]));
   TBUF_X1 i_0_111 (.A(n_0_25), .EN(n_0_54), .Z(cpu_data[28]));
   TBUF_X1 i_0_113 (.A(n_0_24), .EN(n_0_54), .Z(cpu_data[29]));
   TBUF_X1 i_0_115 (.A(n_0_23), .EN(n_0_54), .Z(cpu_data[30]));
   TBUF_X1 i_0_117 (.A(n_0_22), .EN(n_0_54), .Z(cpu_data[31]));
   INV_X1 i_0_118 (.A(n_0_55), .ZN(n_0_54));
   DLH_X1 i_0_119 (.D(n_0_1), .G(n_0_88), .Q(n_0_55));
   DFF_X1 \in_data_reg[31]  (.D(dcm_out_data[31]), .CK(n_0_0), .Q(in_data[31]), 
      .QN());
   DFF_X1 \in_data_reg[30]  (.D(dcm_out_data[30]), .CK(n_0_0), .Q(in_data[30]), 
      .QN());
   DFF_X1 \in_data_reg[29]  (.D(dcm_out_data[29]), .CK(n_0_0), .Q(in_data[29]), 
      .QN());
   DFF_X1 \in_data_reg[28]  (.D(dcm_out_data[28]), .CK(n_0_0), .Q(in_data[28]), 
      .QN());
   DFF_X1 \in_data_reg[27]  (.D(dcm_out_data[27]), .CK(n_0_0), .Q(in_data[27]), 
      .QN());
   DFF_X1 \in_data_reg[26]  (.D(dcm_out_data[26]), .CK(n_0_0), .Q(in_data[26]), 
      .QN());
   DFF_X1 \in_data_reg[25]  (.D(dcm_out_data[25]), .CK(n_0_0), .Q(in_data[25]), 
      .QN());
   DFF_X1 \in_data_reg[24]  (.D(dcm_out_data[24]), .CK(n_0_0), .Q(in_data[24]), 
      .QN());
   DFF_X1 \in_data_reg[23]  (.D(dcm_out_data[23]), .CK(n_0_0), .Q(in_data[23]), 
      .QN());
   DFF_X1 \in_data_reg[22]  (.D(dcm_out_data[22]), .CK(n_0_0), .Q(in_data[22]), 
      .QN());
   DFF_X1 \in_data_reg[21]  (.D(dcm_out_data[21]), .CK(n_0_0), .Q(in_data[21]), 
      .QN());
   DFF_X1 \in_data_reg[20]  (.D(dcm_out_data[20]), .CK(n_0_0), .Q(in_data[20]), 
      .QN());
   DFF_X1 \in_data_reg[19]  (.D(dcm_out_data[19]), .CK(n_0_0), .Q(in_data[19]), 
      .QN());
   DFF_X1 \in_data_reg[18]  (.D(dcm_out_data[18]), .CK(n_0_0), .Q(in_data[18]), 
      .QN());
   DFF_X1 \in_data_reg[17]  (.D(dcm_out_data[17]), .CK(n_0_0), .Q(in_data[17]), 
      .QN());
   DFF_X1 \in_data_reg[16]  (.D(dcm_out_data[16]), .CK(n_0_0), .Q(in_data[16]), 
      .QN());
   DFF_X1 \in_data_reg[15]  (.D(dcm_out_data[15]), .CK(n_0_0), .Q(in_data[15]), 
      .QN());
   DFF_X1 \in_data_reg[14]  (.D(dcm_out_data[14]), .CK(n_0_0), .Q(in_data[14]), 
      .QN());
   DFF_X1 \in_data_reg[13]  (.D(dcm_out_data[13]), .CK(n_0_0), .Q(in_data[13]), 
      .QN());
   DFF_X1 \in_data_reg[12]  (.D(dcm_out_data[12]), .CK(n_0_0), .Q(in_data[12]), 
      .QN());
   DFF_X1 \in_data_reg[11]  (.D(dcm_out_data[11]), .CK(n_0_0), .Q(in_data[11]), 
      .QN());
   DFF_X1 \in_data_reg[10]  (.D(dcm_out_data[10]), .CK(n_0_0), .Q(in_data[10]), 
      .QN());
   DFF_X1 \in_data_reg[9]  (.D(dcm_out_data[9]), .CK(n_0_0), .Q(in_data[9]), 
      .QN());
   DFF_X1 \in_data_reg[8]  (.D(dcm_out_data[8]), .CK(n_0_0), .Q(in_data[8]), 
      .QN());
   DFF_X1 \in_data_reg[7]  (.D(dcm_out_data[7]), .CK(n_0_0), .Q(in_data[7]), 
      .QN());
   DFF_X1 \in_data_reg[6]  (.D(dcm_out_data[6]), .CK(n_0_0), .Q(in_data[6]), 
      .QN());
   DFF_X1 \in_data_reg[5]  (.D(dcm_out_data[5]), .CK(n_0_0), .Q(in_data[5]), 
      .QN());
   DFF_X1 \in_data_reg[4]  (.D(dcm_out_data[4]), .CK(n_0_0), .Q(in_data[4]), 
      .QN());
   DFF_X1 \in_data_reg[3]  (.D(dcm_out_data[3]), .CK(n_0_0), .Q(in_data[3]), 
      .QN());
   DFF_X1 \in_data_reg[2]  (.D(dcm_out_data[2]), .CK(n_0_0), .Q(in_data[2]), 
      .QN());
   DFF_X1 \in_data_reg[1]  (.D(dcm_out_data[1]), .CK(n_0_0), .Q(in_data[1]), 
      .QN());
   DFF_X1 \in_data_reg[0]  (.D(dcm_out_data[0]), .CK(n_0_0), .Q(in_data[0]), 
      .QN());
   MUX2_X1 i_0_0_0 (.A(to_std_logic), .B(n_0), .S(n_0_0_0), .Z(n_0_0_0));
   MUX2_X1 i_0_0_1 (.A(to_std_logic), .B(n_0), .S(n_0_0_1), .Z(n_0_0_1));
   MUX2_X1 i_0_0_2 (.A(to_std_logic), .B(n_0), .S(n_0_0_2), .Z(n_0_0_2));
   MUX2_X1 i_0_0_3 (.A(to_std_logic), .B(n_0), .S(n_0_0_3), .Z(n_0_0_3));
   MUX2_X1 i_0_0_4 (.A(to_std_logic), .B(n_0), .S(n_0_0_4), .Z(n_0_0_4));
   MUX2_X1 i_0_0_5 (.A(to_std_logic), .B(n_0), .S(n_0_0_5), .Z(n_0_0_5));
   MUX2_X1 i_0_0_6 (.A(to_std_logic), .B(n_0), .S(n_0_0_6), .Z(n_0_0_6));
   MUX2_X1 i_0_0_7 (.A(to_std_logic), .B(n_0), .S(n_0_0_7), .Z(n_0_0_7));
   NOR2_X1 i_0_0_8 (.A1(n_0_0_15), .A2(in_state[1]), .ZN(n_0));
   NOR2_X1 i_0_0_9 (.A1(in_state[1]), .A2(in_state[0]), .ZN(to_std_logic));
   OAI211_X1 i_0_0_52 (.A(rst), .B(n_0_0_13), .C1(n_0_0_8), .C2(in_state[1]), 
      .ZN(error_success));
   AOI21_X1 i_0_0_53 (.A(n_0_0_6), .B1(n_0_0_7), .B2(in_state[1]), .ZN(n_0_0_13));
   INV_X1 i_0_0_54 (.A(clk), .ZN(n_0_0));
   INV_X1 i_0_0_10 (.A(in_state[0]), .ZN(n_0_0_15));
   NOR2_X1 i_0_0_11 (.A1(in_state[1]), .A2(n_0_0_50), .ZN(n_0_21));
   INV_X1 i_0_0_12 (.A(dcm_error_success), .ZN(n_0_0_8));
   INV_X1 i_0_0_15 (.A(n_0_0_9), .ZN(n_0_1));
   NAND2_X1 i_0_0_16 (.A1(rst), .A2(n_0_0_0), .ZN(n_0_0_9));
   OAI211_X1 i_0_0_17 (.A(in_state[1]), .B(n_0_0_10), .C1(in_state[0]), .C2(
      n_0_0_11), .ZN(n_0_88));
   NAND2_X1 i_0_0_18 (.A1(rst), .A2(n_0_0_1), .ZN(n_0_0_10));
   INV_X1 i_0_0_19 (.A(n_0_0_12), .ZN(n_0_0_11));
   OR2_X1 i_0_0_20 (.A1(n_0_0_50), .A2(n_0_0_2), .ZN(n_0_0_12));
   INV_X1 i_0_0_21 (.A(n_0_0_14), .ZN(n_0_56));
   NAND2_X1 i_0_0_22 (.A1(in_data[0]), .A2(n_0_0_3), .ZN(n_0_0_14));
   INV_X1 i_0_0_23 (.A(n_0_0_17), .ZN(n_0_57));
   NAND2_X1 i_0_0_24 (.A1(in_data[1]), .A2(n_0_0_3), .ZN(n_0_0_17));
   INV_X1 i_0_0_25 (.A(n_0_0_18), .ZN(n_0_58));
   NAND2_X1 i_0_0_26 (.A1(in_data[2]), .A2(n_0_0_3), .ZN(n_0_0_18));
   INV_X1 i_0_0_27 (.A(n_0_0_19), .ZN(n_0_59));
   NAND2_X1 i_0_0_28 (.A1(in_data[3]), .A2(n_0_0_3), .ZN(n_0_0_19));
   INV_X1 i_0_0_29 (.A(n_0_0_20), .ZN(n_0_60));
   NAND2_X1 i_0_0_30 (.A1(in_data[4]), .A2(n_0_0_3), .ZN(n_0_0_20));
   INV_X1 i_0_0_31 (.A(n_0_0_21), .ZN(n_0_61));
   NAND2_X1 i_0_0_32 (.A1(in_data[5]), .A2(n_0_0_3), .ZN(n_0_0_21));
   INV_X1 i_0_0_33 (.A(n_0_0_22), .ZN(n_0_62));
   NAND2_X1 i_0_0_34 (.A1(in_data[6]), .A2(n_0_0_3), .ZN(n_0_0_22));
   INV_X1 i_0_0_35 (.A(n_0_0_23), .ZN(n_0_63));
   NAND2_X1 i_0_0_36 (.A1(in_data[7]), .A2(n_0_0_3), .ZN(n_0_0_23));
   INV_X1 i_0_0_37 (.A(n_0_0_24), .ZN(n_0_64));
   NAND2_X1 i_0_0_38 (.A1(in_data[8]), .A2(n_0_0_3), .ZN(n_0_0_24));
   INV_X1 i_0_0_39 (.A(n_0_0_25), .ZN(n_0_65));
   NAND2_X1 i_0_0_40 (.A1(in_data[9]), .A2(n_0_0_3), .ZN(n_0_0_25));
   INV_X1 i_0_0_41 (.A(n_0_0_26), .ZN(n_0_66));
   NAND2_X1 i_0_0_42 (.A1(in_data[10]), .A2(n_0_0_3), .ZN(n_0_0_26));
   INV_X1 i_0_0_43 (.A(n_0_0_27), .ZN(n_0_67));
   NAND2_X1 i_0_0_44 (.A1(in_data[11]), .A2(n_0_0_3), .ZN(n_0_0_27));
   INV_X1 i_0_0_45 (.A(n_0_0_28), .ZN(n_0_68));
   NAND2_X1 i_0_0_46 (.A1(in_data[12]), .A2(n_0_0_3), .ZN(n_0_0_28));
   INV_X1 i_0_0_47 (.A(n_0_0_29), .ZN(n_0_69));
   NAND2_X1 i_0_0_48 (.A1(in_data[13]), .A2(n_0_0_3), .ZN(n_0_0_29));
   INV_X1 i_0_0_49 (.A(n_0_0_30), .ZN(n_0_70));
   NAND2_X1 i_0_0_50 (.A1(in_data[14]), .A2(n_0_0_3), .ZN(n_0_0_30));
   INV_X1 i_0_0_51 (.A(n_0_0_31), .ZN(n_0_71));
   NAND2_X1 i_0_0_55 (.A1(in_data[15]), .A2(n_0_0_3), .ZN(n_0_0_31));
   INV_X1 i_0_0_56 (.A(n_0_0_32), .ZN(n_0_72));
   NAND2_X1 i_0_0_57 (.A1(in_data[16]), .A2(n_0_0_3), .ZN(n_0_0_32));
   INV_X1 i_0_0_58 (.A(n_0_0_33), .ZN(n_0_73));
   NAND2_X1 i_0_0_59 (.A1(in_data[17]), .A2(n_0_0_3), .ZN(n_0_0_33));
   INV_X1 i_0_0_60 (.A(n_0_0_34), .ZN(n_0_74));
   NAND2_X1 i_0_0_61 (.A1(in_data[18]), .A2(n_0_0_3), .ZN(n_0_0_34));
   INV_X1 i_0_0_62 (.A(n_0_0_35), .ZN(n_0_75));
   NAND2_X1 i_0_0_63 (.A1(in_data[19]), .A2(n_0_0_3), .ZN(n_0_0_35));
   INV_X1 i_0_0_64 (.A(n_0_0_36), .ZN(n_0_76));
   NAND2_X1 i_0_0_65 (.A1(in_data[20]), .A2(n_0_0_3), .ZN(n_0_0_36));
   INV_X1 i_0_0_66 (.A(n_0_0_37), .ZN(n_0_77));
   NAND2_X1 i_0_0_67 (.A1(in_data[21]), .A2(n_0_0_3), .ZN(n_0_0_37));
   INV_X1 i_0_0_68 (.A(n_0_0_38), .ZN(n_0_78));
   NAND2_X1 i_0_0_69 (.A1(in_data[22]), .A2(n_0_0_3), .ZN(n_0_0_38));
   INV_X1 i_0_0_70 (.A(n_0_0_39), .ZN(n_0_79));
   NAND2_X1 i_0_0_71 (.A1(in_data[23]), .A2(n_0_0_3), .ZN(n_0_0_39));
   INV_X1 i_0_0_72 (.A(n_0_0_40), .ZN(n_0_80));
   NAND2_X1 i_0_0_73 (.A1(in_data[24]), .A2(n_0_0_3), .ZN(n_0_0_40));
   INV_X1 i_0_0_74 (.A(n_0_0_41), .ZN(n_0_81));
   NAND2_X1 i_0_0_75 (.A1(in_data[25]), .A2(n_0_0_3), .ZN(n_0_0_41));
   INV_X1 i_0_0_76 (.A(n_0_0_42), .ZN(n_0_82));
   NAND2_X1 i_0_0_77 (.A1(in_data[26]), .A2(n_0_0_3), .ZN(n_0_0_42));
   INV_X1 i_0_0_78 (.A(n_0_0_43), .ZN(n_0_83));
   NAND2_X1 i_0_0_79 (.A1(in_data[27]), .A2(n_0_0_3), .ZN(n_0_0_43));
   INV_X1 i_0_0_80 (.A(n_0_0_44), .ZN(n_0_84));
   NAND2_X1 i_0_0_81 (.A1(in_data[28]), .A2(n_0_0_3), .ZN(n_0_0_44));
   INV_X1 i_0_0_82 (.A(n_0_0_45), .ZN(n_0_85));
   NAND2_X1 i_0_0_83 (.A1(in_data[29]), .A2(n_0_0_3), .ZN(n_0_0_45));
   INV_X1 i_0_0_84 (.A(n_0_0_46), .ZN(n_0_86));
   NAND2_X1 i_0_0_85 (.A1(in_data[30]), .A2(n_0_0_3), .ZN(n_0_0_46));
   INV_X1 i_0_0_86 (.A(n_0_0_47), .ZN(n_0_87));
   NAND2_X1 i_0_0_87 (.A1(in_data[31]), .A2(n_0_0_3), .ZN(n_0_0_47));
   OAI21_X1 i_0_0_88 (.A(n_0_0_48), .B1(in_state[1]), .B2(n_0_0_50), .ZN(n_0_20));
   NAND2_X1 i_0_0_89 (.A1(in_state[1]), .A2(n_0_0_49), .ZN(n_0_0_48));
   OR3_X1 i_0_0_90 (.A1(n_0_0_50), .A2(n_0_0_4), .A3(n_0_0_5), .ZN(n_0_0_49));
   INV_X1 i_0_0_91 (.A(rst), .ZN(n_0_0_50));
   NAND2_X1 i_0_0_13 (.A1(n_0_0_8), .A2(rst), .ZN(n_0_0_16));
   NAND2_X1 i_0_0_14 (.A1(nau_done), .A2(rst), .ZN(n_0_0_51));
   AOI21_X1 i_0_0_92 (.A(in_state[1]), .B1(n_0_0_16), .B2(n_0_0_51), .ZN(
      interrupt));
endmodule
