library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
use work.common.all;

-----------------------------------------------------------------ENTITY-----------------------------------------------------------------------------------
entity interp is
    generic (
        WORD_LENGTH : integer := 32;
        ADDR_LENGTH : integer := 16;
        MAX_LENGTH  : integer := 64
    );

    port (
        in_state       : in std_logic_vector(1 downto 0); --state signal sent from CPU
        clk            : in std_logic;
        rst            : in std_logic;
        adr            : in std_logic_vector(15 downto 0);
        in_data        : inout std_logic_vector(31 downto 0);
        interp_done_op : out std_logic_vector(1 downto 0);
        interrupt      : out std_logic;
        error_success  : out std_logic
    );
end entity;

-----------------------------------------------------------------ARCHITECTURE-----------------------------------------------------------------------------------
architecture rtl of interp is
-----------------------------------------------------------------SIGNALS-----------------------------------------------------------------------------------
begin
-----------------------------------------------------------------PORT MAPS-----------------------------------------------------------------------------------
-----------------------------------------------------------------PROCESSES-----------------------------------------------------------------------------------
-----------------------------------------------------------------RESET-----------------------------------------------------------------------------------
-----------------------------------------------------------------INITIALIZATION-----------------------------------------------------------------------------------
-----------------------------------------------------------------ERROR HANDLING-----------------------------------------------------------------------------------
-----------------------------------------------------------------MEMORY IO-----------------------------------------------------------------------------------
-----------------------------------------------------------------MATRIX MANIPULATION-----------------------------------------------------------------------------------
-----------------------------------------------------------------UTILITIES-----------------------------------------------------------------------------------
-----------------------------------------------------------------MAIN FSM-----------------------------------------------------------------------------------
end architecture;