/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Thu Apr 23 20:29:01 2020
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 1840813067 */

module datapath(plus, in_b);
   output [63:0]plus;
   input [63:0]in_b;

   XOR2_X1 i_0 (.A(in_b[1]), .B(in_b[0]), .Z(plus[1]));
   AND2_X1 i_1 (.A1(n_61), .A2(n_0), .ZN(plus[2]));
   OAI21_X1 i_2 (.A(in_b[2]), .B1(in_b[1]), .B2(in_b[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(in_b[3]), .B(n_61), .Z(plus[3]));
   XOR2_X1 i_4 (.A(in_b[4]), .B(n_60), .Z(plus[4]));
   XOR2_X1 i_5 (.A(in_b[5]), .B(n_59), .Z(plus[5]));
   AND2_X1 i_6 (.A1(n_58), .A2(n_1), .ZN(plus[6]));
   OAI21_X1 i_7 (.A(in_b[6]), .B1(n_59), .B2(in_b[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(in_b[7]), .B(n_58), .Z(plus[7]));
   XOR2_X1 i_9 (.A(in_b[8]), .B(n_57), .Z(plus[8]));
   AND2_X1 i_10 (.A1(n_56), .A2(n_2), .ZN(plus[9]));
   OAI21_X1 i_11 (.A(in_b[9]), .B1(n_57), .B2(in_b[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(in_b[10]), .B(n_56), .Z(plus[10]));
   XNOR2_X1 i_13 (.A(in_b[11]), .B(n_55), .ZN(plus[11]));
   XOR2_X1 i_14 (.A(in_b[12]), .B(n_54), .Z(plus[12]));
   XNOR2_X1 i_15 (.A(in_b[13]), .B(n_53), .ZN(plus[13]));
   XOR2_X1 i_16 (.A(in_b[14]), .B(n_52), .Z(plus[14]));
   AND2_X1 i_17 (.A1(n_51), .A2(n_3), .ZN(plus[15]));
   OAI21_X1 i_18 (.A(in_b[15]), .B1(n_52), .B2(in_b[14]), .ZN(n_3));
   XOR2_X1 i_19 (.A(in_b[16]), .B(n_51), .Z(plus[16]));
   XOR2_X1 i_20 (.A(in_b[17]), .B(n_50), .Z(plus[17]));
   XOR2_X1 i_21 (.A(in_b[18]), .B(n_49), .Z(plus[18]));
   XNOR2_X1 i_22 (.A(in_b[19]), .B(n_48), .ZN(plus[19]));
   XNOR2_X1 i_23 (.A(in_b[20]), .B(n_47), .ZN(plus[20]));
   XNOR2_X1 i_24 (.A(in_b[21]), .B(n_46), .ZN(plus[21]));
   XOR2_X1 i_25 (.A(in_b[22]), .B(n_45), .Z(plus[22]));
   XOR2_X1 i_26 (.A(in_b[23]), .B(n_44), .Z(plus[23]));
   XNOR2_X1 i_27 (.A(in_b[24]), .B(n_43), .ZN(plus[24]));
   XNOR2_X1 i_28 (.A(in_b[25]), .B(n_42), .ZN(plus[25]));
   XNOR2_X1 i_29 (.A(in_b[26]), .B(n_41), .ZN(plus[26]));
   XOR2_X1 i_30 (.A(in_b[27]), .B(n_40), .Z(plus[27]));
   XOR2_X1 i_31 (.A(in_b[28]), .B(n_39), .Z(plus[28]));
   XNOR2_X1 i_32 (.A(in_b[29]), .B(n_38), .ZN(plus[29]));
   XNOR2_X1 i_33 (.A(in_b[30]), .B(n_37), .ZN(plus[30]));
   XNOR2_X1 i_34 (.A(in_b[31]), .B(n_36), .ZN(plus[31]));
   XOR2_X1 i_35 (.A(in_b[32]), .B(n_35), .Z(plus[32]));
   XOR2_X1 i_36 (.A(in_b[33]), .B(n_34), .Z(plus[33]));
   XNOR2_X1 i_37 (.A(in_b[34]), .B(n_33), .ZN(plus[34]));
   XNOR2_X1 i_38 (.A(in_b[35]), .B(n_32), .ZN(plus[35]));
   XNOR2_X1 i_39 (.A(in_b[36]), .B(n_31), .ZN(plus[36]));
   XOR2_X1 i_40 (.A(in_b[37]), .B(n_30), .Z(plus[37]));
   XOR2_X1 i_41 (.A(in_b[38]), .B(n_29), .Z(plus[38]));
   XNOR2_X1 i_42 (.A(in_b[39]), .B(n_28), .ZN(plus[39]));
   XNOR2_X1 i_43 (.A(in_b[40]), .B(n_27), .ZN(plus[40]));
   XOR2_X1 i_44 (.A(in_b[41]), .B(n_26), .Z(plus[41]));
   XNOR2_X1 i_45 (.A(in_b[42]), .B(n_25), .ZN(plus[42]));
   XOR2_X1 i_46 (.A(in_b[43]), .B(n_24), .Z(plus[43]));
   AND2_X1 i_47 (.A1(n_23), .A2(n_4), .ZN(plus[44]));
   OAI21_X1 i_48 (.A(in_b[44]), .B1(n_24), .B2(in_b[43]), .ZN(n_4));
   XOR2_X1 i_49 (.A(in_b[45]), .B(n_23), .Z(plus[45]));
   XOR2_X1 i_50 (.A(in_b[46]), .B(n_22), .Z(plus[46]));
   XOR2_X1 i_51 (.A(in_b[47]), .B(n_21), .Z(plus[47]));
   XOR2_X1 i_52 (.A(in_b[48]), .B(n_20), .Z(plus[48]));
   XNOR2_X1 i_53 (.A(in_b[49]), .B(n_19), .ZN(plus[49]));
   XNOR2_X1 i_54 (.A(in_b[50]), .B(n_18), .ZN(plus[50]));
   XNOR2_X1 i_55 (.A(in_b[51]), .B(n_17), .ZN(plus[51]));
   XOR2_X1 i_56 (.A(in_b[52]), .B(n_16), .Z(plus[52]));
   XNOR2_X1 i_57 (.A(in_b[53]), .B(n_15), .ZN(plus[53]));
   XNOR2_X1 i_58 (.A(in_b[54]), .B(n_14), .ZN(plus[54]));
   XNOR2_X1 i_59 (.A(in_b[55]), .B(n_13), .ZN(plus[55]));
   XOR2_X1 i_60 (.A(in_b[56]), .B(n_12), .Z(plus[56]));
   AND2_X1 i_61 (.A1(n_11), .A2(n_5), .ZN(plus[57]));
   OAI21_X1 i_62 (.A(in_b[57]), .B1(n_12), .B2(in_b[56]), .ZN(n_5));
   XOR2_X1 i_63 (.A(in_b[58]), .B(n_11), .Z(plus[58]));
   XNOR2_X1 i_64 (.A(in_b[59]), .B(n_10), .ZN(plus[59]));
   XNOR2_X1 i_65 (.A(in_b[60]), .B(n_9), .ZN(plus[60]));
   XOR2_X1 i_66 (.A(in_b[61]), .B(n_8), .Z(plus[61]));
   XNOR2_X1 i_67 (.A(in_b[62]), .B(n_7), .ZN(plus[62]));
   XNOR2_X1 i_68 (.A(in_b[63]), .B(n_6), .ZN(plus[63]));
   NOR3_X1 i_69 (.A1(n_8), .A2(in_b[61]), .A3(in_b[62]), .ZN(n_6));
   NOR2_X1 i_70 (.A1(n_8), .A2(in_b[61]), .ZN(n_7));
   NAND2_X1 i_71 (.A1(n_9), .A2(n_72), .ZN(n_8));
   NOR3_X1 i_72 (.A1(n_11), .A2(in_b[58]), .A3(in_b[59]), .ZN(n_9));
   NOR2_X1 i_73 (.A1(n_11), .A2(in_b[58]), .ZN(n_10));
   OR3_X1 i_74 (.A1(n_12), .A2(in_b[56]), .A3(in_b[57]), .ZN(n_11));
   NAND2_X1 i_75 (.A1(n_13), .A2(n_71), .ZN(n_12));
   NOR4_X1 i_76 (.A1(n_16), .A2(in_b[52]), .A3(in_b[53]), .A4(in_b[54]), 
      .ZN(n_13));
   NOR3_X1 i_77 (.A1(n_16), .A2(in_b[52]), .A3(in_b[53]), .ZN(n_14));
   NOR2_X1 i_78 (.A1(n_16), .A2(in_b[52]), .ZN(n_15));
   NAND2_X1 i_79 (.A1(n_17), .A2(n_70), .ZN(n_16));
   NOR4_X1 i_80 (.A1(n_20), .A2(in_b[48]), .A3(in_b[49]), .A4(in_b[50]), 
      .ZN(n_17));
   NOR3_X1 i_81 (.A1(n_20), .A2(in_b[48]), .A3(in_b[49]), .ZN(n_18));
   NOR2_X1 i_82 (.A1(n_20), .A2(in_b[48]), .ZN(n_19));
   OR2_X1 i_83 (.A1(n_21), .A2(in_b[47]), .ZN(n_20));
   OR2_X1 i_84 (.A1(n_22), .A2(in_b[46]), .ZN(n_21));
   OR2_X1 i_85 (.A1(n_23), .A2(in_b[45]), .ZN(n_22));
   OR3_X1 i_86 (.A1(n_24), .A2(in_b[43]), .A3(in_b[44]), .ZN(n_23));
   NAND2_X1 i_87 (.A1(n_25), .A2(n_69), .ZN(n_24));
   NOR2_X1 i_88 (.A1(n_26), .A2(in_b[41]), .ZN(n_25));
   NAND2_X1 i_89 (.A1(n_27), .A2(n_68), .ZN(n_26));
   NOR3_X1 i_90 (.A1(n_29), .A2(in_b[38]), .A3(in_b[39]), .ZN(n_27));
   NOR2_X1 i_91 (.A1(n_29), .A2(in_b[38]), .ZN(n_28));
   OR2_X1 i_92 (.A1(n_30), .A2(in_b[37]), .ZN(n_29));
   NAND2_X1 i_93 (.A1(n_31), .A2(n_67), .ZN(n_30));
   NOR4_X1 i_94 (.A1(n_34), .A2(in_b[33]), .A3(in_b[34]), .A4(in_b[35]), 
      .ZN(n_31));
   NOR3_X1 i_95 (.A1(n_34), .A2(in_b[33]), .A3(in_b[34]), .ZN(n_32));
   NOR2_X1 i_96 (.A1(n_34), .A2(in_b[33]), .ZN(n_33));
   OR2_X1 i_97 (.A1(n_35), .A2(in_b[32]), .ZN(n_34));
   NAND2_X1 i_98 (.A1(n_36), .A2(n_66), .ZN(n_35));
   NOR4_X1 i_99 (.A1(n_39), .A2(in_b[28]), .A3(in_b[29]), .A4(in_b[30]), 
      .ZN(n_36));
   NOR3_X1 i_100 (.A1(n_39), .A2(in_b[28]), .A3(in_b[29]), .ZN(n_37));
   NOR2_X1 i_101 (.A1(n_39), .A2(in_b[28]), .ZN(n_38));
   OR2_X1 i_102 (.A1(n_40), .A2(in_b[27]), .ZN(n_39));
   NAND2_X1 i_103 (.A1(n_41), .A2(n_65), .ZN(n_40));
   NOR4_X1 i_104 (.A1(n_44), .A2(in_b[23]), .A3(in_b[24]), .A4(in_b[25]), 
      .ZN(n_41));
   NOR3_X1 i_105 (.A1(n_44), .A2(in_b[23]), .A3(in_b[24]), .ZN(n_42));
   NOR2_X1 i_106 (.A1(n_44), .A2(in_b[23]), .ZN(n_43));
   OR2_X1 i_107 (.A1(n_45), .A2(in_b[22]), .ZN(n_44));
   NAND2_X1 i_108 (.A1(n_46), .A2(n_64), .ZN(n_45));
   NOR4_X1 i_109 (.A1(n_49), .A2(in_b[18]), .A3(in_b[19]), .A4(in_b[20]), 
      .ZN(n_46));
   NOR3_X1 i_110 (.A1(n_49), .A2(in_b[18]), .A3(in_b[19]), .ZN(n_47));
   NOR2_X1 i_111 (.A1(n_49), .A2(in_b[18]), .ZN(n_48));
   OR2_X1 i_112 (.A1(n_50), .A2(in_b[17]), .ZN(n_49));
   OR2_X1 i_113 (.A1(n_51), .A2(in_b[16]), .ZN(n_50));
   OR3_X1 i_114 (.A1(n_52), .A2(in_b[14]), .A3(in_b[15]), .ZN(n_51));
   NAND2_X1 i_115 (.A1(n_53), .A2(n_63), .ZN(n_52));
   NOR2_X1 i_116 (.A1(n_54), .A2(in_b[12]), .ZN(n_53));
   NAND2_X1 i_117 (.A1(n_55), .A2(n_62), .ZN(n_54));
   NOR2_X1 i_118 (.A1(n_56), .A2(in_b[10]), .ZN(n_55));
   OR3_X1 i_119 (.A1(n_57), .A2(in_b[8]), .A3(in_b[9]), .ZN(n_56));
   OR2_X1 i_120 (.A1(n_58), .A2(in_b[7]), .ZN(n_57));
   OR3_X1 i_121 (.A1(n_59), .A2(in_b[5]), .A3(in_b[6]), .ZN(n_58));
   OR2_X1 i_122 (.A1(n_60), .A2(in_b[4]), .ZN(n_59));
   OR2_X1 i_123 (.A1(n_61), .A2(in_b[3]), .ZN(n_60));
   OR3_X1 i_124 (.A1(in_b[2]), .A2(in_b[1]), .A3(in_b[0]), .ZN(n_61));
   INV_X1 i_125 (.A(in_b[11]), .ZN(n_62));
   INV_X1 i_126 (.A(in_b[13]), .ZN(n_63));
   INV_X1 i_127 (.A(in_b[21]), .ZN(n_64));
   INV_X1 i_128 (.A(in_b[26]), .ZN(n_65));
   INV_X1 i_129 (.A(in_b[31]), .ZN(n_66));
   INV_X1 i_130 (.A(in_b[36]), .ZN(n_67));
   INV_X1 i_131 (.A(in_b[40]), .ZN(n_68));
   INV_X1 i_132 (.A(in_b[42]), .ZN(n_69));
   INV_X1 i_133 (.A(in_b[51]), .ZN(n_70));
   INV_X1 i_134 (.A(in_b[55]), .ZN(n_71));
   INV_X1 i_135 (.A(in_b[60]), .ZN(n_72));
endmodule

module fpu_adder(mode, clk, rst, enbl, add_sub, in_a, in_b, out_c, done, err, 
      zero, posv);
   input [1:0]mode;
   input clk;
   input rst;
   input enbl;
   input add_sub;
   input [63:0]in_a;
   input [63:0]in_b;
   output [63:0]out_c;
   output done;
   output err;
   output zero;
   output posv;

   wire in_b_signal;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire b;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_1_0;
   wire n_0_1_1;
   wire n_0_1_2;
   wire n_0_125;
   wire n_0_1_3;
   wire n_0_126;
   wire n_0_1_4;
   wire n_0_127;
   wire n_0_1_5;
   wire n_0_128;
   wire n_0_1_6;
   wire n_0_129;
   wire n_0_1_7;
   wire n_0_130;
   wire n_0_1_8;
   wire n_0_131;
   wire n_0_1_9;
   wire n_0_132;
   wire n_0_1_10;
   wire n_0_133;
   wire n_0_1_11;
   wire n_0_134;
   wire n_0_1_12;
   wire n_0_135;
   wire n_0_1_13;
   wire n_0_136;
   wire n_0_1_14;
   wire n_0_137;
   wire n_0_1_15;
   wire n_0_138;
   wire n_0_1_16;
   wire n_0_139;
   wire n_0_1_17;
   wire n_0_140;
   wire n_0_1_18;
   wire n_0_141;
   wire n_0_1_19;
   wire n_0_142;
   wire n_0_1_20;
   wire n_0_143;
   wire n_0_1_21;
   wire n_0_144;
   wire n_0_1_22;
   wire n_0_145;
   wire n_0_1_23;
   wire n_0_146;
   wire n_0_1_24;
   wire n_0_147;
   wire n_0_1_25;
   wire n_0_148;
   wire n_0_1_26;
   wire n_0_149;
   wire n_0_1_27;
   wire n_0_150;
   wire n_0_1_28;
   wire n_0_151;
   wire n_0_1_29;
   wire n_0_152;
   wire n_0_1_30;
   wire n_0_153;
   wire n_0_1_31;
   wire n_0_154;
   wire n_0_1_32;
   wire n_0_155;
   wire n_0_1_33;
   wire n_0_156;
   wire n_0_1_34;
   wire n_0_157;
   wire n_0_1_35;
   wire n_0_158;
   wire n_0_1_36;
   wire n_0_159;
   wire n_0_1_37;
   wire n_0_160;
   wire n_0_1_38;
   wire n_0_161;
   wire n_0_1_39;
   wire n_0_162;
   wire n_0_1_40;
   wire n_0_163;
   wire n_0_1_41;
   wire n_0_164;
   wire n_0_1_42;
   wire n_0_165;
   wire n_0_1_43;
   wire n_0_166;
   wire n_0_1_44;
   wire n_0_167;
   wire n_0_1_45;
   wire n_0_168;
   wire n_0_1_46;
   wire n_0_169;
   wire n_0_1_47;
   wire n_0_170;
   wire n_0_1_48;
   wire n_0_171;
   wire n_0_1_49;
   wire n_0_172;
   wire n_0_1_50;
   wire n_0_173;
   wire n_0_1_51;
   wire n_0_174;
   wire n_0_1_52;
   wire n_0_175;
   wire n_0_1_53;
   wire n_0_176;
   wire n_0_1_54;
   wire n_0_177;
   wire n_0_1_55;
   wire n_0_178;
   wire n_0_1_56;
   wire n_0_179;
   wire n_0_1_57;
   wire n_0_180;
   wire n_0_1_58;
   wire n_0_181;
   wire n_0_1_59;
   wire n_0_182;
   wire n_0_1_60;
   wire n_0_183;
   wire n_0_1_61;
   wire n_0_184;
   wire n_0_1_62;
   wire n_0_185;
   wire n_0_1_63;
   wire n_0_186;
   wire n_0_1_64;
   wire n_0_187;
   wire n_0_1_65;
   wire n_0_188;
   wire n_0_1_66;
   wire n_0_1_67;
   wire n_0_189;
   wire n_0_1_68;
   wire n_0_1_69;
   wire n_0_1_70;
   wire n_0_1_71;
   wire n_0_1_72;
   wire n_0_1_73;
   wire n_0_1_74;
   wire n_0_1_75;
   wire n_0_1_76;
   wire n_0_1_77;
   wire n_0_1_78;
   wire n_0_1_79;
   wire n_0_1_80;
   wire n_0_1_81;
   wire n_0_1_82;
   wire n_0_1_83;
   wire n_0_1_84;
   wire n_0_1_85;
   wire n_0_1_86;
   wire n_0_1_87;
   wire n_0_1_88;
   wire n_0_190;
   wire n_0_191;
   wire n_0_1_89;
   wire n_0_1_90;
   wire n_0_1_91;
   wire n_0_1_92;
   wire FA1_n_0;
   wire n_0_1_93;
   wire n_0_1_94;
   wire n_0_192;
   wire n_0_1_95;
   wire n_0_1_96;
   wire n_0_1_97;
   wire n_0_193;
   wire n_0_1_98;
   wire n_0_1_99;
   wire n_0_1_100;
   wire n_0_1_101;
   wire n_0_1_102;
   wire n_0_194;
   wire n_0_1_103;
   wire n_0_1_104;
   wire n_0_1_105;
   wire n_0_195;
   wire n_0_1_106;
   wire n_0_1_107;
   wire n_0_1_108;
   wire n_0_1_109;
   wire n_0_1_110;
   wire n_0_196;
   wire n_0_1_111;
   wire n_0_1_112;
   wire n_0_1_113;
   wire n_0_197;
   wire n_0_1_114;
   wire n_0_1_115;
   wire n_0_1_116;
   wire n_0_1_117;
   wire n_0_1_118;
   wire n_0_198;
   wire n_0_1_119;
   wire n_0_1_120;
   wire n_0_1_121;
   wire n_0_199;
   wire n_0_1_122;
   wire n_0_1_123;
   wire n_0_1_124;
   wire n_0_1_125;
   wire n_0_1_126;
   wire n_0_200;
   wire n_0_1_127;
   wire n_0_1_128;
   wire n_0_1_129;
   wire n_0_201;
   wire n_0_1_130;
   wire n_0_1_131;
   wire n_0_1_132;
   wire n_0_1_133;
   wire n_0_1_134;
   wire n_0_202;
   wire n_0_1_135;
   wire n_0_1_136;
   wire n_0_1_137;
   wire n_0_203;
   wire n_0_1_138;
   wire n_0_1_139;
   wire n_0_1_140;
   wire n_0_1_141;
   wire n_0_1_142;
   wire n_0_204;
   wire n_0_1_143;
   wire n_0_1_144;
   wire n_0_1_145;
   wire n_0_205;
   wire n_0_1_146;
   wire n_0_1_147;
   wire n_0_1_148;
   wire n_0_1_149;
   wire n_0_1_150;
   wire n_0_206;
   wire n_0_1_151;
   wire n_0_1_152;
   wire n_0_1_153;
   wire n_0_207;
   wire n_0_1_154;
   wire n_0_1_155;
   wire n_0_1_156;
   wire n_0_1_157;
   wire n_0_1_158;
   wire n_0_208;
   wire n_0_1_159;
   wire n_0_1_160;
   wire n_0_1_161;
   wire n_0_209;
   wire n_0_1_162;
   wire n_0_1_163;
   wire n_0_1_164;
   wire n_0_1_165;
   wire n_0_1_166;
   wire n_0_210;
   wire n_0_1_167;
   wire n_0_1_168;
   wire n_0_1_169;
   wire n_0_211;
   wire n_0_1_170;
   wire n_0_1_171;
   wire n_0_1_172;
   wire n_0_1_173;
   wire n_0_1_174;
   wire n_0_212;
   wire n_0_1_175;
   wire n_0_1_176;
   wire n_0_1_177;
   wire n_0_213;
   wire n_0_1_178;
   wire n_0_1_179;
   wire n_0_1_180;
   wire n_0_1_181;
   wire n_0_1_182;
   wire n_0_214;
   wire n_0_1_183;
   wire n_0_1_184;
   wire n_0_1_185;
   wire n_0_215;
   wire n_0_1_186;
   wire n_0_1_187;
   wire n_0_1_188;
   wire n_0_1_189;
   wire n_0_1_190;
   wire n_0_216;
   wire n_0_1_191;
   wire n_0_1_192;
   wire n_0_1_193;
   wire n_0_217;
   wire n_0_1_194;
   wire n_0_1_195;
   wire n_0_1_196;
   wire n_0_1_197;
   wire n_0_1_198;
   wire n_0_218;
   wire n_0_1_199;
   wire n_0_1_200;
   wire n_0_1_201;
   wire n_0_219;
   wire n_0_1_202;
   wire n_0_1_203;
   wire n_0_1_204;
   wire n_0_1_205;
   wire n_0_1_206;
   wire n_0_220;
   wire n_0_1_207;
   wire n_0_1_208;
   wire n_0_1_209;
   wire n_0_221;
   wire n_0_1_210;
   wire n_0_1_211;
   wire n_0_1_212;
   wire n_0_1_213;
   wire n_0_1_214;
   wire n_0_222;
   wire n_0_1_215;
   wire n_0_1_216;
   wire n_0_1_217;
   wire n_0_223;
   wire n_0_1_218;
   wire n_0_1_219;
   wire n_0_1_220;
   wire n_0_1_221;
   wire n_0_1_222;
   wire n_0_224;
   wire n_0_1_223;
   wire n_0_1_224;
   wire n_0_1_225;
   wire n_0_225;
   wire n_0_1_226;
   wire n_0_1_227;
   wire n_0_1_228;
   wire n_0_1_229;
   wire n_0_1_230;
   wire n_0_226;
   wire n_0_1_231;
   wire n_0_1_232;
   wire n_0_1_233;
   wire n_0_227;
   wire n_0_1_234;
   wire n_0_1_235;
   wire n_0_1_236;
   wire n_0_1_237;
   wire n_0_1_238;
   wire n_0_228;
   wire n_0_1_239;
   wire n_0_1_240;
   wire n_0_1_241;
   wire n_0_229;
   wire n_0_1_242;
   wire n_0_1_243;
   wire n_0_1_244;
   wire n_0_1_245;
   wire n_0_1_246;
   wire n_0_230;
   wire n_0_1_247;
   wire n_0_1_248;
   wire n_0_1_249;
   wire n_0_231;
   wire n_0_1_250;
   wire n_0_1_251;
   wire n_0_1_252;
   wire n_0_1_253;
   wire n_0_1_254;
   wire n_0_232;
   wire n_0_1_255;
   wire n_0_1_256;
   wire n_0_1_257;
   wire n_0_233;
   wire n_0_1_258;
   wire n_0_1_259;
   wire n_0_1_260;
   wire n_0_1_261;
   wire n_0_1_262;
   wire n_0_234;
   wire n_0_1_263;
   wire n_0_1_264;
   wire n_0_1_265;
   wire n_0_235;
   wire n_0_1_266;
   wire n_0_1_267;
   wire n_0_1_268;
   wire n_0_1_269;
   wire n_0_1_270;
   wire n_0_236;
   wire n_0_1_271;
   wire n_0_1_272;
   wire n_0_1_273;
   wire n_0_237;
   wire n_0_1_274;
   wire n_0_1_275;
   wire n_0_1_276;
   wire n_0_1_277;
   wire n_0_1_278;
   wire n_0_238;
   wire n_0_1_279;
   wire n_0_1_280;
   wire n_0_1_281;
   wire n_0_239;
   wire n_0_1_282;
   wire n_0_1_283;
   wire n_0_1_284;
   wire n_0_1_285;
   wire n_0_1_286;
   wire n_0_240;
   wire n_0_1_287;
   wire n_0_1_288;
   wire n_0_1_289;
   wire n_0_241;
   wire n_0_1_290;
   wire n_0_1_291;
   wire n_0_1_292;
   wire n_0_1_293;
   wire n_0_1_294;
   wire n_0_242;
   wire n_0_1_295;
   wire n_0_1_296;
   wire n_0_1_297;
   wire n_0_243;
   wire n_0_1_298;
   wire n_0_1_299;
   wire n_0_1_300;
   wire n_0_1_301;
   wire n_0_1_302;
   wire n_0_244;
   wire n_0_1_303;
   wire n_0_1_304;
   wire n_0_1_305;
   wire n_0_245;
   wire n_0_1_306;
   wire n_0_1_307;
   wire n_0_1_308;
   wire n_0_1_309;
   wire n_0_1_310;
   wire n_0_246;
   wire n_0_1_311;
   wire n_0_1_312;
   wire n_0_1_313;
   wire n_0_247;
   wire n_0_1_314;
   wire n_0_1_315;
   wire n_0_1_316;
   wire n_0_1_317;
   wire n_0_1_318;
   wire n_0_248;
   wire n_0_1_319;
   wire n_0_1_320;
   wire n_0_1_321;
   wire n_0_249;
   wire n_0_1_322;
   wire n_0_1_323;
   wire n_0_1_324;
   wire n_0_1_325;
   wire n_0_1_326;
   wire n_0_250;
   wire n_0_1_327;
   wire n_0_1_328;
   wire n_0_1_329;
   wire n_0_251;
   wire n_0_1_330;
   wire n_0_1_331;
   wire n_0_1_332;
   wire n_0_1_333;
   wire n_0_1_334;
   wire n_0_252;
   wire n_0_1_335;
   wire n_0_1_336;
   wire n_0_1_337;
   wire n_0_253;
   wire n_0_1_338;
   wire n_0_1_339;
   wire n_0_1_340;
   wire n_0_254;
   wire n_0_255;

   DLH_X1 posv_reg (.D(n_0_191), .G(n_0_255), .Q(posv));
   DLH_X1 zero_signal_reg (.D(n_0_190), .G(n_0_255), .Q(zero));
   DLH_X1 error_signal_reg (.D(n_0_189), .G(n_0_255), .Q(err));
   DLH_X1 \out_c_signal_reg[63]  (.D(n_0_254), .G(n_0_188), .Q(out_c[63]));
   DLH_X1 \out_c_signal_reg[62]  (.D(n_0_253), .G(n_0_188), .Q(out_c[62]));
   DLH_X1 \out_c_signal_reg[61]  (.D(n_0_252), .G(n_0_188), .Q(out_c[61]));
   DLH_X1 \out_c_signal_reg[60]  (.D(n_0_251), .G(n_0_188), .Q(out_c[60]));
   DLH_X1 \out_c_signal_reg[59]  (.D(n_0_250), .G(n_0_188), .Q(out_c[59]));
   DLH_X1 \out_c_signal_reg[58]  (.D(n_0_249), .G(n_0_188), .Q(out_c[58]));
   DLH_X1 \out_c_signal_reg[57]  (.D(n_0_248), .G(n_0_188), .Q(out_c[57]));
   DLH_X1 \out_c_signal_reg[56]  (.D(n_0_247), .G(n_0_188), .Q(out_c[56]));
   DLH_X1 \out_c_signal_reg[55]  (.D(n_0_246), .G(n_0_188), .Q(out_c[55]));
   DLH_X1 \out_c_signal_reg[54]  (.D(n_0_245), .G(n_0_188), .Q(out_c[54]));
   DLH_X1 \out_c_signal_reg[53]  (.D(n_0_244), .G(n_0_188), .Q(out_c[53]));
   DLH_X1 \out_c_signal_reg[52]  (.D(n_0_243), .G(n_0_188), .Q(out_c[52]));
   DLH_X1 \out_c_signal_reg[51]  (.D(n_0_242), .G(n_0_188), .Q(out_c[51]));
   DLH_X1 \out_c_signal_reg[50]  (.D(n_0_241), .G(n_0_188), .Q(out_c[50]));
   DLH_X1 \out_c_signal_reg[49]  (.D(n_0_240), .G(n_0_188), .Q(out_c[49]));
   DLH_X1 \out_c_signal_reg[48]  (.D(n_0_239), .G(n_0_188), .Q(out_c[48]));
   DLH_X1 \out_c_signal_reg[47]  (.D(n_0_238), .G(n_0_188), .Q(out_c[47]));
   DLH_X1 \out_c_signal_reg[46]  (.D(n_0_237), .G(n_0_188), .Q(out_c[46]));
   DLH_X1 \out_c_signal_reg[45]  (.D(n_0_236), .G(n_0_188), .Q(out_c[45]));
   DLH_X1 \out_c_signal_reg[44]  (.D(n_0_235), .G(n_0_188), .Q(out_c[44]));
   DLH_X1 \out_c_signal_reg[43]  (.D(n_0_234), .G(n_0_188), .Q(out_c[43]));
   DLH_X1 \out_c_signal_reg[42]  (.D(n_0_233), .G(n_0_188), .Q(out_c[42]));
   DLH_X1 \out_c_signal_reg[41]  (.D(n_0_232), .G(n_0_188), .Q(out_c[41]));
   DLH_X1 \out_c_signal_reg[40]  (.D(n_0_231), .G(n_0_188), .Q(out_c[40]));
   DLH_X1 \out_c_signal_reg[39]  (.D(n_0_230), .G(n_0_188), .Q(out_c[39]));
   DLH_X1 \out_c_signal_reg[38]  (.D(n_0_229), .G(n_0_188), .Q(out_c[38]));
   DLH_X1 \out_c_signal_reg[37]  (.D(n_0_228), .G(n_0_188), .Q(out_c[37]));
   DLH_X1 \out_c_signal_reg[36]  (.D(n_0_227), .G(n_0_188), .Q(out_c[36]));
   DLH_X1 \out_c_signal_reg[35]  (.D(n_0_226), .G(n_0_188), .Q(out_c[35]));
   DLH_X1 \out_c_signal_reg[34]  (.D(n_0_225), .G(n_0_188), .Q(out_c[34]));
   DLH_X1 \out_c_signal_reg[33]  (.D(n_0_224), .G(n_0_188), .Q(out_c[33]));
   DLH_X1 \out_c_signal_reg[32]  (.D(n_0_223), .G(n_0_188), .Q(out_c[32]));
   DLH_X1 \out_c_signal_reg[31]  (.D(n_0_222), .G(n_0_188), .Q(out_c[31]));
   DLH_X1 \out_c_signal_reg[30]  (.D(n_0_221), .G(n_0_188), .Q(out_c[30]));
   DLH_X1 \out_c_signal_reg[29]  (.D(n_0_220), .G(n_0_188), .Q(out_c[29]));
   DLH_X1 \out_c_signal_reg[28]  (.D(n_0_219), .G(n_0_188), .Q(out_c[28]));
   DLH_X1 \out_c_signal_reg[27]  (.D(n_0_218), .G(n_0_188), .Q(out_c[27]));
   DLH_X1 \out_c_signal_reg[26]  (.D(n_0_217), .G(n_0_188), .Q(out_c[26]));
   DLH_X1 \out_c_signal_reg[25]  (.D(n_0_216), .G(n_0_188), .Q(out_c[25]));
   DLH_X1 \out_c_signal_reg[24]  (.D(n_0_215), .G(n_0_188), .Q(out_c[24]));
   DLH_X1 \out_c_signal_reg[23]  (.D(n_0_214), .G(n_0_188), .Q(out_c[23]));
   DLH_X1 \out_c_signal_reg[22]  (.D(n_0_213), .G(n_0_188), .Q(out_c[22]));
   DLH_X1 \out_c_signal_reg[21]  (.D(n_0_212), .G(n_0_188), .Q(out_c[21]));
   DLH_X1 \out_c_signal_reg[20]  (.D(n_0_211), .G(n_0_188), .Q(out_c[20]));
   DLH_X1 \out_c_signal_reg[19]  (.D(n_0_210), .G(n_0_188), .Q(out_c[19]));
   DLH_X1 \out_c_signal_reg[18]  (.D(n_0_209), .G(n_0_188), .Q(out_c[18]));
   DLH_X1 \out_c_signal_reg[17]  (.D(n_0_208), .G(n_0_188), .Q(out_c[17]));
   DLH_X1 \out_c_signal_reg[16]  (.D(n_0_207), .G(n_0_188), .Q(out_c[16]));
   DLH_X1 \out_c_signal_reg[15]  (.D(n_0_206), .G(n_0_188), .Q(out_c[15]));
   DLH_X1 \out_c_signal_reg[14]  (.D(n_0_205), .G(n_0_188), .Q(out_c[14]));
   DLH_X1 \out_c_signal_reg[13]  (.D(n_0_204), .G(n_0_188), .Q(out_c[13]));
   DLH_X1 \out_c_signal_reg[12]  (.D(n_0_203), .G(n_0_188), .Q(out_c[12]));
   DLH_X1 \out_c_signal_reg[11]  (.D(n_0_202), .G(n_0_188), .Q(out_c[11]));
   DLH_X1 \out_c_signal_reg[10]  (.D(n_0_201), .G(n_0_188), .Q(out_c[10]));
   DLH_X1 \out_c_signal_reg[9]  (.D(n_0_200), .G(n_0_188), .Q(out_c[9]));
   DLH_X1 \out_c_signal_reg[8]  (.D(n_0_199), .G(n_0_188), .Q(out_c[8]));
   DLH_X1 \out_c_signal_reg[7]  (.D(n_0_198), .G(n_0_188), .Q(out_c[7]));
   DLH_X1 \out_c_signal_reg[6]  (.D(n_0_197), .G(n_0_188), .Q(out_c[6]));
   DLH_X1 \out_c_signal_reg[5]  (.D(n_0_196), .G(n_0_188), .Q(out_c[5]));
   DLH_X1 \out_c_signal_reg[4]  (.D(n_0_195), .G(n_0_188), .Q(out_c[4]));
   DLH_X1 \out_c_signal_reg[3]  (.D(n_0_194), .G(n_0_188), .Q(out_c[3]));
   DLH_X1 \out_c_signal_reg[2]  (.D(n_0_193), .G(n_0_188), .Q(out_c[2]));
   DLH_X1 \out_c_signal_reg[1]  (.D(n_0_192), .G(n_0_188), .Q(out_c[1]));
   DLH_X1 \out_c_signal_reg[0]  (.D(FA1_n_0), .G(n_0_188), .Q(out_c[0]));
   DLH_X1 \in_b_signal_reg[63]  (.D(n_0_187), .G(n_0_188), .Q(in_b_signal));
   DLH_X1 \in_b_signal_reg[62]  (.D(n_0_186), .G(n_0_188), .Q(n_0_0));
   DLH_X1 \in_b_signal_reg[61]  (.D(n_0_185), .G(n_0_188), .Q(n_0_1));
   DLH_X1 \in_b_signal_reg[60]  (.D(n_0_184), .G(n_0_188), .Q(n_0_2));
   DLH_X1 \in_b_signal_reg[59]  (.D(n_0_183), .G(n_0_188), .Q(n_0_3));
   DLH_X1 \in_b_signal_reg[58]  (.D(n_0_182), .G(n_0_188), .Q(n_0_4));
   DLH_X1 \in_b_signal_reg[57]  (.D(n_0_181), .G(n_0_188), .Q(n_0_5));
   DLH_X1 \in_b_signal_reg[56]  (.D(n_0_180), .G(n_0_188), .Q(n_0_6));
   DLH_X1 \in_b_signal_reg[55]  (.D(n_0_179), .G(n_0_188), .Q(n_0_7));
   DLH_X1 \in_b_signal_reg[54]  (.D(n_0_178), .G(n_0_188), .Q(n_0_8));
   DLH_X1 \in_b_signal_reg[53]  (.D(n_0_177), .G(n_0_188), .Q(n_0_9));
   DLH_X1 \in_b_signal_reg[52]  (.D(n_0_176), .G(n_0_188), .Q(n_0_10));
   DLH_X1 \in_b_signal_reg[51]  (.D(n_0_175), .G(n_0_188), .Q(n_0_11));
   DLH_X1 \in_b_signal_reg[50]  (.D(n_0_174), .G(n_0_188), .Q(n_0_12));
   DLH_X1 \in_b_signal_reg[49]  (.D(n_0_173), .G(n_0_188), .Q(n_0_13));
   DLH_X1 \in_b_signal_reg[48]  (.D(n_0_172), .G(n_0_188), .Q(n_0_14));
   DLH_X1 \in_b_signal_reg[47]  (.D(n_0_171), .G(n_0_188), .Q(n_0_15));
   DLH_X1 \in_b_signal_reg[46]  (.D(n_0_170), .G(n_0_188), .Q(n_0_16));
   DLH_X1 \in_b_signal_reg[45]  (.D(n_0_169), .G(n_0_188), .Q(n_0_17));
   DLH_X1 \in_b_signal_reg[44]  (.D(n_0_168), .G(n_0_188), .Q(n_0_18));
   DLH_X1 \in_b_signal_reg[43]  (.D(n_0_167), .G(n_0_188), .Q(n_0_19));
   DLH_X1 \in_b_signal_reg[42]  (.D(n_0_166), .G(n_0_188), .Q(n_0_20));
   DLH_X1 \in_b_signal_reg[41]  (.D(n_0_165), .G(n_0_188), .Q(n_0_21));
   DLH_X1 \in_b_signal_reg[40]  (.D(n_0_164), .G(n_0_188), .Q(n_0_22));
   DLH_X1 \in_b_signal_reg[39]  (.D(n_0_163), .G(n_0_188), .Q(n_0_23));
   DLH_X1 \in_b_signal_reg[38]  (.D(n_0_162), .G(n_0_188), .Q(n_0_24));
   DLH_X1 \in_b_signal_reg[37]  (.D(n_0_161), .G(n_0_188), .Q(n_0_25));
   DLH_X1 \in_b_signal_reg[36]  (.D(n_0_160), .G(n_0_188), .Q(n_0_26));
   DLH_X1 \in_b_signal_reg[35]  (.D(n_0_159), .G(n_0_188), .Q(n_0_27));
   DLH_X1 \in_b_signal_reg[34]  (.D(n_0_158), .G(n_0_188), .Q(n_0_28));
   DLH_X1 \in_b_signal_reg[33]  (.D(n_0_157), .G(n_0_188), .Q(n_0_29));
   DLH_X1 \in_b_signal_reg[32]  (.D(n_0_156), .G(n_0_188), .Q(n_0_30));
   DLH_X1 \in_b_signal_reg[31]  (.D(n_0_155), .G(n_0_188), .Q(n_0_31));
   DLH_X1 \in_b_signal_reg[30]  (.D(n_0_154), .G(n_0_188), .Q(n_0_32));
   DLH_X1 \in_b_signal_reg[29]  (.D(n_0_153), .G(n_0_188), .Q(n_0_33));
   DLH_X1 \in_b_signal_reg[28]  (.D(n_0_152), .G(n_0_188), .Q(n_0_34));
   DLH_X1 \in_b_signal_reg[27]  (.D(n_0_151), .G(n_0_188), .Q(n_0_35));
   DLH_X1 \in_b_signal_reg[26]  (.D(n_0_150), .G(n_0_188), .Q(n_0_36));
   DLH_X1 \in_b_signal_reg[25]  (.D(n_0_149), .G(n_0_188), .Q(n_0_37));
   DLH_X1 \in_b_signal_reg[24]  (.D(n_0_148), .G(n_0_188), .Q(n_0_38));
   DLH_X1 \in_b_signal_reg[23]  (.D(n_0_147), .G(n_0_188), .Q(n_0_39));
   DLH_X1 \in_b_signal_reg[22]  (.D(n_0_146), .G(n_0_188), .Q(n_0_40));
   DLH_X1 \in_b_signal_reg[21]  (.D(n_0_145), .G(n_0_188), .Q(n_0_41));
   DLH_X1 \in_b_signal_reg[20]  (.D(n_0_144), .G(n_0_188), .Q(n_0_42));
   DLH_X1 \in_b_signal_reg[19]  (.D(n_0_143), .G(n_0_188), .Q(n_0_43));
   DLH_X1 \in_b_signal_reg[18]  (.D(n_0_142), .G(n_0_188), .Q(n_0_44));
   DLH_X1 \in_b_signal_reg[17]  (.D(n_0_141), .G(n_0_188), .Q(n_0_45));
   DLH_X1 \in_b_signal_reg[16]  (.D(n_0_140), .G(n_0_188), .Q(n_0_46));
   DLH_X1 \in_b_signal_reg[15]  (.D(n_0_139), .G(n_0_188), .Q(n_0_47));
   DLH_X1 \in_b_signal_reg[14]  (.D(n_0_138), .G(n_0_188), .Q(n_0_48));
   DLH_X1 \in_b_signal_reg[13]  (.D(n_0_137), .G(n_0_188), .Q(n_0_49));
   DLH_X1 \in_b_signal_reg[12]  (.D(n_0_136), .G(n_0_188), .Q(n_0_50));
   DLH_X1 \in_b_signal_reg[11]  (.D(n_0_135), .G(n_0_188), .Q(n_0_51));
   DLH_X1 \in_b_signal_reg[10]  (.D(n_0_134), .G(n_0_188), .Q(n_0_52));
   DLH_X1 \in_b_signal_reg[9]  (.D(n_0_133), .G(n_0_188), .Q(n_0_53));
   DLH_X1 \in_b_signal_reg[8]  (.D(n_0_132), .G(n_0_188), .Q(n_0_54));
   DLH_X1 \in_b_signal_reg[7]  (.D(n_0_131), .G(n_0_188), .Q(n_0_55));
   DLH_X1 \in_b_signal_reg[6]  (.D(n_0_130), .G(n_0_188), .Q(n_0_56));
   DLH_X1 \in_b_signal_reg[5]  (.D(n_0_129), .G(n_0_188), .Q(n_0_57));
   DLH_X1 \in_b_signal_reg[4]  (.D(n_0_128), .G(n_0_188), .Q(n_0_58));
   DLH_X1 \in_b_signal_reg[3]  (.D(n_0_127), .G(n_0_188), .Q(n_0_59));
   DLH_X1 \in_b_signal_reg[2]  (.D(n_0_126), .G(n_0_188), .Q(n_0_60));
   DLH_X1 \in_b_signal_reg[1]  (.D(n_0_125), .G(n_0_188), .Q(b));
   DLH_X1 \in_b_signal_reg[0]  (.D(in_b[0]), .G(n_0_188), .Q(n_0_61));
   datapath i_0_9 (.plus({n_0_124, n_0_123, n_0_122, n_0_121, n_0_120, n_0_119, 
      n_0_118, n_0_117, n_0_116, n_0_115, n_0_114, n_0_113, n_0_112, n_0_111, 
      n_0_110, n_0_109, n_0_108, n_0_107, n_0_106, n_0_105, n_0_104, n_0_103, 
      n_0_102, n_0_101, n_0_100, n_0_99, n_0_98, n_0_97, n_0_96, n_0_95, n_0_94, 
      n_0_93, n_0_92, n_0_91, n_0_90, n_0_89, n_0_88, n_0_87, n_0_86, n_0_85, 
      n_0_84, n_0_83, n_0_82, n_0_81, n_0_80, n_0_79, n_0_78, n_0_77, n_0_76, 
      n_0_75, n_0_74, n_0_73, n_0_72, n_0_71, n_0_70, n_0_69, n_0_68, n_0_67, 
      n_0_66, n_0_65, n_0_64, n_0_63, n_0_62, uc_0}), .in_b(in_b));
   NAND2_X1 i_0_0_0 (.A1(n_0_0_0), .A2(n_0_0_1), .ZN(done));
   INV_X1 i_0_0_1 (.A(enbl), .ZN(n_0_0_0));
   INV_X1 i_0_0_2 (.A(rst), .ZN(n_0_0_1));
   NAND2_X1 i_0_1_0 (.A1(add_sub), .A2(enbl), .ZN(n_0_1_0));
   INV_X1 i_0_1_1 (.A(n_0_1_0), .ZN(n_0_1_1));
   OAI22_X1 i_0_1_2 (.A1(n_0_1_1), .A2(in_b[1]), .B1(n_0_1_0), .B2(n_0_62), 
      .ZN(n_0_1_2));
   INV_X1 i_0_1_3 (.A(n_0_1_2), .ZN(n_0_125));
   OAI22_X1 i_0_1_4 (.A1(n_0_1_1), .A2(in_b[2]), .B1(n_0_1_0), .B2(n_0_63), 
      .ZN(n_0_1_3));
   INV_X1 i_0_1_5 (.A(n_0_1_3), .ZN(n_0_126));
   OAI22_X1 i_0_1_6 (.A1(n_0_1_1), .A2(in_b[3]), .B1(n_0_1_0), .B2(n_0_64), 
      .ZN(n_0_1_4));
   INV_X1 i_0_1_7 (.A(n_0_1_4), .ZN(n_0_127));
   OAI22_X1 i_0_1_8 (.A1(n_0_1_1), .A2(in_b[4]), .B1(n_0_1_0), .B2(n_0_65), 
      .ZN(n_0_1_5));
   INV_X1 i_0_1_9 (.A(n_0_1_5), .ZN(n_0_128));
   OAI22_X1 i_0_1_10 (.A1(n_0_1_1), .A2(in_b[5]), .B1(n_0_1_0), .B2(n_0_66), 
      .ZN(n_0_1_6));
   INV_X1 i_0_1_11 (.A(n_0_1_6), .ZN(n_0_129));
   OAI22_X1 i_0_1_12 (.A1(n_0_1_1), .A2(in_b[6]), .B1(n_0_1_0), .B2(n_0_67), 
      .ZN(n_0_1_7));
   INV_X1 i_0_1_13 (.A(n_0_1_7), .ZN(n_0_130));
   OAI22_X1 i_0_1_14 (.A1(n_0_1_1), .A2(in_b[7]), .B1(n_0_1_0), .B2(n_0_68), 
      .ZN(n_0_1_8));
   INV_X1 i_0_1_15 (.A(n_0_1_8), .ZN(n_0_131));
   OAI22_X1 i_0_1_16 (.A1(n_0_1_1), .A2(in_b[8]), .B1(n_0_1_0), .B2(n_0_69), 
      .ZN(n_0_1_9));
   INV_X1 i_0_1_17 (.A(n_0_1_9), .ZN(n_0_132));
   OAI22_X1 i_0_1_18 (.A1(n_0_1_1), .A2(in_b[9]), .B1(n_0_1_0), .B2(n_0_70), 
      .ZN(n_0_1_10));
   INV_X1 i_0_1_19 (.A(n_0_1_10), .ZN(n_0_133));
   OAI22_X1 i_0_1_20 (.A1(n_0_1_1), .A2(in_b[10]), .B1(n_0_1_0), .B2(n_0_71), 
      .ZN(n_0_1_11));
   INV_X1 i_0_1_21 (.A(n_0_1_11), .ZN(n_0_134));
   OAI22_X1 i_0_1_22 (.A1(n_0_1_1), .A2(in_b[11]), .B1(n_0_1_0), .B2(n_0_72), 
      .ZN(n_0_1_12));
   INV_X1 i_0_1_23 (.A(n_0_1_12), .ZN(n_0_135));
   OAI22_X1 i_0_1_24 (.A1(n_0_1_1), .A2(in_b[12]), .B1(n_0_1_0), .B2(n_0_73), 
      .ZN(n_0_1_13));
   INV_X1 i_0_1_25 (.A(n_0_1_13), .ZN(n_0_136));
   OAI22_X1 i_0_1_26 (.A1(n_0_1_1), .A2(in_b[13]), .B1(n_0_1_0), .B2(n_0_74), 
      .ZN(n_0_1_14));
   INV_X1 i_0_1_27 (.A(n_0_1_14), .ZN(n_0_137));
   OAI22_X1 i_0_1_28 (.A1(n_0_1_1), .A2(in_b[14]), .B1(n_0_1_0), .B2(n_0_75), 
      .ZN(n_0_1_15));
   INV_X1 i_0_1_29 (.A(n_0_1_15), .ZN(n_0_138));
   OAI22_X1 i_0_1_30 (.A1(n_0_1_1), .A2(in_b[15]), .B1(n_0_1_0), .B2(n_0_76), 
      .ZN(n_0_1_16));
   INV_X1 i_0_1_31 (.A(n_0_1_16), .ZN(n_0_139));
   OAI22_X1 i_0_1_32 (.A1(n_0_1_1), .A2(in_b[16]), .B1(n_0_1_0), .B2(n_0_77), 
      .ZN(n_0_1_17));
   INV_X1 i_0_1_33 (.A(n_0_1_17), .ZN(n_0_140));
   OAI22_X1 i_0_1_34 (.A1(n_0_1_1), .A2(in_b[17]), .B1(n_0_1_0), .B2(n_0_78), 
      .ZN(n_0_1_18));
   INV_X1 i_0_1_35 (.A(n_0_1_18), .ZN(n_0_141));
   OAI22_X1 i_0_1_36 (.A1(n_0_1_1), .A2(in_b[18]), .B1(n_0_1_0), .B2(n_0_79), 
      .ZN(n_0_1_19));
   INV_X1 i_0_1_37 (.A(n_0_1_19), .ZN(n_0_142));
   OAI22_X1 i_0_1_38 (.A1(n_0_1_1), .A2(in_b[19]), .B1(n_0_1_0), .B2(n_0_80), 
      .ZN(n_0_1_20));
   INV_X1 i_0_1_39 (.A(n_0_1_20), .ZN(n_0_143));
   OAI22_X1 i_0_1_40 (.A1(n_0_1_1), .A2(in_b[20]), .B1(n_0_1_0), .B2(n_0_81), 
      .ZN(n_0_1_21));
   INV_X1 i_0_1_41 (.A(n_0_1_21), .ZN(n_0_144));
   OAI22_X1 i_0_1_42 (.A1(n_0_1_1), .A2(in_b[21]), .B1(n_0_1_0), .B2(n_0_82), 
      .ZN(n_0_1_22));
   INV_X1 i_0_1_43 (.A(n_0_1_22), .ZN(n_0_145));
   OAI22_X1 i_0_1_44 (.A1(n_0_1_1), .A2(in_b[22]), .B1(n_0_1_0), .B2(n_0_83), 
      .ZN(n_0_1_23));
   INV_X1 i_0_1_45 (.A(n_0_1_23), .ZN(n_0_146));
   OAI22_X1 i_0_1_46 (.A1(n_0_1_1), .A2(in_b[23]), .B1(n_0_1_0), .B2(n_0_84), 
      .ZN(n_0_1_24));
   INV_X1 i_0_1_47 (.A(n_0_1_24), .ZN(n_0_147));
   OAI22_X1 i_0_1_48 (.A1(n_0_1_1), .A2(in_b[24]), .B1(n_0_1_0), .B2(n_0_85), 
      .ZN(n_0_1_25));
   INV_X1 i_0_1_49 (.A(n_0_1_25), .ZN(n_0_148));
   OAI22_X1 i_0_1_50 (.A1(n_0_1_1), .A2(in_b[25]), .B1(n_0_1_0), .B2(n_0_86), 
      .ZN(n_0_1_26));
   INV_X1 i_0_1_51 (.A(n_0_1_26), .ZN(n_0_149));
   OAI22_X1 i_0_1_52 (.A1(n_0_1_1), .A2(in_b[26]), .B1(n_0_1_0), .B2(n_0_87), 
      .ZN(n_0_1_27));
   INV_X1 i_0_1_53 (.A(n_0_1_27), .ZN(n_0_150));
   OAI22_X1 i_0_1_54 (.A1(n_0_1_1), .A2(in_b[27]), .B1(n_0_1_0), .B2(n_0_88), 
      .ZN(n_0_1_28));
   INV_X1 i_0_1_55 (.A(n_0_1_28), .ZN(n_0_151));
   OAI22_X1 i_0_1_56 (.A1(n_0_1_1), .A2(in_b[28]), .B1(n_0_1_0), .B2(n_0_89), 
      .ZN(n_0_1_29));
   INV_X1 i_0_1_57 (.A(n_0_1_29), .ZN(n_0_152));
   OAI22_X1 i_0_1_58 (.A1(n_0_1_1), .A2(in_b[29]), .B1(n_0_1_0), .B2(n_0_90), 
      .ZN(n_0_1_30));
   INV_X1 i_0_1_59 (.A(n_0_1_30), .ZN(n_0_153));
   OAI22_X1 i_0_1_60 (.A1(n_0_1_1), .A2(in_b[30]), .B1(n_0_1_0), .B2(n_0_91), 
      .ZN(n_0_1_31));
   INV_X1 i_0_1_61 (.A(n_0_1_31), .ZN(n_0_154));
   OAI22_X1 i_0_1_62 (.A1(n_0_1_1), .A2(in_b[31]), .B1(n_0_1_0), .B2(n_0_92), 
      .ZN(n_0_1_32));
   INV_X1 i_0_1_63 (.A(n_0_1_32), .ZN(n_0_155));
   OAI22_X1 i_0_1_64 (.A1(n_0_1_1), .A2(in_b[32]), .B1(n_0_1_0), .B2(n_0_93), 
      .ZN(n_0_1_33));
   INV_X1 i_0_1_65 (.A(n_0_1_33), .ZN(n_0_156));
   OAI22_X1 i_0_1_66 (.A1(n_0_1_1), .A2(in_b[33]), .B1(n_0_1_0), .B2(n_0_94), 
      .ZN(n_0_1_34));
   INV_X1 i_0_1_67 (.A(n_0_1_34), .ZN(n_0_157));
   OAI22_X1 i_0_1_68 (.A1(n_0_1_1), .A2(in_b[34]), .B1(n_0_1_0), .B2(n_0_95), 
      .ZN(n_0_1_35));
   INV_X1 i_0_1_69 (.A(n_0_1_35), .ZN(n_0_158));
   OAI22_X1 i_0_1_70 (.A1(n_0_1_1), .A2(in_b[35]), .B1(n_0_1_0), .B2(n_0_96), 
      .ZN(n_0_1_36));
   INV_X1 i_0_1_71 (.A(n_0_1_36), .ZN(n_0_159));
   OAI22_X1 i_0_1_72 (.A1(n_0_1_1), .A2(in_b[36]), .B1(n_0_1_0), .B2(n_0_97), 
      .ZN(n_0_1_37));
   INV_X1 i_0_1_73 (.A(n_0_1_37), .ZN(n_0_160));
   OAI22_X1 i_0_1_74 (.A1(n_0_1_1), .A2(in_b[37]), .B1(n_0_1_0), .B2(n_0_98), 
      .ZN(n_0_1_38));
   INV_X1 i_0_1_75 (.A(n_0_1_38), .ZN(n_0_161));
   OAI22_X1 i_0_1_76 (.A1(n_0_1_1), .A2(in_b[38]), .B1(n_0_1_0), .B2(n_0_99), 
      .ZN(n_0_1_39));
   INV_X1 i_0_1_77 (.A(n_0_1_39), .ZN(n_0_162));
   OAI22_X1 i_0_1_78 (.A1(n_0_1_1), .A2(in_b[39]), .B1(n_0_1_0), .B2(n_0_100), 
      .ZN(n_0_1_40));
   INV_X1 i_0_1_79 (.A(n_0_1_40), .ZN(n_0_163));
   OAI22_X1 i_0_1_80 (.A1(n_0_1_1), .A2(in_b[40]), .B1(n_0_1_0), .B2(n_0_101), 
      .ZN(n_0_1_41));
   INV_X1 i_0_1_81 (.A(n_0_1_41), .ZN(n_0_164));
   OAI22_X1 i_0_1_82 (.A1(n_0_1_1), .A2(in_b[41]), .B1(n_0_1_0), .B2(n_0_102), 
      .ZN(n_0_1_42));
   INV_X1 i_0_1_83 (.A(n_0_1_42), .ZN(n_0_165));
   OAI22_X1 i_0_1_84 (.A1(n_0_1_1), .A2(in_b[42]), .B1(n_0_1_0), .B2(n_0_103), 
      .ZN(n_0_1_43));
   INV_X1 i_0_1_85 (.A(n_0_1_43), .ZN(n_0_166));
   OAI22_X1 i_0_1_86 (.A1(n_0_1_1), .A2(in_b[43]), .B1(n_0_1_0), .B2(n_0_104), 
      .ZN(n_0_1_44));
   INV_X1 i_0_1_87 (.A(n_0_1_44), .ZN(n_0_167));
   OAI22_X1 i_0_1_88 (.A1(n_0_1_1), .A2(in_b[44]), .B1(n_0_1_0), .B2(n_0_105), 
      .ZN(n_0_1_45));
   INV_X1 i_0_1_89 (.A(n_0_1_45), .ZN(n_0_168));
   OAI22_X1 i_0_1_90 (.A1(n_0_1_1), .A2(in_b[45]), .B1(n_0_1_0), .B2(n_0_106), 
      .ZN(n_0_1_46));
   INV_X1 i_0_1_91 (.A(n_0_1_46), .ZN(n_0_169));
   OAI22_X1 i_0_1_92 (.A1(n_0_1_1), .A2(in_b[46]), .B1(n_0_1_0), .B2(n_0_107), 
      .ZN(n_0_1_47));
   INV_X1 i_0_1_93 (.A(n_0_1_47), .ZN(n_0_170));
   OAI22_X1 i_0_1_94 (.A1(n_0_1_1), .A2(in_b[47]), .B1(n_0_1_0), .B2(n_0_108), 
      .ZN(n_0_1_48));
   INV_X1 i_0_1_95 (.A(n_0_1_48), .ZN(n_0_171));
   OAI22_X1 i_0_1_96 (.A1(n_0_1_1), .A2(in_b[48]), .B1(n_0_1_0), .B2(n_0_109), 
      .ZN(n_0_1_49));
   INV_X1 i_0_1_97 (.A(n_0_1_49), .ZN(n_0_172));
   OAI22_X1 i_0_1_98 (.A1(n_0_1_1), .A2(in_b[49]), .B1(n_0_1_0), .B2(n_0_110), 
      .ZN(n_0_1_50));
   INV_X1 i_0_1_99 (.A(n_0_1_50), .ZN(n_0_173));
   OAI22_X1 i_0_1_100 (.A1(n_0_1_1), .A2(in_b[50]), .B1(n_0_1_0), .B2(n_0_111), 
      .ZN(n_0_1_51));
   INV_X1 i_0_1_101 (.A(n_0_1_51), .ZN(n_0_174));
   OAI22_X1 i_0_1_102 (.A1(n_0_1_1), .A2(in_b[51]), .B1(n_0_1_0), .B2(n_0_112), 
      .ZN(n_0_1_52));
   INV_X1 i_0_1_103 (.A(n_0_1_52), .ZN(n_0_175));
   OAI22_X1 i_0_1_104 (.A1(n_0_1_1), .A2(in_b[52]), .B1(n_0_1_0), .B2(n_0_113), 
      .ZN(n_0_1_53));
   INV_X1 i_0_1_105 (.A(n_0_1_53), .ZN(n_0_176));
   OAI22_X1 i_0_1_106 (.A1(n_0_1_1), .A2(in_b[53]), .B1(n_0_1_0), .B2(n_0_114), 
      .ZN(n_0_1_54));
   INV_X1 i_0_1_107 (.A(n_0_1_54), .ZN(n_0_177));
   OAI22_X1 i_0_1_108 (.A1(n_0_1_1), .A2(in_b[54]), .B1(n_0_1_0), .B2(n_0_115), 
      .ZN(n_0_1_55));
   INV_X1 i_0_1_109 (.A(n_0_1_55), .ZN(n_0_178));
   OAI22_X1 i_0_1_110 (.A1(n_0_1_1), .A2(in_b[55]), .B1(n_0_1_0), .B2(n_0_116), 
      .ZN(n_0_1_56));
   INV_X1 i_0_1_111 (.A(n_0_1_56), .ZN(n_0_179));
   OAI22_X1 i_0_1_112 (.A1(n_0_1_1), .A2(in_b[56]), .B1(n_0_1_0), .B2(n_0_117), 
      .ZN(n_0_1_57));
   INV_X1 i_0_1_113 (.A(n_0_1_57), .ZN(n_0_180));
   OAI22_X1 i_0_1_114 (.A1(n_0_1_1), .A2(in_b[57]), .B1(n_0_1_0), .B2(n_0_118), 
      .ZN(n_0_1_58));
   INV_X1 i_0_1_115 (.A(n_0_1_58), .ZN(n_0_181));
   OAI22_X1 i_0_1_116 (.A1(n_0_1_1), .A2(in_b[58]), .B1(n_0_1_0), .B2(n_0_119), 
      .ZN(n_0_1_59));
   INV_X1 i_0_1_117 (.A(n_0_1_59), .ZN(n_0_182));
   OAI22_X1 i_0_1_118 (.A1(n_0_1_1), .A2(in_b[59]), .B1(n_0_1_0), .B2(n_0_120), 
      .ZN(n_0_1_60));
   INV_X1 i_0_1_119 (.A(n_0_1_60), .ZN(n_0_183));
   OAI22_X1 i_0_1_120 (.A1(n_0_1_1), .A2(in_b[60]), .B1(n_0_1_0), .B2(n_0_121), 
      .ZN(n_0_1_61));
   INV_X1 i_0_1_121 (.A(n_0_1_61), .ZN(n_0_184));
   OAI22_X1 i_0_1_122 (.A1(n_0_1_1), .A2(in_b[61]), .B1(n_0_1_0), .B2(n_0_122), 
      .ZN(n_0_1_62));
   INV_X1 i_0_1_123 (.A(n_0_1_62), .ZN(n_0_185));
   OAI22_X1 i_0_1_124 (.A1(n_0_1_1), .A2(in_b[62]), .B1(n_0_1_0), .B2(n_0_123), 
      .ZN(n_0_1_63));
   INV_X1 i_0_1_125 (.A(n_0_1_63), .ZN(n_0_186));
   OAI22_X1 i_0_1_126 (.A1(n_0_1_1), .A2(in_b[63]), .B1(n_0_1_0), .B2(n_0_124), 
      .ZN(n_0_1_64));
   INV_X1 i_0_1_127 (.A(n_0_1_64), .ZN(n_0_187));
   INV_X1 i_0_1_128 (.A(rst), .ZN(n_0_1_65));
   AND2_X1 i_0_1_129 (.A1(n_0_1_65), .A2(enbl), .ZN(n_0_188));
   OAI21_X1 i_0_1_130 (.A(n_0_1_65), .B1(in_b_signal), .B2(out_c[63]), .ZN(
      n_0_1_66));
   XOR2_X1 i_0_1_131 (.A(in_a[63]), .B(in_b_signal), .Z(n_0_1_67));
   AOI211_X1 i_0_1_132 (.A(n_0_1_66), .B(n_0_1_67), .C1(in_b_signal), .C2(
      out_c[63]), .ZN(n_0_189));
   NOR4_X1 i_0_1_133 (.A1(out_c[42]), .A2(out_c[41]), .A3(out_c[47]), .A4(
      out_c[44]), .ZN(n_0_1_68));
   NOR4_X1 i_0_1_134 (.A1(out_c[35]), .A2(out_c[32]), .A3(out_c[38]), .A4(
      out_c[37]), .ZN(n_0_1_69));
   NOR4_X1 i_0_1_135 (.A1(out_c[59]), .A2(out_c[56]), .A3(out_c[62]), .A4(
      out_c[61]), .ZN(n_0_1_70));
   NOR4_X1 i_0_1_136 (.A1(out_c[50]), .A2(out_c[49]), .A3(out_c[55]), .A4(
      out_c[52]), .ZN(n_0_1_71));
   NAND4_X1 i_0_1_137 (.A1(n_0_1_68), .A2(n_0_1_69), .A3(n_0_1_70), .A4(n_0_1_71), 
      .ZN(n_0_1_72));
   NOR4_X1 i_0_1_138 (.A1(out_c[11]), .A2(out_c[8]), .A3(out_c[14]), .A4(
      out_c[13]), .ZN(n_0_1_73));
   NOR4_X1 i_0_1_139 (.A1(out_c[2]), .A2(out_c[1]), .A3(out_c[7]), .A4(out_c[4]), 
      .ZN(n_0_1_74));
   NOR4_X1 i_0_1_140 (.A1(out_c[26]), .A2(out_c[25]), .A3(out_c[31]), .A4(
      out_c[28]), .ZN(n_0_1_75));
   NOR4_X1 i_0_1_141 (.A1(out_c[19]), .A2(out_c[16]), .A3(out_c[22]), .A4(
      out_c[21]), .ZN(n_0_1_76));
   NAND4_X1 i_0_1_142 (.A1(n_0_1_73), .A2(n_0_1_74), .A3(n_0_1_75), .A4(n_0_1_76), 
      .ZN(n_0_1_77));
   NOR4_X1 i_0_1_143 (.A1(out_c[10]), .A2(out_c[9]), .A3(out_c[15]), .A4(
      out_c[12]), .ZN(n_0_1_78));
   NOR4_X1 i_0_1_144 (.A1(out_c[3]), .A2(out_c[0]), .A3(out_c[6]), .A4(out_c[5]), 
      .ZN(n_0_1_79));
   NOR4_X1 i_0_1_145 (.A1(out_c[27]), .A2(out_c[24]), .A3(out_c[30]), .A4(
      out_c[29]), .ZN(n_0_1_80));
   NOR4_X1 i_0_1_146 (.A1(out_c[18]), .A2(out_c[17]), .A3(out_c[23]), .A4(
      out_c[20]), .ZN(n_0_1_81));
   NAND4_X1 i_0_1_147 (.A1(n_0_1_78), .A2(n_0_1_79), .A3(n_0_1_80), .A4(n_0_1_81), 
      .ZN(n_0_1_82));
   OR3_X1 i_0_1_148 (.A1(n_0_1_72), .A2(n_0_1_77), .A3(n_0_1_82), .ZN(n_0_1_83));
   NOR4_X1 i_0_1_149 (.A1(out_c[43]), .A2(out_c[40]), .A3(out_c[46]), .A4(
      out_c[45]), .ZN(n_0_1_84));
   NOR4_X1 i_0_1_150 (.A1(out_c[34]), .A2(out_c[33]), .A3(out_c[39]), .A4(
      out_c[36]), .ZN(n_0_1_85));
   NOR4_X1 i_0_1_151 (.A1(out_c[58]), .A2(out_c[57]), .A3(out_c[60]), .A4(
      out_c[63]), .ZN(n_0_1_86));
   NOR4_X1 i_0_1_152 (.A1(out_c[51]), .A2(out_c[48]), .A3(out_c[54]), .A4(
      out_c[53]), .ZN(n_0_1_87));
   NAND4_X1 i_0_1_153 (.A1(n_0_1_84), .A2(n_0_1_85), .A3(n_0_1_86), .A4(n_0_1_87), 
      .ZN(n_0_1_88));
   OAI21_X1 i_0_1_154 (.A(n_0_1_65), .B1(n_0_1_83), .B2(n_0_1_88), .ZN(n_0_190));
   NOR3_X1 i_0_1_155 (.A1(zero), .A2(rst), .A3(out_c[63]), .ZN(n_0_191));
   NAND2_X1 i_0_1_156 (.A1(n_0_61), .A2(in_a[0]), .ZN(n_0_1_89));
   INV_X1 i_0_1_157 (.A(n_0_1_89), .ZN(n_0_1_90));
   INV_X1 i_0_1_158 (.A(n_0_61), .ZN(n_0_1_91));
   INV_X1 i_0_1_159 (.A(in_a[0]), .ZN(n_0_1_92));
   AOI21_X1 i_0_1_160 (.A(n_0_1_90), .B1(n_0_1_91), .B2(n_0_1_92), .ZN(FA1_n_0));
   NAND2_X1 i_0_1_161 (.A1(b), .A2(in_a[1]), .ZN(n_0_1_93));
   OAI21_X1 i_0_1_162 (.A(n_0_1_93), .B1(b), .B2(in_a[1]), .ZN(n_0_1_94));
   XOR2_X1 i_0_1_163 (.A(n_0_1_94), .B(n_0_1_89), .Z(n_0_192));
   OAI21_X1 i_0_1_164 (.A(n_0_1_93), .B1(n_0_1_94), .B2(n_0_1_89), .ZN(n_0_1_95));
   NAND2_X1 i_0_1_165 (.A1(n_0_60), .A2(in_a[2]), .ZN(n_0_1_96));
   OAI21_X1 i_0_1_166 (.A(n_0_1_96), .B1(n_0_60), .B2(in_a[2]), .ZN(n_0_1_97));
   XNOR2_X1 i_0_1_167 (.A(n_0_1_95), .B(n_0_1_97), .ZN(n_0_193));
   INV_X1 i_0_1_168 (.A(n_0_1_96), .ZN(n_0_1_98));
   INV_X1 i_0_1_169 (.A(n_0_1_97), .ZN(n_0_1_99));
   AOI21_X1 i_0_1_170 (.A(n_0_1_98), .B1(n_0_1_95), .B2(n_0_1_99), .ZN(n_0_1_100));
   NAND2_X1 i_0_1_171 (.A1(n_0_59), .A2(in_a[3]), .ZN(n_0_1_101));
   OAI21_X1 i_0_1_172 (.A(n_0_1_101), .B1(n_0_59), .B2(in_a[3]), .ZN(n_0_1_102));
   XOR2_X1 i_0_1_173 (.A(n_0_1_100), .B(n_0_1_102), .Z(n_0_194));
   OAI21_X1 i_0_1_174 (.A(n_0_1_101), .B1(n_0_1_100), .B2(n_0_1_102), .ZN(
      n_0_1_103));
   NAND2_X1 i_0_1_175 (.A1(n_0_58), .A2(in_a[4]), .ZN(n_0_1_104));
   OAI21_X1 i_0_1_176 (.A(n_0_1_104), .B1(n_0_58), .B2(in_a[4]), .ZN(n_0_1_105));
   XNOR2_X1 i_0_1_177 (.A(n_0_1_103), .B(n_0_1_105), .ZN(n_0_195));
   INV_X1 i_0_1_178 (.A(n_0_1_104), .ZN(n_0_1_106));
   INV_X1 i_0_1_179 (.A(n_0_1_105), .ZN(n_0_1_107));
   AOI21_X1 i_0_1_180 (.A(n_0_1_106), .B1(n_0_1_103), .B2(n_0_1_107), .ZN(
      n_0_1_108));
   NAND2_X1 i_0_1_181 (.A1(n_0_57), .A2(in_a[5]), .ZN(n_0_1_109));
   OAI21_X1 i_0_1_182 (.A(n_0_1_109), .B1(n_0_57), .B2(in_a[5]), .ZN(n_0_1_110));
   XOR2_X1 i_0_1_183 (.A(n_0_1_108), .B(n_0_1_110), .Z(n_0_196));
   OAI21_X1 i_0_1_184 (.A(n_0_1_109), .B1(n_0_1_108), .B2(n_0_1_110), .ZN(
      n_0_1_111));
   NAND2_X1 i_0_1_185 (.A1(n_0_56), .A2(in_a[6]), .ZN(n_0_1_112));
   OAI21_X1 i_0_1_186 (.A(n_0_1_112), .B1(n_0_56), .B2(in_a[6]), .ZN(n_0_1_113));
   XNOR2_X1 i_0_1_187 (.A(n_0_1_111), .B(n_0_1_113), .ZN(n_0_197));
   INV_X1 i_0_1_188 (.A(n_0_1_112), .ZN(n_0_1_114));
   INV_X1 i_0_1_189 (.A(n_0_1_113), .ZN(n_0_1_115));
   AOI21_X1 i_0_1_190 (.A(n_0_1_114), .B1(n_0_1_111), .B2(n_0_1_115), .ZN(
      n_0_1_116));
   NAND2_X1 i_0_1_191 (.A1(n_0_55), .A2(in_a[7]), .ZN(n_0_1_117));
   OAI21_X1 i_0_1_192 (.A(n_0_1_117), .B1(n_0_55), .B2(in_a[7]), .ZN(n_0_1_118));
   XOR2_X1 i_0_1_193 (.A(n_0_1_116), .B(n_0_1_118), .Z(n_0_198));
   OAI21_X1 i_0_1_194 (.A(n_0_1_117), .B1(n_0_1_116), .B2(n_0_1_118), .ZN(
      n_0_1_119));
   NAND2_X1 i_0_1_195 (.A1(n_0_54), .A2(in_a[8]), .ZN(n_0_1_120));
   OAI21_X1 i_0_1_196 (.A(n_0_1_120), .B1(n_0_54), .B2(in_a[8]), .ZN(n_0_1_121));
   XNOR2_X1 i_0_1_197 (.A(n_0_1_119), .B(n_0_1_121), .ZN(n_0_199));
   INV_X1 i_0_1_198 (.A(n_0_1_120), .ZN(n_0_1_122));
   INV_X1 i_0_1_199 (.A(n_0_1_121), .ZN(n_0_1_123));
   AOI21_X1 i_0_1_200 (.A(n_0_1_122), .B1(n_0_1_119), .B2(n_0_1_123), .ZN(
      n_0_1_124));
   NAND2_X1 i_0_1_201 (.A1(n_0_53), .A2(in_a[9]), .ZN(n_0_1_125));
   OAI21_X1 i_0_1_202 (.A(n_0_1_125), .B1(n_0_53), .B2(in_a[9]), .ZN(n_0_1_126));
   XOR2_X1 i_0_1_203 (.A(n_0_1_124), .B(n_0_1_126), .Z(n_0_200));
   OAI21_X1 i_0_1_204 (.A(n_0_1_125), .B1(n_0_1_124), .B2(n_0_1_126), .ZN(
      n_0_1_127));
   NAND2_X1 i_0_1_205 (.A1(n_0_52), .A2(in_a[10]), .ZN(n_0_1_128));
   OAI21_X1 i_0_1_206 (.A(n_0_1_128), .B1(n_0_52), .B2(in_a[10]), .ZN(n_0_1_129));
   XNOR2_X1 i_0_1_207 (.A(n_0_1_127), .B(n_0_1_129), .ZN(n_0_201));
   INV_X1 i_0_1_208 (.A(n_0_1_128), .ZN(n_0_1_130));
   INV_X1 i_0_1_209 (.A(n_0_1_129), .ZN(n_0_1_131));
   AOI21_X1 i_0_1_210 (.A(n_0_1_130), .B1(n_0_1_127), .B2(n_0_1_131), .ZN(
      n_0_1_132));
   NAND2_X1 i_0_1_211 (.A1(n_0_51), .A2(in_a[11]), .ZN(n_0_1_133));
   OAI21_X1 i_0_1_212 (.A(n_0_1_133), .B1(n_0_51), .B2(in_a[11]), .ZN(n_0_1_134));
   XOR2_X1 i_0_1_213 (.A(n_0_1_132), .B(n_0_1_134), .Z(n_0_202));
   OAI21_X1 i_0_1_214 (.A(n_0_1_133), .B1(n_0_1_132), .B2(n_0_1_134), .ZN(
      n_0_1_135));
   NAND2_X1 i_0_1_215 (.A1(n_0_50), .A2(in_a[12]), .ZN(n_0_1_136));
   OAI21_X1 i_0_1_216 (.A(n_0_1_136), .B1(n_0_50), .B2(in_a[12]), .ZN(n_0_1_137));
   XNOR2_X1 i_0_1_217 (.A(n_0_1_135), .B(n_0_1_137), .ZN(n_0_203));
   INV_X1 i_0_1_218 (.A(n_0_1_136), .ZN(n_0_1_138));
   INV_X1 i_0_1_219 (.A(n_0_1_137), .ZN(n_0_1_139));
   AOI21_X1 i_0_1_220 (.A(n_0_1_138), .B1(n_0_1_135), .B2(n_0_1_139), .ZN(
      n_0_1_140));
   NAND2_X1 i_0_1_221 (.A1(n_0_49), .A2(in_a[13]), .ZN(n_0_1_141));
   OAI21_X1 i_0_1_222 (.A(n_0_1_141), .B1(n_0_49), .B2(in_a[13]), .ZN(n_0_1_142));
   XOR2_X1 i_0_1_223 (.A(n_0_1_140), .B(n_0_1_142), .Z(n_0_204));
   OAI21_X1 i_0_1_224 (.A(n_0_1_141), .B1(n_0_1_140), .B2(n_0_1_142), .ZN(
      n_0_1_143));
   NAND2_X1 i_0_1_225 (.A1(n_0_48), .A2(in_a[14]), .ZN(n_0_1_144));
   OAI21_X1 i_0_1_226 (.A(n_0_1_144), .B1(n_0_48), .B2(in_a[14]), .ZN(n_0_1_145));
   XNOR2_X1 i_0_1_227 (.A(n_0_1_143), .B(n_0_1_145), .ZN(n_0_205));
   INV_X1 i_0_1_228 (.A(n_0_1_144), .ZN(n_0_1_146));
   INV_X1 i_0_1_229 (.A(n_0_1_145), .ZN(n_0_1_147));
   AOI21_X1 i_0_1_230 (.A(n_0_1_146), .B1(n_0_1_143), .B2(n_0_1_147), .ZN(
      n_0_1_148));
   NAND2_X1 i_0_1_231 (.A1(n_0_47), .A2(in_a[15]), .ZN(n_0_1_149));
   OAI21_X1 i_0_1_232 (.A(n_0_1_149), .B1(n_0_47), .B2(in_a[15]), .ZN(n_0_1_150));
   XOR2_X1 i_0_1_233 (.A(n_0_1_148), .B(n_0_1_150), .Z(n_0_206));
   OAI21_X1 i_0_1_234 (.A(n_0_1_149), .B1(n_0_1_148), .B2(n_0_1_150), .ZN(
      n_0_1_151));
   NAND2_X1 i_0_1_235 (.A1(n_0_46), .A2(in_a[16]), .ZN(n_0_1_152));
   OAI21_X1 i_0_1_236 (.A(n_0_1_152), .B1(n_0_46), .B2(in_a[16]), .ZN(n_0_1_153));
   XNOR2_X1 i_0_1_237 (.A(n_0_1_151), .B(n_0_1_153), .ZN(n_0_207));
   INV_X1 i_0_1_238 (.A(n_0_1_152), .ZN(n_0_1_154));
   INV_X1 i_0_1_239 (.A(n_0_1_153), .ZN(n_0_1_155));
   AOI21_X1 i_0_1_240 (.A(n_0_1_154), .B1(n_0_1_151), .B2(n_0_1_155), .ZN(
      n_0_1_156));
   NAND2_X1 i_0_1_241 (.A1(n_0_45), .A2(in_a[17]), .ZN(n_0_1_157));
   OAI21_X1 i_0_1_242 (.A(n_0_1_157), .B1(n_0_45), .B2(in_a[17]), .ZN(n_0_1_158));
   XOR2_X1 i_0_1_243 (.A(n_0_1_156), .B(n_0_1_158), .Z(n_0_208));
   OAI21_X1 i_0_1_244 (.A(n_0_1_157), .B1(n_0_1_156), .B2(n_0_1_158), .ZN(
      n_0_1_159));
   NAND2_X1 i_0_1_245 (.A1(n_0_44), .A2(in_a[18]), .ZN(n_0_1_160));
   OAI21_X1 i_0_1_246 (.A(n_0_1_160), .B1(n_0_44), .B2(in_a[18]), .ZN(n_0_1_161));
   XNOR2_X1 i_0_1_247 (.A(n_0_1_159), .B(n_0_1_161), .ZN(n_0_209));
   INV_X1 i_0_1_248 (.A(n_0_1_160), .ZN(n_0_1_162));
   INV_X1 i_0_1_249 (.A(n_0_1_161), .ZN(n_0_1_163));
   AOI21_X1 i_0_1_250 (.A(n_0_1_162), .B1(n_0_1_159), .B2(n_0_1_163), .ZN(
      n_0_1_164));
   NAND2_X1 i_0_1_251 (.A1(n_0_43), .A2(in_a[19]), .ZN(n_0_1_165));
   OAI21_X1 i_0_1_252 (.A(n_0_1_165), .B1(n_0_43), .B2(in_a[19]), .ZN(n_0_1_166));
   XOR2_X1 i_0_1_253 (.A(n_0_1_164), .B(n_0_1_166), .Z(n_0_210));
   OAI21_X1 i_0_1_254 (.A(n_0_1_165), .B1(n_0_1_164), .B2(n_0_1_166), .ZN(
      n_0_1_167));
   NAND2_X1 i_0_1_255 (.A1(n_0_42), .A2(in_a[20]), .ZN(n_0_1_168));
   OAI21_X1 i_0_1_256 (.A(n_0_1_168), .B1(n_0_42), .B2(in_a[20]), .ZN(n_0_1_169));
   XNOR2_X1 i_0_1_257 (.A(n_0_1_167), .B(n_0_1_169), .ZN(n_0_211));
   INV_X1 i_0_1_258 (.A(n_0_1_168), .ZN(n_0_1_170));
   INV_X1 i_0_1_259 (.A(n_0_1_169), .ZN(n_0_1_171));
   AOI21_X1 i_0_1_260 (.A(n_0_1_170), .B1(n_0_1_167), .B2(n_0_1_171), .ZN(
      n_0_1_172));
   NAND2_X1 i_0_1_261 (.A1(n_0_41), .A2(in_a[21]), .ZN(n_0_1_173));
   OAI21_X1 i_0_1_262 (.A(n_0_1_173), .B1(n_0_41), .B2(in_a[21]), .ZN(n_0_1_174));
   XOR2_X1 i_0_1_263 (.A(n_0_1_172), .B(n_0_1_174), .Z(n_0_212));
   OAI21_X1 i_0_1_264 (.A(n_0_1_173), .B1(n_0_1_172), .B2(n_0_1_174), .ZN(
      n_0_1_175));
   NAND2_X1 i_0_1_265 (.A1(n_0_40), .A2(in_a[22]), .ZN(n_0_1_176));
   OAI21_X1 i_0_1_266 (.A(n_0_1_176), .B1(n_0_40), .B2(in_a[22]), .ZN(n_0_1_177));
   XNOR2_X1 i_0_1_267 (.A(n_0_1_175), .B(n_0_1_177), .ZN(n_0_213));
   INV_X1 i_0_1_268 (.A(n_0_1_176), .ZN(n_0_1_178));
   INV_X1 i_0_1_269 (.A(n_0_1_177), .ZN(n_0_1_179));
   AOI21_X1 i_0_1_270 (.A(n_0_1_178), .B1(n_0_1_175), .B2(n_0_1_179), .ZN(
      n_0_1_180));
   NAND2_X1 i_0_1_271 (.A1(n_0_39), .A2(in_a[23]), .ZN(n_0_1_181));
   OAI21_X1 i_0_1_272 (.A(n_0_1_181), .B1(n_0_39), .B2(in_a[23]), .ZN(n_0_1_182));
   XOR2_X1 i_0_1_273 (.A(n_0_1_180), .B(n_0_1_182), .Z(n_0_214));
   OAI21_X1 i_0_1_274 (.A(n_0_1_181), .B1(n_0_1_180), .B2(n_0_1_182), .ZN(
      n_0_1_183));
   NAND2_X1 i_0_1_275 (.A1(n_0_38), .A2(in_a[24]), .ZN(n_0_1_184));
   OAI21_X1 i_0_1_276 (.A(n_0_1_184), .B1(n_0_38), .B2(in_a[24]), .ZN(n_0_1_185));
   XNOR2_X1 i_0_1_277 (.A(n_0_1_183), .B(n_0_1_185), .ZN(n_0_215));
   INV_X1 i_0_1_278 (.A(n_0_1_184), .ZN(n_0_1_186));
   INV_X1 i_0_1_279 (.A(n_0_1_185), .ZN(n_0_1_187));
   AOI21_X1 i_0_1_280 (.A(n_0_1_186), .B1(n_0_1_183), .B2(n_0_1_187), .ZN(
      n_0_1_188));
   NAND2_X1 i_0_1_281 (.A1(n_0_37), .A2(in_a[25]), .ZN(n_0_1_189));
   OAI21_X1 i_0_1_282 (.A(n_0_1_189), .B1(n_0_37), .B2(in_a[25]), .ZN(n_0_1_190));
   XOR2_X1 i_0_1_283 (.A(n_0_1_188), .B(n_0_1_190), .Z(n_0_216));
   OAI21_X1 i_0_1_284 (.A(n_0_1_189), .B1(n_0_1_188), .B2(n_0_1_190), .ZN(
      n_0_1_191));
   NAND2_X1 i_0_1_285 (.A1(n_0_36), .A2(in_a[26]), .ZN(n_0_1_192));
   OAI21_X1 i_0_1_286 (.A(n_0_1_192), .B1(n_0_36), .B2(in_a[26]), .ZN(n_0_1_193));
   XNOR2_X1 i_0_1_287 (.A(n_0_1_191), .B(n_0_1_193), .ZN(n_0_217));
   INV_X1 i_0_1_288 (.A(n_0_1_192), .ZN(n_0_1_194));
   INV_X1 i_0_1_289 (.A(n_0_1_193), .ZN(n_0_1_195));
   AOI21_X1 i_0_1_290 (.A(n_0_1_194), .B1(n_0_1_191), .B2(n_0_1_195), .ZN(
      n_0_1_196));
   NAND2_X1 i_0_1_291 (.A1(n_0_35), .A2(in_a[27]), .ZN(n_0_1_197));
   OAI21_X1 i_0_1_292 (.A(n_0_1_197), .B1(n_0_35), .B2(in_a[27]), .ZN(n_0_1_198));
   XOR2_X1 i_0_1_293 (.A(n_0_1_196), .B(n_0_1_198), .Z(n_0_218));
   OAI21_X1 i_0_1_294 (.A(n_0_1_197), .B1(n_0_1_196), .B2(n_0_1_198), .ZN(
      n_0_1_199));
   NAND2_X1 i_0_1_295 (.A1(n_0_34), .A2(in_a[28]), .ZN(n_0_1_200));
   OAI21_X1 i_0_1_296 (.A(n_0_1_200), .B1(n_0_34), .B2(in_a[28]), .ZN(n_0_1_201));
   XNOR2_X1 i_0_1_297 (.A(n_0_1_199), .B(n_0_1_201), .ZN(n_0_219));
   INV_X1 i_0_1_298 (.A(n_0_1_200), .ZN(n_0_1_202));
   INV_X1 i_0_1_299 (.A(n_0_1_201), .ZN(n_0_1_203));
   AOI21_X1 i_0_1_300 (.A(n_0_1_202), .B1(n_0_1_199), .B2(n_0_1_203), .ZN(
      n_0_1_204));
   NAND2_X1 i_0_1_301 (.A1(n_0_33), .A2(in_a[29]), .ZN(n_0_1_205));
   OAI21_X1 i_0_1_302 (.A(n_0_1_205), .B1(n_0_33), .B2(in_a[29]), .ZN(n_0_1_206));
   XOR2_X1 i_0_1_303 (.A(n_0_1_204), .B(n_0_1_206), .Z(n_0_220));
   OAI21_X1 i_0_1_304 (.A(n_0_1_205), .B1(n_0_1_204), .B2(n_0_1_206), .ZN(
      n_0_1_207));
   NAND2_X1 i_0_1_305 (.A1(n_0_32), .A2(in_a[30]), .ZN(n_0_1_208));
   OAI21_X1 i_0_1_306 (.A(n_0_1_208), .B1(n_0_32), .B2(in_a[30]), .ZN(n_0_1_209));
   XNOR2_X1 i_0_1_307 (.A(n_0_1_207), .B(n_0_1_209), .ZN(n_0_221));
   INV_X1 i_0_1_308 (.A(n_0_1_208), .ZN(n_0_1_210));
   INV_X1 i_0_1_309 (.A(n_0_1_209), .ZN(n_0_1_211));
   AOI21_X1 i_0_1_310 (.A(n_0_1_210), .B1(n_0_1_207), .B2(n_0_1_211), .ZN(
      n_0_1_212));
   NAND2_X1 i_0_1_311 (.A1(n_0_31), .A2(in_a[31]), .ZN(n_0_1_213));
   OAI21_X1 i_0_1_312 (.A(n_0_1_213), .B1(n_0_31), .B2(in_a[31]), .ZN(n_0_1_214));
   XOR2_X1 i_0_1_313 (.A(n_0_1_212), .B(n_0_1_214), .Z(n_0_222));
   OAI21_X1 i_0_1_314 (.A(n_0_1_213), .B1(n_0_1_212), .B2(n_0_1_214), .ZN(
      n_0_1_215));
   NAND2_X1 i_0_1_315 (.A1(n_0_30), .A2(in_a[32]), .ZN(n_0_1_216));
   OAI21_X1 i_0_1_316 (.A(n_0_1_216), .B1(n_0_30), .B2(in_a[32]), .ZN(n_0_1_217));
   XNOR2_X1 i_0_1_317 (.A(n_0_1_215), .B(n_0_1_217), .ZN(n_0_223));
   INV_X1 i_0_1_318 (.A(n_0_1_216), .ZN(n_0_1_218));
   INV_X1 i_0_1_319 (.A(n_0_1_217), .ZN(n_0_1_219));
   AOI21_X1 i_0_1_320 (.A(n_0_1_218), .B1(n_0_1_215), .B2(n_0_1_219), .ZN(
      n_0_1_220));
   NAND2_X1 i_0_1_321 (.A1(n_0_29), .A2(in_a[33]), .ZN(n_0_1_221));
   OAI21_X1 i_0_1_322 (.A(n_0_1_221), .B1(n_0_29), .B2(in_a[33]), .ZN(n_0_1_222));
   XOR2_X1 i_0_1_323 (.A(n_0_1_220), .B(n_0_1_222), .Z(n_0_224));
   OAI21_X1 i_0_1_324 (.A(n_0_1_221), .B1(n_0_1_220), .B2(n_0_1_222), .ZN(
      n_0_1_223));
   NAND2_X1 i_0_1_325 (.A1(n_0_28), .A2(in_a[34]), .ZN(n_0_1_224));
   OAI21_X1 i_0_1_326 (.A(n_0_1_224), .B1(n_0_28), .B2(in_a[34]), .ZN(n_0_1_225));
   XNOR2_X1 i_0_1_327 (.A(n_0_1_223), .B(n_0_1_225), .ZN(n_0_225));
   INV_X1 i_0_1_328 (.A(n_0_1_224), .ZN(n_0_1_226));
   INV_X1 i_0_1_329 (.A(n_0_1_225), .ZN(n_0_1_227));
   AOI21_X1 i_0_1_330 (.A(n_0_1_226), .B1(n_0_1_223), .B2(n_0_1_227), .ZN(
      n_0_1_228));
   NAND2_X1 i_0_1_331 (.A1(n_0_27), .A2(in_a[35]), .ZN(n_0_1_229));
   OAI21_X1 i_0_1_332 (.A(n_0_1_229), .B1(n_0_27), .B2(in_a[35]), .ZN(n_0_1_230));
   XOR2_X1 i_0_1_333 (.A(n_0_1_228), .B(n_0_1_230), .Z(n_0_226));
   OAI21_X1 i_0_1_334 (.A(n_0_1_229), .B1(n_0_1_228), .B2(n_0_1_230), .ZN(
      n_0_1_231));
   NAND2_X1 i_0_1_335 (.A1(n_0_26), .A2(in_a[36]), .ZN(n_0_1_232));
   OAI21_X1 i_0_1_336 (.A(n_0_1_232), .B1(n_0_26), .B2(in_a[36]), .ZN(n_0_1_233));
   XNOR2_X1 i_0_1_337 (.A(n_0_1_231), .B(n_0_1_233), .ZN(n_0_227));
   INV_X1 i_0_1_338 (.A(n_0_1_232), .ZN(n_0_1_234));
   INV_X1 i_0_1_339 (.A(n_0_1_233), .ZN(n_0_1_235));
   AOI21_X1 i_0_1_340 (.A(n_0_1_234), .B1(n_0_1_231), .B2(n_0_1_235), .ZN(
      n_0_1_236));
   NAND2_X1 i_0_1_341 (.A1(n_0_25), .A2(in_a[37]), .ZN(n_0_1_237));
   OAI21_X1 i_0_1_342 (.A(n_0_1_237), .B1(n_0_25), .B2(in_a[37]), .ZN(n_0_1_238));
   XOR2_X1 i_0_1_343 (.A(n_0_1_236), .B(n_0_1_238), .Z(n_0_228));
   OAI21_X1 i_0_1_344 (.A(n_0_1_237), .B1(n_0_1_236), .B2(n_0_1_238), .ZN(
      n_0_1_239));
   NAND2_X1 i_0_1_345 (.A1(n_0_24), .A2(in_a[38]), .ZN(n_0_1_240));
   OAI21_X1 i_0_1_346 (.A(n_0_1_240), .B1(n_0_24), .B2(in_a[38]), .ZN(n_0_1_241));
   XNOR2_X1 i_0_1_347 (.A(n_0_1_239), .B(n_0_1_241), .ZN(n_0_229));
   INV_X1 i_0_1_348 (.A(n_0_1_240), .ZN(n_0_1_242));
   INV_X1 i_0_1_349 (.A(n_0_1_241), .ZN(n_0_1_243));
   AOI21_X1 i_0_1_350 (.A(n_0_1_242), .B1(n_0_1_239), .B2(n_0_1_243), .ZN(
      n_0_1_244));
   NAND2_X1 i_0_1_351 (.A1(n_0_23), .A2(in_a[39]), .ZN(n_0_1_245));
   OAI21_X1 i_0_1_352 (.A(n_0_1_245), .B1(n_0_23), .B2(in_a[39]), .ZN(n_0_1_246));
   XOR2_X1 i_0_1_353 (.A(n_0_1_244), .B(n_0_1_246), .Z(n_0_230));
   OAI21_X1 i_0_1_354 (.A(n_0_1_245), .B1(n_0_1_244), .B2(n_0_1_246), .ZN(
      n_0_1_247));
   NAND2_X1 i_0_1_355 (.A1(n_0_22), .A2(in_a[40]), .ZN(n_0_1_248));
   OAI21_X1 i_0_1_356 (.A(n_0_1_248), .B1(n_0_22), .B2(in_a[40]), .ZN(n_0_1_249));
   XNOR2_X1 i_0_1_357 (.A(n_0_1_247), .B(n_0_1_249), .ZN(n_0_231));
   INV_X1 i_0_1_358 (.A(n_0_1_248), .ZN(n_0_1_250));
   INV_X1 i_0_1_359 (.A(n_0_1_249), .ZN(n_0_1_251));
   AOI21_X1 i_0_1_360 (.A(n_0_1_250), .B1(n_0_1_247), .B2(n_0_1_251), .ZN(
      n_0_1_252));
   NAND2_X1 i_0_1_361 (.A1(n_0_21), .A2(in_a[41]), .ZN(n_0_1_253));
   OAI21_X1 i_0_1_362 (.A(n_0_1_253), .B1(n_0_21), .B2(in_a[41]), .ZN(n_0_1_254));
   XOR2_X1 i_0_1_363 (.A(n_0_1_252), .B(n_0_1_254), .Z(n_0_232));
   OAI21_X1 i_0_1_364 (.A(n_0_1_253), .B1(n_0_1_252), .B2(n_0_1_254), .ZN(
      n_0_1_255));
   NAND2_X1 i_0_1_365 (.A1(n_0_20), .A2(in_a[42]), .ZN(n_0_1_256));
   OAI21_X1 i_0_1_366 (.A(n_0_1_256), .B1(n_0_20), .B2(in_a[42]), .ZN(n_0_1_257));
   XNOR2_X1 i_0_1_367 (.A(n_0_1_255), .B(n_0_1_257), .ZN(n_0_233));
   INV_X1 i_0_1_368 (.A(n_0_1_256), .ZN(n_0_1_258));
   INV_X1 i_0_1_369 (.A(n_0_1_257), .ZN(n_0_1_259));
   AOI21_X1 i_0_1_370 (.A(n_0_1_258), .B1(n_0_1_255), .B2(n_0_1_259), .ZN(
      n_0_1_260));
   NAND2_X1 i_0_1_371 (.A1(n_0_19), .A2(in_a[43]), .ZN(n_0_1_261));
   OAI21_X1 i_0_1_372 (.A(n_0_1_261), .B1(n_0_19), .B2(in_a[43]), .ZN(n_0_1_262));
   XOR2_X1 i_0_1_373 (.A(n_0_1_260), .B(n_0_1_262), .Z(n_0_234));
   OAI21_X1 i_0_1_374 (.A(n_0_1_261), .B1(n_0_1_260), .B2(n_0_1_262), .ZN(
      n_0_1_263));
   NAND2_X1 i_0_1_375 (.A1(n_0_18), .A2(in_a[44]), .ZN(n_0_1_264));
   OAI21_X1 i_0_1_376 (.A(n_0_1_264), .B1(n_0_18), .B2(in_a[44]), .ZN(n_0_1_265));
   XNOR2_X1 i_0_1_377 (.A(n_0_1_263), .B(n_0_1_265), .ZN(n_0_235));
   INV_X1 i_0_1_378 (.A(n_0_1_264), .ZN(n_0_1_266));
   INV_X1 i_0_1_379 (.A(n_0_1_265), .ZN(n_0_1_267));
   AOI21_X1 i_0_1_380 (.A(n_0_1_266), .B1(n_0_1_263), .B2(n_0_1_267), .ZN(
      n_0_1_268));
   NAND2_X1 i_0_1_381 (.A1(n_0_17), .A2(in_a[45]), .ZN(n_0_1_269));
   OAI21_X1 i_0_1_382 (.A(n_0_1_269), .B1(n_0_17), .B2(in_a[45]), .ZN(n_0_1_270));
   XOR2_X1 i_0_1_383 (.A(n_0_1_268), .B(n_0_1_270), .Z(n_0_236));
   OAI21_X1 i_0_1_384 (.A(n_0_1_269), .B1(n_0_1_268), .B2(n_0_1_270), .ZN(
      n_0_1_271));
   NAND2_X1 i_0_1_385 (.A1(n_0_16), .A2(in_a[46]), .ZN(n_0_1_272));
   OAI21_X1 i_0_1_386 (.A(n_0_1_272), .B1(n_0_16), .B2(in_a[46]), .ZN(n_0_1_273));
   XNOR2_X1 i_0_1_387 (.A(n_0_1_271), .B(n_0_1_273), .ZN(n_0_237));
   INV_X1 i_0_1_388 (.A(n_0_1_272), .ZN(n_0_1_274));
   INV_X1 i_0_1_389 (.A(n_0_1_273), .ZN(n_0_1_275));
   AOI21_X1 i_0_1_390 (.A(n_0_1_274), .B1(n_0_1_271), .B2(n_0_1_275), .ZN(
      n_0_1_276));
   NAND2_X1 i_0_1_391 (.A1(n_0_15), .A2(in_a[47]), .ZN(n_0_1_277));
   OAI21_X1 i_0_1_392 (.A(n_0_1_277), .B1(n_0_15), .B2(in_a[47]), .ZN(n_0_1_278));
   XOR2_X1 i_0_1_393 (.A(n_0_1_276), .B(n_0_1_278), .Z(n_0_238));
   OAI21_X1 i_0_1_394 (.A(n_0_1_277), .B1(n_0_1_276), .B2(n_0_1_278), .ZN(
      n_0_1_279));
   NAND2_X1 i_0_1_395 (.A1(n_0_14), .A2(in_a[48]), .ZN(n_0_1_280));
   OAI21_X1 i_0_1_396 (.A(n_0_1_280), .B1(n_0_14), .B2(in_a[48]), .ZN(n_0_1_281));
   XNOR2_X1 i_0_1_397 (.A(n_0_1_279), .B(n_0_1_281), .ZN(n_0_239));
   INV_X1 i_0_1_398 (.A(n_0_1_280), .ZN(n_0_1_282));
   INV_X1 i_0_1_399 (.A(n_0_1_281), .ZN(n_0_1_283));
   AOI21_X1 i_0_1_400 (.A(n_0_1_282), .B1(n_0_1_279), .B2(n_0_1_283), .ZN(
      n_0_1_284));
   NAND2_X1 i_0_1_401 (.A1(n_0_13), .A2(in_a[49]), .ZN(n_0_1_285));
   OAI21_X1 i_0_1_402 (.A(n_0_1_285), .B1(n_0_13), .B2(in_a[49]), .ZN(n_0_1_286));
   XOR2_X1 i_0_1_403 (.A(n_0_1_284), .B(n_0_1_286), .Z(n_0_240));
   OAI21_X1 i_0_1_404 (.A(n_0_1_285), .B1(n_0_1_284), .B2(n_0_1_286), .ZN(
      n_0_1_287));
   NAND2_X1 i_0_1_405 (.A1(n_0_12), .A2(in_a[50]), .ZN(n_0_1_288));
   OAI21_X1 i_0_1_406 (.A(n_0_1_288), .B1(n_0_12), .B2(in_a[50]), .ZN(n_0_1_289));
   XNOR2_X1 i_0_1_407 (.A(n_0_1_287), .B(n_0_1_289), .ZN(n_0_241));
   INV_X1 i_0_1_408 (.A(n_0_1_288), .ZN(n_0_1_290));
   INV_X1 i_0_1_409 (.A(n_0_1_289), .ZN(n_0_1_291));
   AOI21_X1 i_0_1_410 (.A(n_0_1_290), .B1(n_0_1_287), .B2(n_0_1_291), .ZN(
      n_0_1_292));
   NAND2_X1 i_0_1_411 (.A1(n_0_11), .A2(in_a[51]), .ZN(n_0_1_293));
   OAI21_X1 i_0_1_412 (.A(n_0_1_293), .B1(n_0_11), .B2(in_a[51]), .ZN(n_0_1_294));
   XOR2_X1 i_0_1_413 (.A(n_0_1_292), .B(n_0_1_294), .Z(n_0_242));
   OAI21_X1 i_0_1_414 (.A(n_0_1_293), .B1(n_0_1_292), .B2(n_0_1_294), .ZN(
      n_0_1_295));
   NAND2_X1 i_0_1_415 (.A1(n_0_10), .A2(in_a[52]), .ZN(n_0_1_296));
   OAI21_X1 i_0_1_416 (.A(n_0_1_296), .B1(n_0_10), .B2(in_a[52]), .ZN(n_0_1_297));
   XNOR2_X1 i_0_1_417 (.A(n_0_1_295), .B(n_0_1_297), .ZN(n_0_243));
   INV_X1 i_0_1_418 (.A(n_0_1_296), .ZN(n_0_1_298));
   INV_X1 i_0_1_419 (.A(n_0_1_297), .ZN(n_0_1_299));
   AOI21_X1 i_0_1_420 (.A(n_0_1_298), .B1(n_0_1_295), .B2(n_0_1_299), .ZN(
      n_0_1_300));
   NAND2_X1 i_0_1_421 (.A1(n_0_9), .A2(in_a[53]), .ZN(n_0_1_301));
   OAI21_X1 i_0_1_422 (.A(n_0_1_301), .B1(n_0_9), .B2(in_a[53]), .ZN(n_0_1_302));
   XOR2_X1 i_0_1_423 (.A(n_0_1_300), .B(n_0_1_302), .Z(n_0_244));
   OAI21_X1 i_0_1_424 (.A(n_0_1_301), .B1(n_0_1_300), .B2(n_0_1_302), .ZN(
      n_0_1_303));
   NAND2_X1 i_0_1_425 (.A1(n_0_8), .A2(in_a[54]), .ZN(n_0_1_304));
   OAI21_X1 i_0_1_426 (.A(n_0_1_304), .B1(n_0_8), .B2(in_a[54]), .ZN(n_0_1_305));
   XNOR2_X1 i_0_1_427 (.A(n_0_1_303), .B(n_0_1_305), .ZN(n_0_245));
   INV_X1 i_0_1_428 (.A(n_0_1_304), .ZN(n_0_1_306));
   INV_X1 i_0_1_429 (.A(n_0_1_305), .ZN(n_0_1_307));
   AOI21_X1 i_0_1_430 (.A(n_0_1_306), .B1(n_0_1_303), .B2(n_0_1_307), .ZN(
      n_0_1_308));
   NAND2_X1 i_0_1_431 (.A1(n_0_7), .A2(in_a[55]), .ZN(n_0_1_309));
   OAI21_X1 i_0_1_432 (.A(n_0_1_309), .B1(n_0_7), .B2(in_a[55]), .ZN(n_0_1_310));
   XOR2_X1 i_0_1_433 (.A(n_0_1_308), .B(n_0_1_310), .Z(n_0_246));
   OAI21_X1 i_0_1_434 (.A(n_0_1_309), .B1(n_0_1_308), .B2(n_0_1_310), .ZN(
      n_0_1_311));
   NAND2_X1 i_0_1_435 (.A1(n_0_6), .A2(in_a[56]), .ZN(n_0_1_312));
   OAI21_X1 i_0_1_436 (.A(n_0_1_312), .B1(n_0_6), .B2(in_a[56]), .ZN(n_0_1_313));
   XNOR2_X1 i_0_1_437 (.A(n_0_1_311), .B(n_0_1_313), .ZN(n_0_247));
   INV_X1 i_0_1_438 (.A(n_0_1_312), .ZN(n_0_1_314));
   INV_X1 i_0_1_439 (.A(n_0_1_313), .ZN(n_0_1_315));
   AOI21_X1 i_0_1_440 (.A(n_0_1_314), .B1(n_0_1_311), .B2(n_0_1_315), .ZN(
      n_0_1_316));
   NAND2_X1 i_0_1_441 (.A1(n_0_5), .A2(in_a[57]), .ZN(n_0_1_317));
   OAI21_X1 i_0_1_442 (.A(n_0_1_317), .B1(n_0_5), .B2(in_a[57]), .ZN(n_0_1_318));
   XOR2_X1 i_0_1_443 (.A(n_0_1_316), .B(n_0_1_318), .Z(n_0_248));
   OAI21_X1 i_0_1_444 (.A(n_0_1_317), .B1(n_0_1_316), .B2(n_0_1_318), .ZN(
      n_0_1_319));
   NAND2_X1 i_0_1_445 (.A1(n_0_4), .A2(in_a[58]), .ZN(n_0_1_320));
   OAI21_X1 i_0_1_446 (.A(n_0_1_320), .B1(n_0_4), .B2(in_a[58]), .ZN(n_0_1_321));
   XNOR2_X1 i_0_1_447 (.A(n_0_1_319), .B(n_0_1_321), .ZN(n_0_249));
   INV_X1 i_0_1_448 (.A(n_0_1_320), .ZN(n_0_1_322));
   INV_X1 i_0_1_449 (.A(n_0_1_321), .ZN(n_0_1_323));
   AOI21_X1 i_0_1_450 (.A(n_0_1_322), .B1(n_0_1_319), .B2(n_0_1_323), .ZN(
      n_0_1_324));
   NAND2_X1 i_0_1_451 (.A1(n_0_3), .A2(in_a[59]), .ZN(n_0_1_325));
   OAI21_X1 i_0_1_452 (.A(n_0_1_325), .B1(n_0_3), .B2(in_a[59]), .ZN(n_0_1_326));
   XOR2_X1 i_0_1_453 (.A(n_0_1_324), .B(n_0_1_326), .Z(n_0_250));
   OAI21_X1 i_0_1_454 (.A(n_0_1_325), .B1(n_0_1_324), .B2(n_0_1_326), .ZN(
      n_0_1_327));
   NAND2_X1 i_0_1_455 (.A1(n_0_2), .A2(in_a[60]), .ZN(n_0_1_328));
   OAI21_X1 i_0_1_456 (.A(n_0_1_328), .B1(n_0_2), .B2(in_a[60]), .ZN(n_0_1_329));
   XNOR2_X1 i_0_1_457 (.A(n_0_1_327), .B(n_0_1_329), .ZN(n_0_251));
   INV_X1 i_0_1_458 (.A(n_0_1_328), .ZN(n_0_1_330));
   INV_X1 i_0_1_459 (.A(n_0_1_329), .ZN(n_0_1_331));
   AOI21_X1 i_0_1_460 (.A(n_0_1_330), .B1(n_0_1_327), .B2(n_0_1_331), .ZN(
      n_0_1_332));
   NAND2_X1 i_0_1_461 (.A1(n_0_1), .A2(in_a[61]), .ZN(n_0_1_333));
   OAI21_X1 i_0_1_462 (.A(n_0_1_333), .B1(n_0_1), .B2(in_a[61]), .ZN(n_0_1_334));
   XOR2_X1 i_0_1_463 (.A(n_0_1_332), .B(n_0_1_334), .Z(n_0_252));
   OAI21_X1 i_0_1_464 (.A(n_0_1_333), .B1(n_0_1_332), .B2(n_0_1_334), .ZN(
      n_0_1_335));
   NAND2_X1 i_0_1_465 (.A1(n_0_0), .A2(in_a[62]), .ZN(n_0_1_336));
   OAI21_X1 i_0_1_466 (.A(n_0_1_336), .B1(n_0_0), .B2(in_a[62]), .ZN(n_0_1_337));
   XNOR2_X1 i_0_1_467 (.A(n_0_1_335), .B(n_0_1_337), .ZN(n_0_253));
   INV_X1 i_0_1_468 (.A(n_0_1_336), .ZN(n_0_1_338));
   INV_X1 i_0_1_469 (.A(n_0_1_337), .ZN(n_0_1_339));
   AOI21_X1 i_0_1_470 (.A(n_0_1_338), .B1(n_0_1_335), .B2(n_0_1_339), .ZN(
      n_0_1_340));
   XNOR2_X1 i_0_1_471 (.A(n_0_1_340), .B(n_0_1_67), .ZN(n_0_254));
   BUF_X1 rt_shieldBuf__1 (.A(done), .Z(n_0_255));
endmodule
