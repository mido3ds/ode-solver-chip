/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sat Apr 25 20:22:51 2020
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 1629102782 */

module half_adder__3_147(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   INV_X1 i_2 (.A(a), .ZN(f));
endmodule

module half_adder__3_144(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_141(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_138(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_135(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_132(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_129(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   XOR2_X1 i_1_0 (.A(a), .B(b), .Z(f));
endmodule

module incrementor__3_148(a, enbl, c);
   input [6:0]a;
   input enbl;
   output [6:0]c;

   half_adder__3_147 half_adder_0_0_half_adder_0_i (.a(a[0]), .b(), .cout(), 
      .f(c[0]));
   half_adder__3_144 half_adder_0_1_half_adder_0_i (.a(a[1]), .b(a[0]), .cout(
      n_0), .f(c[1]));
   half_adder__3_141 half_adder_0_2_half_adder_0_i (.a(a[2]), .b(n_0), .cout(n_1), 
      .f(c[2]));
   half_adder__3_138 half_adder_0_3_half_adder_0_i (.a(a[3]), .b(n_1), .cout(n_2), 
      .f(c[3]));
   half_adder__3_135 half_adder_0_4_half_adder_0_i (.a(a[4]), .b(n_2), .cout(n_3), 
      .f(c[4]));
   half_adder__3_132 half_adder_0_5_half_adder_0_i (.a(a[5]), .b(n_3), .cout(n_4), 
      .f(c[5]));
   half_adder__3_129 half_adder_0_6_half_adder_0_i (.a(a[6]), .b(n_4), .cout(), 
      .f(c[6]));
endmodule

module full_adder__3_125(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;

   INV_X1 i_0_0 (.A(n_0_4), .ZN(cout));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(f));
   NAND2_X1 i_0_2 (.A1(n_0_1), .A2(n_0_4), .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(n_0_3), .A2(n_0_2), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(a), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(b), .ZN(n_0_3));
   NAND2_X1 i_0_6 (.A1(b), .A2(a), .ZN(n_0_4));
endmodule

module full_adder__3_121(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;

   NAND2_X1 i_0_0 (.A1(n_0_3), .A2(n_0_9), .ZN(cout));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(f));
   NAND2_X1 i_0_2 (.A1(n_0_1), .A2(n_0_3), .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(n_0_2), .A2(n_0_5), .ZN(n_0_1));
   INV_X1 i_0_4 (.A(cin), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(cin), .A2(n_0_4), .ZN(n_0_3));
   INV_X1 i_0_6 (.A(n_0_5), .ZN(n_0_4));
   NAND2_X1 i_0_7 (.A1(n_0_6), .A2(n_0_9), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(n_0_8), .A2(n_0_7), .ZN(n_0_6));
   INV_X1 i_0_9 (.A(a), .ZN(n_0_7));
   INV_X1 i_0_10 (.A(b), .ZN(n_0_8));
   NAND2_X1 i_0_11 (.A1(b), .A2(a), .ZN(n_0_9));
endmodule

module full_adder__3_117(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_2;
   wire n_0_3;
   wire n_0_1;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(cin), .B1(a), .B2(b), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
   INV_X1 i_0_0 (.A(n_0_2), .ZN(f));
   NAND2_X1 i_0_1 (.A1(n_0_4), .A2(n_0_3), .ZN(n_0_2));
   NAND2_X1 i_0_4 (.A1(cin), .A2(n_0_1), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(n_0_5), .ZN(n_0_1));
   NAND2_X1 i_0_6 (.A1(n_0_6), .A2(n_0_5), .ZN(n_0_4));
   XNOR2_X1 i_0_7 (.A(b), .B(a), .ZN(n_0_5));
   INV_X1 i_0_8 (.A(cin), .ZN(n_0_6));
endmodule

module full_adder__3_113(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__3_109(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__3_105(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__3_101(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
endmodule

module int_adder__3_126(a, b, cin, enbl, c, cout);
   input [6:0]a;
   input [2:0]b;
   input cin;
   input enbl;
   output [6:0]c;
   output cout;

   full_adder__3_125 full_adder_0_0_full_adder_0_i (.a(a[0]), .b(b[0]), .cin(), 
      .f(c[0]), .cout(n_0));
   full_adder__3_121 full_adder_0_1_full_adder_0_i (.a(a[1]), .b(b[1]), .cin(n_0), 
      .f(c[1]), .cout(n_1));
   full_adder__3_117 full_adder_0_2_full_adder_0_i (.a(a[2]), .b(b[2]), .cin(n_1), 
      .f(c[2]), .cout(n_2));
   full_adder__3_113 full_adder_0_3_full_adder_0_i (.a(a[3]), .b(), .cin(n_2), 
      .f(c[3]), .cout(n_3));
   full_adder__3_109 full_adder_0_4_full_adder_0_i (.a(a[4]), .b(), .cin(n_3), 
      .f(c[4]), .cout(n_4));
   full_adder__3_105 full_adder_0_5_full_adder_0_i (.a(a[5]), .b(), .cin(n_4), 
      .f(c[5]), .cout(n_5));
   full_adder__3_101 full_adder_0_6_full_adder_0_i (.a(a[6]), .b(), .cin(n_5), 
      .f(c[6]), .cout());
endmodule

module range_extractor__3_149(in_a, in_size, out_a, out_b);
   input [6:0]in_a;
   input [2:0]in_size;
   output [6:0]out_a;
   output [6:0]out_b;

   incrementor__3_148 inc (.a(in_a), .enbl(), .c(out_a));
   int_adder__3_126 add (.a(out_a), .b(in_size), .cin(), .enbl(), .c(out_b), 
      .cout());
endmodule

module full_adder__3_79(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   INV_X1 i_3 (.A(a), .ZN(f));
endmodule

module full_adder(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
endmodule

module int_adder__parameterized0(a, b, cin, enbl, c, cout);
   input [6:0]a;
   input [5:0]b;
   input cin;
   input enbl;
   output [6:0]c;
   output cout;

   full_adder__3_79 full_adder_0_5_full_adder_0_i (.a(a[5]), .b(), .cin(), 
      .f(c[5]), .cout());
   full_adder full_adder_0_6_full_adder_0_i (.a(a[6]), .b(), .cin(a[5]), 
      .f(c[6]), .cout());
endmodule

module full_adder__3_51(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XNOR2_X1 i_0_0 (.A(b), .B(a), .ZN(f));
   OR2_X1 i_0_1 (.A1(b), .A2(a), .ZN(cout));
endmodule

module full_adder__3_55(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(n_0_0));
   XOR2_X1 i_0_1 (.A(n_0_0), .B(cin), .Z(f));
endmodule

module int_adder__parameterized1(a, b, cin, enbl, c, cout);
   input [6:0]a;
   input [6:0]b;
   input cin;
   input enbl;
   output [6:0]c;
   output cout;

   full_adder__3_51 full_adder_0_5_full_adder_0_i (.a(a[5]), .b(b[5]), .cin(), 
      .f(c[5]), .cout(n_0));
   full_adder__3_55 full_adder_0_6_full_adder_0_i (.a(a[6]), .b(b[6]), .cin(n_0), 
      .f(c[6]), .cout());
endmodule

module half_adder__3_199(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   INV_X1 i_2 (.A(a), .ZN(f));
endmodule

module half_adder__3_196(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;

   INV_X1 i_0_0 (.A(n_0_0), .ZN(f));
   NAND2_X1 i_0_1 (.A1(n_0_1), .A2(n_0_4), .ZN(n_0_0));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(n_0_3), .ZN(n_0_1));
   INV_X1 i_0_3 (.A(a), .ZN(n_0_2));
   INV_X1 i_0_4 (.A(b), .ZN(n_0_3));
   INV_X1 i_0_5 (.A(n_0_4), .ZN(cout));
   NAND2_X1 i_0_6 (.A1(a), .A2(b), .ZN(n_0_4));
endmodule

module half_adder__3_193(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   INV_X1 i_0_1 (.A(n_0_0), .ZN(f));
   NAND2_X1 i_0_2 (.A1(n_0_2), .A2(n_0_1), .ZN(n_0_0));
   NAND2_X1 i_0_3 (.A1(a), .A2(b), .ZN(n_0_1));
   NAND2_X1 i_0_4 (.A1(n_0_3), .A2(n_0_4), .ZN(n_0_2));
   INV_X1 i_0_5 (.A(a), .ZN(n_0_3));
   INV_X1 i_0_6 (.A(b), .ZN(n_0_4));
endmodule

module half_adder__3_190(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_187(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_184(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_181(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   XOR2_X1 i_1_0 (.A(a), .B(b), .Z(f));
endmodule

module incrementor__3_200(a, enbl, c);
   input [6:0]a;
   input enbl;
   output [6:0]c;

   half_adder__3_199 half_adder_0_0_half_adder_0_i (.a(a[0]), .b(), .cout(), 
      .f(c[0]));
   half_adder__3_196 half_adder_0_1_half_adder_0_i (.a(a[1]), .b(a[0]), .cout(
      n_0), .f(c[1]));
   half_adder__3_193 half_adder_0_2_half_adder_0_i (.a(a[2]), .b(n_0), .cout(n_1), 
      .f(c[2]));
   half_adder__3_190 half_adder_0_3_half_adder_0_i (.a(a[3]), .b(n_1), .cout(n_2), 
      .f(c[3]));
   half_adder__3_187 half_adder_0_4_half_adder_0_i (.a(a[4]), .b(n_2), .cout(n_3), 
      .f(c[4]));
   half_adder__3_184 half_adder_0_5_half_adder_0_i (.a(a[5]), .b(n_3), .cout(n_4), 
      .f(c[5]));
   half_adder__3_181 half_adder_0_6_half_adder_0_i (.a(a[6]), .b(n_4), .cout(), 
      .f(c[6]));
endmodule

module full_adder__3_177(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(f));
   AND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(cout));
endmodule

module full_adder__3_173(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;

   NAND2_X1 i_0_0 (.A1(n_0_2), .A2(n_0_6), .ZN(cout));
   NOR2_X1 i_0_1 (.A1(n_0_1), .A2(n_0_0), .ZN(f));
   AOI21_X1 i_0_2 (.A(cin), .B1(n_0_3), .B2(n_0_6), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_2), .ZN(n_0_1));
   NAND3_X1 i_0_4 (.A1(n_0_3), .A2(cin), .A3(n_0_6), .ZN(n_0_2));
   NAND2_X1 i_0_5 (.A1(n_0_4), .A2(n_0_5), .ZN(n_0_3));
   INV_X1 i_0_6 (.A(a), .ZN(n_0_4));
   INV_X1 i_0_7 (.A(b), .ZN(n_0_5));
   NAND2_X1 i_0_8 (.A1(a), .A2(b), .ZN(n_0_6));
endmodule

module full_adder__3_169(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(f));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(cin), .B1(a), .B2(b), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module full_adder__3_165(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__3_161(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__3_157(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__3_153(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
endmodule

module int_adder__3_178(a, b, cin, enbl, c, cout);
   input [6:0]a;
   input [2:0]b;
   input cin;
   input enbl;
   output [6:0]c;
   output cout;

   full_adder__3_177 full_adder_0_0_full_adder_0_i (.a(a[0]), .b(b[0]), .cin(), 
      .f(c[0]), .cout(n_0));
   full_adder__3_173 full_adder_0_1_full_adder_0_i (.a(a[1]), .b(b[1]), .cin(n_0), 
      .f(c[1]), .cout(n_1));
   full_adder__3_169 full_adder_0_2_full_adder_0_i (.a(a[2]), .b(b[2]), .cin(n_1), 
      .f(c[2]), .cout(n_2));
   full_adder__3_165 full_adder_0_3_full_adder_0_i (.a(a[3]), .b(), .cin(n_2), 
      .f(c[3]), .cout(n_3));
   full_adder__3_161 full_adder_0_4_full_adder_0_i (.a(a[4]), .b(), .cin(n_3), 
      .f(c[4]), .cout(n_4));
   full_adder__3_157 full_adder_0_5_full_adder_0_i (.a(a[5]), .b(), .cin(n_4), 
      .f(c[5]), .cout(n_5));
   full_adder__3_153 full_adder_0_6_full_adder_0_i (.a(a[6]), .b(), .cin(n_5), 
      .f(c[6]), .cout());
endmodule

module range_extractor__3_201(in_a, in_size, out_a, out_b);
   input [6:0]in_a;
   input [2:0]in_size;
   output [6:0]out_a;
   output [6:0]out_b;

   incrementor__3_200 inc (.a(in_a), .enbl(), .c(out_a));
   int_adder__3_178 add (.a(out_a), .b(in_size), .cin(), .enbl(), .c(out_b), 
      .cout());
endmodule

module half_adder__3_251(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   INV_X1 i_2 (.A(a), .ZN(f));
endmodule

module half_adder__3_248(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_245(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_242(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_239(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_236(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_233(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   XOR2_X1 i_1_0 (.A(a), .B(b), .Z(f));
endmodule

module incrementor__3_252(a, enbl, c);
   input [6:0]a;
   input enbl;
   output [6:0]c;

   half_adder__3_251 half_adder_0_0_half_adder_0_i (.a(a[0]), .b(), .cout(), 
      .f(c[0]));
   half_adder__3_248 half_adder_0_1_half_adder_0_i (.a(a[1]), .b(a[0]), .cout(
      n_0), .f(c[1]));
   half_adder__3_245 half_adder_0_2_half_adder_0_i (.a(a[2]), .b(n_0), .cout(n_1), 
      .f(c[2]));
   half_adder__3_242 half_adder_0_3_half_adder_0_i (.a(a[3]), .b(n_1), .cout(n_2), 
      .f(c[3]));
   half_adder__3_239 half_adder_0_4_half_adder_0_i (.a(a[4]), .b(n_2), .cout(n_3), 
      .f(c[4]));
   half_adder__3_236 half_adder_0_5_half_adder_0_i (.a(a[5]), .b(n_3), .cout(n_4), 
      .f(c[5]));
   half_adder__3_233 half_adder_0_6_half_adder_0_i (.a(a[6]), .b(n_4), .cout(), 
      .f(c[6]));
endmodule

module full_adder__3_229(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(f));
   AND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(cout));
endmodule

module full_adder__3_225(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(f));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(cin), .B1(a), .B2(b), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module full_adder__3_221(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(f));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(cin), .B1(a), .B2(b), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module full_adder__3_217(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__3_213(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__3_209(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__3_205(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
endmodule

module int_adder__3_230(a, b, cin, enbl, c, cout);
   input [6:0]a;
   input [2:0]b;
   input cin;
   input enbl;
   output [6:0]c;
   output cout;

   full_adder__3_229 full_adder_0_0_full_adder_0_i (.a(a[0]), .b(b[0]), .cin(), 
      .f(c[0]), .cout(n_0));
   full_adder__3_225 full_adder_0_1_full_adder_0_i (.a(a[1]), .b(b[1]), .cin(n_0), 
      .f(c[1]), .cout(n_1));
   full_adder__3_221 full_adder_0_2_full_adder_0_i (.a(a[2]), .b(b[2]), .cin(n_1), 
      .f(c[2]), .cout(n_2));
   full_adder__3_217 full_adder_0_3_full_adder_0_i (.a(a[3]), .b(), .cin(n_2), 
      .f(c[3]), .cout(n_3));
   full_adder__3_213 full_adder_0_4_full_adder_0_i (.a(a[4]), .b(), .cin(n_3), 
      .f(c[4]), .cout(n_4));
   full_adder__3_209 full_adder_0_5_full_adder_0_i (.a(a[5]), .b(), .cin(n_4), 
      .f(c[5]), .cout(n_5));
   full_adder__3_205 full_adder_0_6_full_adder_0_i (.a(a[6]), .b(), .cin(n_5), 
      .f(c[6]), .cout());
endmodule

module range_extractor__3_253(in_a, in_size, out_a, out_b);
   input [6:0]in_a;
   input [2:0]in_size;
   output [6:0]out_a;
   output [6:0]out_b;

   incrementor__3_252 inc (.a(in_a), .enbl(), .c(out_a));
   int_adder__3_230 add (.a(out_a), .b(in_size), .cin(), .enbl(), .c(out_b), 
      .cout());
endmodule

module half_adder__3_303(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   INV_X1 i_2 (.A(a), .ZN(f));
endmodule

module half_adder__3_300(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_297(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_294(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_291(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_288(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_285(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   XOR2_X1 i_1_0 (.A(a), .B(b), .Z(f));
endmodule

module incrementor__3_304(a, enbl, c);
   input [6:0]a;
   input enbl;
   output [6:0]c;

   half_adder__3_303 half_adder_0_0_half_adder_0_i (.a(a[0]), .b(), .cout(), 
      .f(c[0]));
   half_adder__3_300 half_adder_0_1_half_adder_0_i (.a(a[1]), .b(a[0]), .cout(
      n_0), .f(c[1]));
   half_adder__3_297 half_adder_0_2_half_adder_0_i (.a(a[2]), .b(n_0), .cout(n_1), 
      .f(c[2]));
   half_adder__3_294 half_adder_0_3_half_adder_0_i (.a(a[3]), .b(n_1), .cout(n_2), 
      .f(c[3]));
   half_adder__3_291 half_adder_0_4_half_adder_0_i (.a(a[4]), .b(n_2), .cout(n_3), 
      .f(c[4]));
   half_adder__3_288 half_adder_0_5_half_adder_0_i (.a(a[5]), .b(n_3), .cout(n_4), 
      .f(c[5]));
   half_adder__3_285 half_adder_0_6_half_adder_0_i (.a(a[6]), .b(n_4), .cout(), 
      .f(c[6]));
endmodule

module full_adder__3_281(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(f));
   AND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(cout));
endmodule

module full_adder__3_277(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(f));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(cin), .B1(a), .B2(b), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module full_adder__3_273(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(f));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(cin), .B1(a), .B2(b), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module full_adder__3_269(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__3_265(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__3_261(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__3_257(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
endmodule

module int_adder__3_282(a, b, cin, enbl, c, cout);
   input [6:0]a;
   input [2:0]b;
   input cin;
   input enbl;
   output [6:0]c;
   output cout;

   full_adder__3_281 full_adder_0_0_full_adder_0_i (.a(a[0]), .b(b[0]), .cin(), 
      .f(c[0]), .cout(n_0));
   full_adder__3_277 full_adder_0_1_full_adder_0_i (.a(a[1]), .b(b[1]), .cin(n_0), 
      .f(c[1]), .cout(n_1));
   full_adder__3_273 full_adder_0_2_full_adder_0_i (.a(a[2]), .b(b[2]), .cin(n_1), 
      .f(c[2]), .cout(n_2));
   full_adder__3_269 full_adder_0_3_full_adder_0_i (.a(a[3]), .b(), .cin(n_2), 
      .f(c[3]), .cout(n_3));
   full_adder__3_265 full_adder_0_4_full_adder_0_i (.a(a[4]), .b(), .cin(n_3), 
      .f(c[4]), .cout(n_4));
   full_adder__3_261 full_adder_0_5_full_adder_0_i (.a(a[5]), .b(), .cin(n_4), 
      .f(c[5]), .cout(n_5));
   full_adder__3_257 full_adder_0_6_full_adder_0_i (.a(a[6]), .b(), .cin(n_5), 
      .f(c[6]), .cout());
endmodule

module range_extractor__3_305(in_a, in_size, out_a, out_b);
   input [6:0]in_a;
   input [2:0]in_size;
   output [6:0]out_a;
   output [6:0]out_b;

   incrementor__3_304 inc (.a(in_a), .enbl(), .c(out_a));
   int_adder__3_282 add (.a(out_a), .b(in_size), .cin(), .enbl(), .c(out_b), 
      .cout());
endmodule

module half_adder__3_355(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   INV_X1 i_2 (.A(a), .ZN(f));
endmodule

module half_adder__3_352(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_349(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_346(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_343(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_340(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_337(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   XOR2_X1 i_1_0 (.A(a), .B(b), .Z(f));
endmodule

module incrementor__3_356(a, enbl, c);
   input [6:0]a;
   input enbl;
   output [6:0]c;

   half_adder__3_355 half_adder_0_0_half_adder_0_i (.a(a[0]), .b(), .cout(), 
      .f(c[0]));
   half_adder__3_352 half_adder_0_1_half_adder_0_i (.a(a[1]), .b(a[0]), .cout(
      n_0), .f(c[1]));
   half_adder__3_349 half_adder_0_2_half_adder_0_i (.a(a[2]), .b(n_0), .cout(n_1), 
      .f(c[2]));
   half_adder__3_346 half_adder_0_3_half_adder_0_i (.a(a[3]), .b(n_1), .cout(n_2), 
      .f(c[3]));
   half_adder__3_343 half_adder_0_4_half_adder_0_i (.a(a[4]), .b(n_2), .cout(n_3), 
      .f(c[4]));
   half_adder__3_340 half_adder_0_5_half_adder_0_i (.a(a[5]), .b(n_3), .cout(n_4), 
      .f(c[5]));
   half_adder__3_337 half_adder_0_6_half_adder_0_i (.a(a[6]), .b(n_4), .cout(), 
      .f(c[6]));
endmodule

module full_adder__3_333(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(f));
   AND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(cout));
endmodule

module full_adder__3_329(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(f));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(cin), .B1(a), .B2(b), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module full_adder__3_325(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(f));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(cin), .B1(a), .B2(b), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module full_adder__3_321(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__3_317(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__3_313(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__3_309(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
endmodule

module int_adder__3_334(a, b, cin, enbl, c, cout);
   input [6:0]a;
   input [2:0]b;
   input cin;
   input enbl;
   output [6:0]c;
   output cout;

   full_adder__3_333 full_adder_0_0_full_adder_0_i (.a(a[0]), .b(b[0]), .cin(), 
      .f(c[0]), .cout(n_0));
   full_adder__3_329 full_adder_0_1_full_adder_0_i (.a(a[1]), .b(b[1]), .cin(n_0), 
      .f(c[1]), .cout(n_1));
   full_adder__3_325 full_adder_0_2_full_adder_0_i (.a(a[2]), .b(b[2]), .cin(n_1), 
      .f(c[2]), .cout(n_2));
   full_adder__3_321 full_adder_0_3_full_adder_0_i (.a(a[3]), .b(), .cin(n_2), 
      .f(c[3]), .cout(n_3));
   full_adder__3_317 full_adder_0_4_full_adder_0_i (.a(a[4]), .b(), .cin(n_3), 
      .f(c[4]), .cout(n_4));
   full_adder__3_313 full_adder_0_5_full_adder_0_i (.a(a[5]), .b(), .cin(n_4), 
      .f(c[5]), .cout(n_5));
   full_adder__3_309 full_adder_0_6_full_adder_0_i (.a(a[6]), .b(), .cin(n_5), 
      .f(c[6]), .cout());
endmodule

module range_extractor__3_357(in_a, in_size, out_a, out_b);
   input [6:0]in_a;
   input [2:0]in_size;
   output [6:0]out_a;
   output [6:0]out_b;

   incrementor__3_356 inc (.a(in_a), .enbl(), .c(out_a));
   int_adder__3_334 add (.a(out_a), .b(in_size), .cin(), .enbl(), .c(out_b), 
      .cout());
endmodule

module half_adder__3_407(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   INV_X1 i_2 (.A(a), .ZN(f));
endmodule

module half_adder__3_404(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_401(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_398(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_395(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_392(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_389(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   XOR2_X1 i_1_0 (.A(a), .B(b), .Z(f));
endmodule

module incrementor__3_408(a, enbl, c);
   input [6:0]a;
   input enbl;
   output [6:0]c;

   half_adder__3_407 half_adder_0_0_half_adder_0_i (.a(a[0]), .b(), .cout(), 
      .f(c[0]));
   half_adder__3_404 half_adder_0_1_half_adder_0_i (.a(a[1]), .b(a[0]), .cout(
      n_0), .f(c[1]));
   half_adder__3_401 half_adder_0_2_half_adder_0_i (.a(a[2]), .b(n_0), .cout(n_1), 
      .f(c[2]));
   half_adder__3_398 half_adder_0_3_half_adder_0_i (.a(a[3]), .b(n_1), .cout(n_2), 
      .f(c[3]));
   half_adder__3_395 half_adder_0_4_half_adder_0_i (.a(a[4]), .b(n_2), .cout(n_3), 
      .f(c[4]));
   half_adder__3_392 half_adder_0_5_half_adder_0_i (.a(a[5]), .b(n_3), .cout(n_4), 
      .f(c[5]));
   half_adder__3_389 half_adder_0_6_half_adder_0_i (.a(a[6]), .b(n_4), .cout(), 
      .f(c[6]));
endmodule

module full_adder__3_385(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(f));
   AND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(cout));
endmodule

module full_adder__3_381(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(f));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(cin), .B1(a), .B2(b), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module full_adder__3_377(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(f));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(cin), .B1(a), .B2(b), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module full_adder__3_373(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__3_369(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__3_365(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__3_361(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
endmodule

module int_adder__3_386(a, b, cin, enbl, c, cout);
   input [6:0]a;
   input [2:0]b;
   input cin;
   input enbl;
   output [6:0]c;
   output cout;

   full_adder__3_385 full_adder_0_0_full_adder_0_i (.a(a[0]), .b(b[0]), .cin(), 
      .f(c[0]), .cout(n_0));
   full_adder__3_381 full_adder_0_1_full_adder_0_i (.a(a[1]), .b(b[1]), .cin(n_0), 
      .f(c[1]), .cout(n_1));
   full_adder__3_377 full_adder_0_2_full_adder_0_i (.a(a[2]), .b(b[2]), .cin(n_1), 
      .f(c[2]), .cout(n_2));
   full_adder__3_373 full_adder_0_3_full_adder_0_i (.a(a[3]), .b(), .cin(n_2), 
      .f(c[3]), .cout(n_3));
   full_adder__3_369 full_adder_0_4_full_adder_0_i (.a(a[4]), .b(), .cin(n_3), 
      .f(c[4]), .cout(n_4));
   full_adder__3_365 full_adder_0_5_full_adder_0_i (.a(a[5]), .b(), .cin(n_4), 
      .f(c[5]), .cout(n_5));
   full_adder__3_361 full_adder_0_6_full_adder_0_i (.a(a[6]), .b(), .cin(n_5), 
      .f(c[6]), .cout());
endmodule

module range_extractor__3_409(in_a, in_size, out_a, out_b);
   input [6:0]in_a;
   input [2:0]in_size;
   output [6:0]out_a;
   output [6:0]out_b;

   incrementor__3_408 inc (.a(in_a), .enbl(), .c(out_a));
   int_adder__3_386 add (.a(out_a), .b(in_size), .cin(), .enbl(), .c(out_b), 
      .cout());
endmodule

module half_adder__3_459(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   INV_X1 i_2 (.A(a), .ZN(f));
endmodule

module half_adder__3_456(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_453(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_450(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_447(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_444(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_441(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   XOR2_X1 i_1_0 (.A(a), .B(b), .Z(f));
endmodule

module incrementor__3_460(a, enbl, c);
   input [6:0]a;
   input enbl;
   output [6:0]c;

   half_adder__3_459 half_adder_0_0_half_adder_0_i (.a(a[0]), .b(), .cout(), 
      .f(c[0]));
   half_adder__3_456 half_adder_0_1_half_adder_0_i (.a(a[1]), .b(a[0]), .cout(
      n_0), .f(c[1]));
   half_adder__3_453 half_adder_0_2_half_adder_0_i (.a(a[2]), .b(n_0), .cout(n_1), 
      .f(c[2]));
   half_adder__3_450 half_adder_0_3_half_adder_0_i (.a(a[3]), .b(n_1), .cout(n_2), 
      .f(c[3]));
   half_adder__3_447 half_adder_0_4_half_adder_0_i (.a(a[4]), .b(n_2), .cout(n_3), 
      .f(c[4]));
   half_adder__3_444 half_adder_0_5_half_adder_0_i (.a(a[5]), .b(n_3), .cout(n_4), 
      .f(c[5]));
   half_adder__3_441 half_adder_0_6_half_adder_0_i (.a(a[6]), .b(n_4), .cout(), 
      .f(c[6]));
endmodule

module full_adder__3_437(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(f));
   AND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(cout));
endmodule

module full_adder__3_433(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(f));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(cin), .B1(a), .B2(b), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module full_adder__3_429(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(f));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(cin), .B1(a), .B2(b), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module full_adder__3_425(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__3_421(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__3_417(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__3_413(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
endmodule

module int_adder__3_438(a, b, cin, enbl, c, cout);
   input [6:0]a;
   input [2:0]b;
   input cin;
   input enbl;
   output [6:0]c;
   output cout;

   full_adder__3_437 full_adder_0_0_full_adder_0_i (.a(a[0]), .b(b[0]), .cin(), 
      .f(c[0]), .cout(n_0));
   full_adder__3_433 full_adder_0_1_full_adder_0_i (.a(a[1]), .b(b[1]), .cin(n_0), 
      .f(c[1]), .cout(n_1));
   full_adder__3_429 full_adder_0_2_full_adder_0_i (.a(a[2]), .b(b[2]), .cin(n_1), 
      .f(c[2]), .cout(n_2));
   full_adder__3_425 full_adder_0_3_full_adder_0_i (.a(a[3]), .b(), .cin(n_2), 
      .f(c[3]), .cout(n_3));
   full_adder__3_421 full_adder_0_4_full_adder_0_i (.a(a[4]), .b(), .cin(n_3), 
      .f(c[4]), .cout(n_4));
   full_adder__3_417 full_adder_0_5_full_adder_0_i (.a(a[5]), .b(), .cin(n_4), 
      .f(c[5]), .cout(n_5));
   full_adder__3_413 full_adder_0_6_full_adder_0_i (.a(a[6]), .b(), .cin(n_5), 
      .f(c[6]), .cout());
endmodule

module range_extractor__3_461(in_a, in_size, out_a, out_b);
   input [6:0]in_a;
   input [2:0]in_size;
   output [6:0]out_a;
   output [6:0]out_b;

   incrementor__3_460 inc (.a(in_a), .enbl(), .c(out_a));
   int_adder__3_438 add (.a(out_a), .b(in_size), .cin(), .enbl(), .c(out_b), 
      .cout());
endmodule

module half_adder__3_82(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   INV_X1 i_2 (.A(a), .ZN(f));
endmodule

module half_adder__3_85(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_88(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_91(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_94(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder__3_97(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   AND2_X1 i_0_0 (.A1(a), .A2(b), .ZN(cout));
   XOR2_X1 i_0_1 (.A(a), .B(b), .Z(f));
endmodule

module half_adder(a, b, cout, f);
   input a;
   input b;
   output cout;
   output f;

   XOR2_X1 i_1_0 (.A(a), .B(b), .Z(f));
endmodule

module incrementor(a, enbl, c);
   input [6:0]a;
   input enbl;
   output [6:0]c;

   half_adder__3_82 half_adder_0_0_half_adder_0_i (.a(a[0]), .b(), .cout(), 
      .f(c[0]));
   half_adder__3_85 half_adder_0_1_half_adder_0_i (.a(a[1]), .b(a[0]), .cout(n_0), 
      .f(c[1]));
   half_adder__3_88 half_adder_0_2_half_adder_0_i (.a(a[2]), .b(n_0), .cout(n_1), 
      .f(c[2]));
   half_adder__3_91 half_adder_0_3_half_adder_0_i (.a(a[3]), .b(n_1), .cout(n_2), 
      .f(c[3]));
   half_adder__3_94 half_adder_0_4_half_adder_0_i (.a(a[4]), .b(n_2), .cout(n_3), 
      .f(c[4]));
   half_adder__3_97 half_adder_0_5_half_adder_0_i (.a(a[5]), .b(n_3), .cout(n_4), 
      .f(c[5]));
   half_adder half_adder_0_6_half_adder_0_i (.a(a[6]), .b(n_4), .cout(), 
      .f(c[6]));
endmodule

module full_adder__3_3(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(f));
   AND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(cout));
endmodule

module full_adder__3_7(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(f));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(cin), .B1(a), .B2(b), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module full_adder__3_11(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(f));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(cin), .B1(a), .B2(b), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module full_adder__3_15(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__3_19(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__3_23(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__3_27(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
endmodule

module int_adder(a, b, cin, enbl, c, cout);
   input [6:0]a;
   input [2:0]b;
   input cin;
   input enbl;
   output [6:0]c;
   output cout;

   full_adder__3_3 full_adder_0_0_full_adder_0_i (.a(a[0]), .b(b[0]), .cin(), 
      .f(c[0]), .cout(n_0));
   full_adder__3_7 full_adder_0_1_full_adder_0_i (.a(a[1]), .b(b[1]), .cin(n_0), 
      .f(c[1]), .cout(n_1));
   full_adder__3_11 full_adder_0_2_full_adder_0_i (.a(a[2]), .b(b[2]), .cin(n_1), 
      .f(c[2]), .cout(n_2));
   full_adder__3_15 full_adder_0_3_full_adder_0_i (.a(a[3]), .b(), .cin(n_2), 
      .f(c[3]), .cout(n_3));
   full_adder__3_19 full_adder_0_4_full_adder_0_i (.a(a[4]), .b(), .cin(n_3), 
      .f(c[4]), .cout(n_4));
   full_adder__3_23 full_adder_0_5_full_adder_0_i (.a(a[5]), .b(), .cin(n_4), 
      .f(c[5]), .cout(n_5));
   full_adder__3_27 full_adder_0_6_full_adder_0_i (.a(a[6]), .b(), .cin(n_5), 
      .f(c[6]), .cout());
endmodule

module range_extractor(in_a, in_size, out_a, out_b);
   input [6:0]in_a;
   input [2:0]in_size;
   output [6:0]out_a;
   output [6:0]out_b;

   incrementor inc (.a(in_a), .enbl(), .c(out_a));
   int_adder add (.a(out_a), .b(in_size), .cin(), .enbl(), .c(out_b), .cout());
endmodule

module decompressor(in_data, rst, enbl_in, clk, state_wait, out_ready, out_data, 
      error_success, buf_test);
   input [31:0]in_data;
   input rst;
   input enbl_in;
   input clk;
   input state_wait;
   output out_ready;
   output [31:0]out_data;
   output error_success;
   output [127:0]buf_test;

   wire n_8_0_5;
   wire n_8_0_4;
   wire n_8_0_0;
   wire n_8_0_3;
   wire n_8_0_1;
   wire n_8_0_2;
   wire n_8_0_6;
   wire n_8_0_7;
   wire n_8_0_8;
   wire n_8_0_9;
   wire n_8_0_10;
   wire n_8_0_11;
   wire n_8_0_12;
   wire n_8_0_13;
   wire n_8_0_14;
   wire n_8_0_15;
   wire n_8_0_16;
   wire n_8_0_17;
   wire n_8_0_18;
   wire n_8_0_19;
   wire n_8_0_20;
   wire n_8_0_21;
   wire n_8_0_22;
   wire n_8_0_23;
   wire n_8_0_24;
   wire n_8_0_25;
   wire n_8_0_26;
   wire n_8_0_27;
   wire n_8_0_28;
   wire n_8_0_29;
   wire n_8_0_30;
   wire n_8_0_31;
   wire n_8_0_32;
   wire n_8_0_33;
   wire n_8_0_34;
   wire n_8_0_35;
   wire n_8_0_36;
   wire n_8_0_37;
   wire n_8_0_38;
   wire n_8_0_39;
   wire n_8_0_40;
   wire n_8_0_41;
   wire n_8_0_42;
   wire n_8_0_43;
   wire n_8_0_44;
   wire n_8_0_45;
   wire n_8_0_46;
   wire n_8_0_47;
   wire n_8_0_48;
   wire n_8_0_49;
   wire n_8_0_50;
   wire n_8_0_51;
   wire n_8_0_52;
   wire n_8_0_53;
   wire n_8_0_54;
   wire n_8_0_55;
   wire n_8_0_56;
   wire n_8_0_57;
   wire n_8_0_58;
   wire n_8_0_59;
   wire n_8_0_60;
   wire n_8_0_61;
   wire n_8_0_62;
   wire n_8_0_63;
   wire n_8_0_64;
   wire n_8_0_65;
   wire n_8_0_66;
   wire n_8_0_67;
   wire n_8_0_68;
   wire n_8_0_69;
   wire n_8_0_70;
   wire n_8_0_71;
   wire n_8_0_72;
   wire n_8_0_73;
   wire n_8_0_74;
   wire n_8_0_75;
   wire n_8_0_76;
   wire n_8_0_77;
   wire n_8_0_78;
   wire n_8_0_79;
   wire n_8_0_80;
   wire n_8_0_81;
   wire n_8_0_82;
   wire n_8_0_83;
   wire n_8_0_84;
   wire n_8_0_85;
   wire n_8_0_86;
   wire n_8_0_87;
   wire n_8_0_88;
   wire n_8_0_89;
   wire n_8_0_90;
   wire n_8_0_91;
   wire n_8_0_92;
   wire n_8_0_93;
   wire n_8_0_94;
   wire n_8_0_95;
   wire n_8_0_96;
   wire n_8_0_97;
   wire n_8_0_98;
   wire n_8_0_99;
   wire n_8_0_100;
   wire n_8_0_101;
   wire n_8_0_102;
   wire n_8_0_103;
   wire n_8_0_104;
   wire n_8_0_105;
   wire n_8_0_106;
   wire n_8_0_107;
   wire n_8_0_108;
   wire n_8_0_109;
   wire n_8_0_110;
   wire n_8_0_111;
   wire n_8_0_112;
   wire n_8_0_113;
   wire n_8_0_114;
   wire n_8_0_115;
   wire n_8_0_116;
   wire n_8_0_117;
   wire n_8_0_118;
   wire n_8_0_119;
   wire n_8_0_120;
   wire n_8_0_121;
   wire n_8_0_122;
   wire n_8_0_123;
   wire n_8_0_124;
   wire n_8_0_125;
   wire n_8_0_126;
   wire n_8_0_127;
   wire n_8_0_128;
   wire n_8_0_129;
   wire n_8_0_130;
   wire n_8_0_131;
   wire n_8_0_132;
   wire n_8_0_133;
   wire n_8_0_134;
   wire n_8_0_135;
   wire n_8_0_136;
   wire n_8_0_137;
   wire n_8_0_138;
   wire n_8_0_139;
   wire n_8_0_140;
   wire n_8_0_141;
   wire n_8_0_142;
   wire n_8_0_143;
   wire n_8_0_144;
   wire n_8_0_145;
   wire n_8_0_146;
   wire n_8_0_147;
   wire n_8_0_148;
   wire n_8_0_149;
   wire n_8_0_150;
   wire n_8_0_151;
   wire n_8_0_152;
   wire n_8_0_153;
   wire n_8_0_154;
   wire n_8_0_155;
   wire n_8_0_156;
   wire n_8_0_157;
   wire n_8_0_158;
   wire n_8_0_159;
   wire n_8_0_160;
   wire n_8_0_161;
   wire n_8_0_162;
   wire n_8_0_163;
   wire n_8_0_164;
   wire n_8_0_165;
   wire n_8_0_166;
   wire n_8_0_167;
   wire n_8_0_168;
   wire n_8_0_169;
   wire n_8_0_170;
   wire n_8_0_171;
   wire n_8_0_172;
   wire n_8_0_173;
   wire n_8_0_174;
   wire n_8_0_175;
   wire n_8_0_176;
   wire n_8_0_177;
   wire n_8_0_178;
   wire n_8_0_179;
   wire n_8_0_180;
   wire n_8_0_181;
   wire n_8_0_182;
   wire n_8_0_183;
   wire n_8_0_184;
   wire n_8_0_185;
   wire n_8_0_186;
   wire n_8_0_187;
   wire n_8_0_188;
   wire n_8_0_189;
   wire n_8_0_190;
   wire n_8_0_191;
   wire n_8_0_192;
   wire n_8_0_193;
   wire n_8_0_194;
   wire n_8_0_195;
   wire n_8_0_196;
   wire n_8_0_197;
   wire n_8_0_198;
   wire n_8_0_199;
   wire n_8_0_200;
   wire n_8_0_201;
   wire n_8_0_202;
   wire n_8_0_203;
   wire n_8_0_204;
   wire n_8_0_205;
   wire n_8_0_206;
   wire n_8_0_207;
   wire n_8_0_208;
   wire n_8_0_209;
   wire n_8_0_210;
   wire n_8_0_211;
   wire n_8_0_212;
   wire n_8_0_213;
   wire n_8_0_214;
   wire n_8_0_215;
   wire n_8_0_216;
   wire n_8_0_217;
   wire n_8_0_218;
   wire n_8_0_219;
   wire n_8_0_220;
   wire n_8_0_221;
   wire n_8_0_222;
   wire n_8_0_223;
   wire n_8_0_224;
   wire n_8_0_225;
   wire n_8_0_226;
   wire n_8_0_227;
   wire n_8_0_228;
   wire n_8_0_229;
   wire n_8_0_230;
   wire n_8_0_231;
   wire n_8_0_232;
   wire n_8_0_233;
   wire n_8_0_234;
   wire n_8_0_235;
   wire n_8_0_236;
   wire n_8_0_237;
   wire n_8_0_238;
   wire n_8_0_239;
   wire n_8_0_240;
   wire n_8_0_241;
   wire n_8_0_242;
   wire n_8_0_243;
   wire n_8_0_244;
   wire n_8_0_245;
   wire n_8_0_246;
   wire n_8_0_247;
   wire n_8_0_248;
   wire n_8_0_249;
   wire n_8_0_250;
   wire n_8_0_251;
   wire n_8_0_252;
   wire n_8_0_253;
   wire n_8_0_254;
   wire n_8_0_255;
   wire n_8_0_256;
   wire n_8_0_257;
   wire n_8_0_258;
   wire n_8_0_259;
   wire n_8_0_260;
   wire n_8_0_261;
   wire n_8_0_262;
   wire n_8_0_263;
   wire n_8_0_264;
   wire n_8_0_265;
   wire n_8_0_266;
   wire n_8_0_267;
   wire n_8_0_268;
   wire n_8_0_269;
   wire n_8_0_270;
   wire n_8_0_271;
   wire n_8_0_272;
   wire n_8_0_273;
   wire n_8_0_274;
   wire n_8_0_275;
   wire n_8_0_276;
   wire n_8_0_277;
   wire n_8_0_278;
   wire n_8_0_279;
   wire n_8_0_280;
   wire n_8_0_281;
   wire n_8_0_282;
   wire n_8_0_283;
   wire n_8_0_284;
   wire n_8_0_285;
   wire n_8_0_286;
   wire n_8_0_287;
   wire n_8_0_288;
   wire n_8_0_289;
   wire n_8_0_290;
   wire n_8_0_291;
   wire n_8_0_292;
   wire n_8_0_293;
   wire n_8_0_294;
   wire n_8_0_295;
   wire n_8_0_296;
   wire n_8_0_297;
   wire n_8_0_298;
   wire n_8_0_299;
   wire n_8_0_300;
   wire n_8_0_301;
   wire n_8_0_302;
   wire n_8_0_303;
   wire n_8_0_304;
   wire n_8_0_305;
   wire n_8_0_306;
   wire n_8_0_307;
   wire n_8_0_308;
   wire n_8_0_309;
   wire n_8_0_310;
   wire n_8_0_311;
   wire n_8_0_312;
   wire n_8_0_313;
   wire n_8_0_314;
   wire n_8_0_315;
   wire n_8_0_316;
   wire n_8_0_317;
   wire n_8_0_318;
   wire n_8_0_319;
   wire n_8_0_320;
   wire n_8_0_321;
   wire n_8_0_322;
   wire n_8_0_323;
   wire n_8_0_324;
   wire n_8_0_325;
   wire n_8_0_326;
   wire n_8_0_327;
   wire n_8_0_328;
   wire n_8_0_329;
   wire n_8_0_330;
   wire n_8_0_331;
   wire n_8_0_332;
   wire n_8_0_333;
   wire n_8_0_334;
   wire n_8_0_335;
   wire n_8_0_336;
   wire n_8_0_337;
   wire n_8_0_338;
   wire n_8_0_339;
   wire n_8_0_340;
   wire n_8_0_341;
   wire n_8_0_342;
   wire n_8_0_343;
   wire n_8_0_344;
   wire n_8_0_345;
   wire n_8_0_346;
   wire n_8_0_347;
   wire n_8_0_348;
   wire n_8_0_349;
   wire n_8_0_350;
   wire n_8_0_351;
   wire n_8_0_352;
   wire n_8_0_353;
   wire n_8_0_354;
   wire n_8_0_355;
   wire n_8_0_356;
   wire n_8_0_357;
   wire n_8_0_358;
   wire n_8_0_359;
   wire n_8_0_360;
   wire n_8_0_361;
   wire n_8_0_362;
   wire n_8_0_363;
   wire n_8_0_364;
   wire n_8_0_365;
   wire n_8_0_366;
   wire n_8_0_367;
   wire n_8_0_368;
   wire n_8_0_369;
   wire n_8_0_370;
   wire n_8_0_371;
   wire n_8_0_372;
   wire n_8_0_373;
   wire n_8_0_374;
   wire n_8_0_375;
   wire n_8_0_376;
   wire n_8_0_377;
   wire n_8_0_378;
   wire n_8_0_379;
   wire n_8_0_380;
   wire n_8_0_381;
   wire n_8_0_382;
   wire n_8_0_383;
   wire n_8_0_384;
   wire n_8_0_385;
   wire n_8_0_386;
   wire n_8_0_387;
   wire n_8_0_388;
   wire n_8_0_389;
   wire n_8_0_390;
   wire n_8_0_391;
   wire n_8_0_392;
   wire n_8_0_393;
   wire n_8_0_394;
   wire n_8_0_395;
   wire n_8_0_396;
   wire n_8_0_397;
   wire n_8_0_398;
   wire n_8_0_399;
   wire n_8_0_400;
   wire n_8_0_401;
   wire n_8_0_402;
   wire n_8_0_403;
   wire n_8_0_404;
   wire n_8_0_405;
   wire n_8_0_406;
   wire n_8_0_407;
   wire n_8_0_408;
   wire n_8_0_409;
   wire n_8_0_410;
   wire n_8_0_411;
   wire n_8_0_412;
   wire n_8_0_413;
   wire n_8_0_414;
   wire n_8_0_415;
   wire n_8_0_416;
   wire n_8_0_417;
   wire n_8_0_418;
   wire n_8_0_419;
   wire n_8_0_420;
   wire n_8_0_421;
   wire n_8_0_422;
   wire n_8_0_423;
   wire n_8_0_424;
   wire n_8_0_425;
   wire n_8_0_426;
   wire n_8_0_427;
   wire n_8_0_428;
   wire n_8_0_429;
   wire n_8_0_430;
   wire n_8_0_431;
   wire n_8_0_432;
   wire n_8_0_433;
   wire n_8_0_434;
   wire n_8_0_435;
   wire n_8_0_436;
   wire n_8_0_437;
   wire n_8_0_438;
   wire n_8_0_439;
   wire n_8_0_440;
   wire n_8_0_441;
   wire n_8_0_442;
   wire n_8_0_443;
   wire n_8_0_444;
   wire n_8_0_445;
   wire n_8_0_446;
   wire n_8_0_447;
   wire n_8_0_448;
   wire n_8_0_449;
   wire n_8_0_450;
   wire n_8_0_451;
   wire n_8_0_452;
   wire n_8_0_453;
   wire n_8_0_454;
   wire n_8_0_455;
   wire n_8_0_456;
   wire n_8_0_457;
   wire n_8_0_458;
   wire n_8_0_459;
   wire n_8_0_460;
   wire n_8_0_461;
   wire n_8_0_462;
   wire n_8_0_463;
   wire n_8_0_464;
   wire n_8_0_465;
   wire n_8_0_466;
   wire n_8_0_467;
   wire n_8_0_468;
   wire n_8_0_469;
   wire n_8_0_470;
   wire n_8_0_471;
   wire n_8_0_472;
   wire n_8_0_473;
   wire n_8_0_474;
   wire n_8_0_475;
   wire n_8_0_476;
   wire n_8_0_477;
   wire n_8_0_478;
   wire n_8_0_479;
   wire n_8_0_480;
   wire n_8_0_481;
   wire n_8_0_482;
   wire n_8_0_483;
   wire n_8_0_484;
   wire n_8_0_485;
   wire n_8_0_486;
   wire n_8_0_487;
   wire n_8_0_488;
   wire n_8_0_489;
   wire n_8_0_490;
   wire n_8_0_491;
   wire n_8_0_492;
   wire n_8_0_493;
   wire n_8_0_494;
   wire n_8_0_495;
   wire n_8_0_496;
   wire n_8_0_497;
   wire n_8_0_498;
   wire n_8_0_499;
   wire n_8_0_500;
   wire n_8_0_501;
   wire n_8_0_502;
   wire n_8_0_503;
   wire n_8_0_504;
   wire n_8_0_505;
   wire n_8_0_506;
   wire n_8_0_507;
   wire n_8_0_508;
   wire n_8_0_509;
   wire n_8_0_510;
   wire n_8_0_511;
   wire n_8_0_512;
   wire n_8_0_513;
   wire n_8_0_514;
   wire n_8_0_515;
   wire n_8_0_516;
   wire n_8_0_517;
   wire n_8_0_518;
   wire n_8_0_519;
   wire n_8_0_520;
   wire n_8_0_521;
   wire n_8_0_522;
   wire n_8_0_523;
   wire n_8_0_524;
   wire n_8_0_525;
   wire n_8_0_526;
   wire n_8_0_527;
   wire n_8_0_528;
   wire n_8_0_529;
   wire n_8_0_530;
   wire n_8_0_531;
   wire n_8_0_532;
   wire n_8_0_533;
   wire n_8_0_534;
   wire n_8_0_535;
   wire n_8_0_536;
   wire n_8_0_537;
   wire n_8_0_538;
   wire n_8_0_539;
   wire n_8_0_540;
   wire n_8_0_541;
   wire n_8_0_542;
   wire n_8_0_543;
   wire n_8_0_544;
   wire n_8_0_545;
   wire n_8_0_546;
   wire n_8_0_547;
   wire n_8_0_548;
   wire n_8_0_549;
   wire n_8_0_550;
   wire n_8_0_551;
   wire n_8_0_552;
   wire n_8_0_553;
   wire n_8_0_554;
   wire n_8_0_555;
   wire n_8_0_556;
   wire n_8_0_557;
   wire n_8_0_558;
   wire n_8_0_559;
   wire n_8_0_560;
   wire n_8_0_561;
   wire n_8_0_562;
   wire n_8_0_563;
   wire n_8_0_564;
   wire n_8_0_565;
   wire n_8_0_566;
   wire n_8_0_567;
   wire n_8_0_568;
   wire n_8_0_569;
   wire n_8_0_570;
   wire n_8_0_571;
   wire n_8_0_572;
   wire n_8_0_573;
   wire n_8_0_574;
   wire n_8_0_575;
   wire n_8_0_576;
   wire n_8_0_577;
   wire n_8_0_578;
   wire n_8_0_579;
   wire n_8_0_580;
   wire n_8_0_581;
   wire n_8_0_582;
   wire n_8_0_583;
   wire n_8_0_584;
   wire n_8_0_585;
   wire n_8_0_586;
   wire n_8_0_587;
   wire n_8_0_588;
   wire n_8_0_589;
   wire n_8_0_590;
   wire n_8_0_591;
   wire n_8_0_592;
   wire n_8_0_593;
   wire n_8_0_594;
   wire n_8_0_595;
   wire n_8_0_596;
   wire n_8_0_597;
   wire n_8_0_598;
   wire n_8_0_599;
   wire n_8_0_600;
   wire n_8_0_601;
   wire n_8_0_602;
   wire n_8_0_603;
   wire n_8_0_604;
   wire n_8_0_605;
   wire n_8_0_606;
   wire n_8_0_607;
   wire n_8_0_608;
   wire n_8_0_609;
   wire n_8_0_610;
   wire n_8_0_611;
   wire n_8_0_612;
   wire n_8_0_613;
   wire n_8_0_614;
   wire n_8_0_615;
   wire n_8_0_616;
   wire n_8_0_617;
   wire n_8_0_618;
   wire n_8_0_619;
   wire n_8_0_620;
   wire n_8_0_621;
   wire n_8_0_622;
   wire n_8_0_623;
   wire n_8_0_624;
   wire n_8_0_625;
   wire n_8_0_626;
   wire n_8_0_627;
   wire n_8_0_628;
   wire n_8_0_629;
   wire n_8_0_630;
   wire n_8_0_631;
   wire n_8_0_632;
   wire n_8_0_633;
   wire n_8_0_634;
   wire n_8_0_635;
   wire n_8_0_636;
   wire n_8_0_637;
   wire n_8_0_638;
   wire n_8_0_639;
   wire n_8_0_640;
   wire n_8_0_641;
   wire n_8_0_642;
   wire n_8_0_643;
   wire n_8_0_644;
   wire n_8_0_645;
   wire n_8_0_646;
   wire n_8_0_647;
   wire n_8_0_648;
   wire n_8_0_649;
   wire n_8_0_650;
   wire n_8_0_651;
   wire n_8_0_652;
   wire n_8_0_653;
   wire n_8_0_654;
   wire n_8_0_655;
   wire n_8_0_656;
   wire n_8_0_657;
   wire n_8_0_658;
   wire n_8_0_659;
   wire n_8_0_660;
   wire n_8_0_661;
   wire n_8_0_662;
   wire n_8_0_663;
   wire n_8_0_664;
   wire n_8_0_665;
   wire n_8_0_666;
   wire n_8_0_667;
   wire n_8_0_668;
   wire n_8_0_669;
   wire n_8_0_670;
   wire n_8_0_671;
   wire n_8_0_672;
   wire n_8_0_673;
   wire n_8_0_674;
   wire n_8_0_675;
   wire n_8_0_676;
   wire n_8_0_677;
   wire n_8_0_678;
   wire n_8_0_679;
   wire n_8_0_680;
   wire n_8_0_681;
   wire n_8_0_682;
   wire n_8_0_683;
   wire n_8_0_684;
   wire n_8_0_685;
   wire n_8_0_686;
   wire n_8_0_687;
   wire n_8_0_688;
   wire n_8_0_689;
   wire n_8_0_690;
   wire n_8_0_691;
   wire n_8_0_692;
   wire n_8_0_693;
   wire n_8_0_694;
   wire n_8_0_695;
   wire n_8_0_696;
   wire n_8_0_697;
   wire n_8_0_698;
   wire n_8_0_699;
   wire n_8_0_700;
   wire n_8_0_701;
   wire n_8_0_702;
   wire n_8_0_703;
   wire n_8_0_704;
   wire n_8_0_705;
   wire n_8_0_706;
   wire n_8_0_707;
   wire n_8_0_708;
   wire n_8_0_709;
   wire n_8_0_710;
   wire n_8_0_711;
   wire n_8_0_712;
   wire n_8_0_713;
   wire n_8_0_714;
   wire n_8_0_715;
   wire n_8_0_716;
   wire n_8_0_717;
   wire n_8_0_718;
   wire n_8_0_719;
   wire n_8_0_720;
   wire n_8_0_721;
   wire n_8_0_722;
   wire n_8_0_723;
   wire n_8_0_724;
   wire n_8_0_725;
   wire n_8_0_726;
   wire n_8_0_727;
   wire n_8_0_728;
   wire n_8_0_729;
   wire n_8_0_730;
   wire n_8_0_731;
   wire n_8_0_732;
   wire n_8_0_733;
   wire n_8_0_734;
   wire n_8_0_735;
   wire n_8_0_736;
   wire n_8_0_737;
   wire n_8_0_738;
   wire n_8_0_739;
   wire n_8_0_740;
   wire n_8_0_741;
   wire n_8_0_742;
   wire n_8_0_743;
   wire n_8_0_744;
   wire n_8_0_745;
   wire n_8_0_746;
   wire n_8_0_747;
   wire n_8_0_748;
   wire n_8_0_749;
   wire n_8_0_750;
   wire n_8_0_751;
   wire n_8_0_752;
   wire n_8_0_753;
   wire n_8_0_754;
   wire n_8_0_755;
   wire n_8_0_756;
   wire n_8_0_757;
   wire n_8_0_758;
   wire n_8_0_759;
   wire n_8_0_760;
   wire n_8_0_761;
   wire n_8_0_762;
   wire n_8_0_763;
   wire n_8_0_764;
   wire n_8_0_765;
   wire n_8_0_766;
   wire n_8_0_767;
   wire n_8_0_768;
   wire n_8_0_769;
   wire n_8_0_770;
   wire n_8_0_771;
   wire n_8_0_772;
   wire n_8_0_773;
   wire n_8_0_774;
   wire n_8_0_775;
   wire n_8_0_776;
   wire n_8_0_777;
   wire n_8_0_778;
   wire n_8_0_779;
   wire n_8_0_780;
   wire n_8_0_781;
   wire n_8_0_782;
   wire n_8_0_783;
   wire n_8_0_784;
   wire n_8_0_785;
   wire n_8_0_786;
   wire n_8_0_787;
   wire n_8_0_788;
   wire n_8_0_789;
   wire n_8_0_790;
   wire n_8_0_791;
   wire n_8_0_792;
   wire n_8_0_793;
   wire n_8_0_794;
   wire n_8_0_795;
   wire n_8_0_796;
   wire n_8_0_797;
   wire n_8_0_798;
   wire n_8_0_799;
   wire n_8_0_800;
   wire n_8_0_801;
   wire n_8_0_802;
   wire n_8_0_803;
   wire n_8_0_804;
   wire n_8_0_805;
   wire n_8_0_806;
   wire n_8_0_807;
   wire n_8_0_808;
   wire n_8_0_809;
   wire n_8_0_810;
   wire n_8_0_811;
   wire n_8_0_812;
   wire n_8_0_813;
   wire n_8_0_814;
   wire n_8_0_815;
   wire n_8_0_816;
   wire n_8_0_817;
   wire n_8_0_818;
   wire n_8_0_819;
   wire n_8_0_820;
   wire n_8_0_821;
   wire n_8_0_822;
   wire n_8_0_823;
   wire n_8_0_824;
   wire n_8_0_825;
   wire n_8_0_826;
   wire n_8_0_827;
   wire n_8_0_828;
   wire n_8_0_829;
   wire n_8_0_830;
   wire n_8_0_831;
   wire n_8_0_832;
   wire n_8_0_833;
   wire n_8_0_834;
   wire n_8_0_835;
   wire n_8_0_836;
   wire n_8_0_837;
   wire n_8_0_838;
   wire n_8_0_839;
   wire n_8_0_840;
   wire n_8_0_841;
   wire n_8_0_842;
   wire n_8_0_843;
   wire n_8_0_844;
   wire n_8_0_845;
   wire n_8_0_846;
   wire n_8_0_847;
   wire n_8_0_848;
   wire n_8_0_849;
   wire n_8_0_850;
   wire n_8_0_851;
   wire n_8_0_852;
   wire n_8_0_853;
   wire n_8_0_854;
   wire n_8_0_855;
   wire n_8_0_856;
   wire n_8_0_857;
   wire n_8_0_858;
   wire n_8_0_859;
   wire n_8_0_860;
   wire n_8_0_861;
   wire n_8_0_862;
   wire n_8_0_863;
   wire n_8_0_864;
   wire n_8_0_865;
   wire n_8_0_866;
   wire n_8_0_867;
   wire n_8_0_868;
   wire n_8_0_869;
   wire n_8_0_870;
   wire n_8_0_871;
   wire n_8_0_872;
   wire n_8_0_873;
   wire n_8_0_874;
   wire n_8_0_875;
   wire n_8_0_876;
   wire n_8_0_877;
   wire n_8_0_878;
   wire n_8_0_879;
   wire n_8_0_880;
   wire n_8_0_881;
   wire n_8_0_882;
   wire n_8_0_883;
   wire n_8_0_884;
   wire n_8_0_885;
   wire n_8_0_886;
   wire n_8_0_887;
   wire n_8_0_888;
   wire n_8_0_889;
   wire n_8_0_890;
   wire n_8_0_891;
   wire n_8_0_892;
   wire n_8_0_893;
   wire n_8_0_894;
   wire n_8_0_895;
   wire n_8_0_896;
   wire n_8_0_897;
   wire n_8_0_898;
   wire n_8_0_899;
   wire n_8_0_900;
   wire n_8_0_901;
   wire n_8_0_902;
   wire n_8_0_903;
   wire n_8_0_904;
   wire n_8_0_905;
   wire n_8_0_906;
   wire n_8_0_907;
   wire n_8_0_908;
   wire n_8_0_909;
   wire n_8_0_910;
   wire n_8_0_911;
   wire n_8_0_912;
   wire n_8_0_913;
   wire n_8_0_914;
   wire n_8_0_915;
   wire n_8_0_916;
   wire n_8_0_917;
   wire n_8_0_918;
   wire n_8_0_919;
   wire n_8_0_920;
   wire n_8_0_921;
   wire n_8_0_922;
   wire n_8_0_923;
   wire n_8_0_924;
   wire n_8_0_925;
   wire n_8_0_926;
   wire n_8_0_927;
   wire n_8_0_928;
   wire n_8_0_929;
   wire n_8_0_930;
   wire n_8_0_931;
   wire n_8_0_932;
   wire n_8_0_933;
   wire n_8_0_934;
   wire n_8_0_935;
   wire n_8_0_936;
   wire n_8_0_937;
   wire n_8_0_938;
   wire n_8_0_939;
   wire n_8_0_940;
   wire n_8_0_941;
   wire n_8_0_942;
   wire n_8_0_943;
   wire n_8_0_944;
   wire n_8_0_945;
   wire n_8_0_946;
   wire n_8_0_947;
   wire n_8_0_948;
   wire n_8_0_949;
   wire n_8_0_950;
   wire n_8_0_951;
   wire n_8_0_952;
   wire n_8_0_953;
   wire n_8_0_954;
   wire n_8_0_955;
   wire n_8_0_956;
   wire n_8_0_957;
   wire n_8_0_958;
   wire n_8_0_959;
   wire n_8_0_960;
   wire n_8_0_961;
   wire n_8_0_962;
   wire n_8_0_963;
   wire n_8_0_964;
   wire n_8_0_965;
   wire n_8_0_966;
   wire n_8_0_967;
   wire n_8_0_968;
   wire n_8_0_969;
   wire n_8_0_970;
   wire n_8_0_971;
   wire n_8_0_972;
   wire n_8_0_973;
   wire n_8_0_974;
   wire n_8_0_975;
   wire n_8_0_976;
   wire n_8_0_977;
   wire n_8_0_978;
   wire n_8_0_979;
   wire n_8_0_980;
   wire n_8_0_981;
   wire n_8_0_982;
   wire n_8_0_983;
   wire n_8_0_984;
   wire n_8_0_985;
   wire n_8_0_986;
   wire n_8_0_987;
   wire n_8_0_988;
   wire n_8_0_989;
   wire n_8_0_990;
   wire n_8_0_991;
   wire n_8_0_992;
   wire n_8_0_993;
   wire n_8_0_994;
   wire n_8_0_995;
   wire n_8_0_996;
   wire n_8_0_997;
   wire n_8_0_998;
   wire n_8_0_999;
   wire n_8_0_1416;
   wire n_8_0_1000;
   wire n_8_0_1001;
   wire n_8_0_1002;
   wire n_8_0_1003;
   wire n_8_0_1004;
   wire n_8_0_1005;
   wire n_8_0_1006;
   wire n_8_0_1007;
   wire n_8_0_1008;
   wire n_8_0_1009;
   wire n_8_0_1010;
   wire n_8_0_1011;
   wire n_8_0_1012;
   wire n_8_0_1013;
   wire n_8_0_1014;
   wire n_8_0_1015;
   wire n_8_0_1016;
   wire n_8_0_1017;
   wire n_8_0_1018;
   wire n_8_0_1019;
   wire n_8_0_1020;
   wire n_8_0_1021;
   wire n_8_0_1022;
   wire n_8_0_1023;
   wire n_8_0_1024;
   wire n_8_0_1025;
   wire n_8_0_1026;
   wire n_8_0_1027;
   wire n_8_0_1028;
   wire n_8_0_1029;
   wire n_8_0_1030;
   wire n_8_0_1031;
   wire n_8_0_1032;
   wire n_8_0_1033;
   wire n_8_0_1034;
   wire n_8_0_1035;
   wire n_8_0_1036;
   wire n_8_0_1037;
   wire n_8_0_1038;
   wire n_8_0_1039;
   wire n_8_0_1040;
   wire n_8_0_1041;
   wire n_8_0_1042;
   wire n_8_0_1043;
   wire n_8_0_1044;
   wire n_8_0_1045;
   wire n_8_0_1046;
   wire n_8_0_1047;
   wire n_8_0_1417;
   wire n_8_0_1048;
   wire n_8_0_1049;
   wire n_8_0_1050;
   wire n_8_0_1051;
   wire n_8_0_1052;
   wire n_8_0_1053;
   wire n_8_0_1054;
   wire n_8_0_1055;
   wire n_8_0_1056;
   wire n_8_0_1057;
   wire n_8_0_1058;
   wire n_8_0_1059;
   wire n_8_0_1060;
   wire n_8_0_1061;
   wire n_8_0_1062;
   wire n_8_0_1063;
   wire n_8_0_1064;
   wire n_8_0_1065;
   wire n_8_0_1066;
   wire n_8_0_1067;
   wire n_8_0_1068;
   wire n_8_0_1069;
   wire n_8_0_1070;
   wire n_8_0_1071;
   wire n_8_0_1072;
   wire n_8_0_1073;
   wire n_8_0_1074;
   wire n_8_0_1418;
   wire n_8_0_1075;
   wire n_8_0_1076;
   wire n_8_0_1077;
   wire n_8_0_1078;
   wire n_8_0_1079;
   wire n_8_0_1080;
   wire n_8_0_1081;
   wire n_8_0_1082;
   wire n_8_0_1083;
   wire n_8_0_1084;
   wire n_8_0_1085;
   wire n_8_0_1086;
   wire n_8_0_1087;
   wire n_8_0_1088;
   wire n_8_0_1089;
   wire n_8_0_1090;
   wire n_8_0_1091;
   wire n_8_0_1092;
   wire n_8_0_1093;
   wire n_8_0_1094;
   wire n_8_0_1095;
   wire n_8_0_1096;
   wire n_8_0_1097;
   wire n_8_0_1098;
   wire n_8_0_1099;
   wire n_8_0_1100;
   wire n_8_0_1101;
   wire n_8_0_1102;
   wire n_8_0_1103;
   wire n_8_0_1104;
   wire n_8_0_1105;
   wire n_8_0_1106;
   wire n_8_0_1107;
   wire n_8_0_1108;
   wire n_8_0_1109;
   wire n_8_0_1110;
   wire n_8_0_1111;
   wire n_8_0_1112;
   wire n_8_0_1113;
   wire n_8_0_1114;
   wire n_8_0_1115;
   wire n_8_0_1116;
   wire n_8_0_1117;
   wire n_8_0_1118;
   wire n_8_0_1119;
   wire n_8_0_1120;
   wire n_8_0_1121;
   wire n_8_0_1122;
   wire n_8_0_1123;
   wire n_8_0_1124;
   wire n_8_0_1125;
   wire n_8_0_1126;
   wire n_8_0_1127;
   wire n_8_0_1128;
   wire n_8_0_1129;
   wire n_8_0_1130;
   wire n_8_0_1131;
   wire n_8_0_1132;
   wire n_8_0_1133;
   wire n_8_0_1134;
   wire n_8_0_1135;
   wire n_8_0_1136;
   wire n_8_0_1137;
   wire n_8_0_1138;
   wire n_8_0_1139;
   wire n_8_0_1140;
   wire n_8_0_1141;
   wire n_8_0_1142;
   wire n_8_0_1143;
   wire n_8_0_1144;
   wire n_8_0_1145;
   wire n_8_0_1146;
   wire n_8_0_1147;
   wire n_8_0_1148;
   wire n_8_0_1149;
   wire n_8_0_1150;
   wire n_8_0_1151;
   wire n_8_0_1152;
   wire n_8_0_1153;
   wire n_8_0_1154;
   wire n_8_0_1155;
   wire n_8_0_1156;
   wire n_8_0_1157;
   wire n_8_0_1158;
   wire n_8_0_1159;
   wire n_8_0_1160;
   wire n_8_0_1161;
   wire n_8_0_1162;
   wire n_8_0_1163;
   wire n_8_0_1164;
   wire n_8_0_1165;
   wire n_8_0_1166;
   wire n_8_0_1419;
   wire n_8_0_1420;
   wire n_8_0_1421;
   wire n_8_0_1422;
   wire n_8_0_1423;
   wire n_8_0_1424;
   wire n_8_0_1425;
   wire n_8_0_1426;
   wire n_8_0_1427;
   wire n_8_0_1428;
   wire n_8_0_1429;
   wire n_8_0_1430;
   wire n_8_0_1431;
   wire n_8_0_1432;
   wire n_8_0_1433;
   wire n_8_0_1434;
   wire n_8_0_1435;
   wire n_8_0_1436;
   wire n_8_0_1437;
   wire n_8_0_1438;
   wire n_8_0_1439;
   wire n_8_0_1440;
   wire n_8_0_1441;
   wire n_8_0_1442;
   wire n_8_0_1443;
   wire n_8_0_1444;
   wire n_8_0_1445;
   wire n_8_0_1446;
   wire n_8_0_1447;
   wire n_8_0_1448;
   wire n_8_0_1449;
   wire n_8_0_1450;
   wire n_8_0_1451;
   wire n_8_0_1452;
   wire n_8_0_1453;
   wire n_8_0_1454;
   wire n_8_0_1455;
   wire n_8_0_1456;
   wire n_8_0_1457;
   wire n_8_0_1458;
   wire n_8_0_1459;
   wire n_8_0_1460;
   wire n_8_0_1461;
   wire n_8_0_1462;
   wire n_8_0_1463;
   wire n_8_0_1464;
   wire n_8_0_1465;
   wire n_8_0_1466;
   wire n_8_0_1467;
   wire n_8_0_1468;
   wire n_8_0_1469;
   wire n_8_0_1470;
   wire n_8_0_1471;
   wire n_8_0_1472;
   wire n_8_0_1473;
   wire n_8_0_1474;
   wire n_8_0_1475;
   wire n_8_0_1476;
   wire n_8_0_1477;
   wire n_8_0_1478;
   wire n_8_0_1479;
   wire n_8_0_1480;
   wire n_8_0_1481;
   wire n_8_0_1482;
   wire n_8_0_1483;
   wire n_8_0_1485;
   wire n_8_0_1486;
   wire n_8_0_1487;
   wire n_8_0_1488;
   wire n_8_0_1489;
   wire n_8_0_1490;
   wire n_8_0_1491;
   wire n_8_0_1492;
   wire n_8_0_1493;
   wire n_8_0_1494;
   wire n_8_0_1495;
   wire n_8_0_1496;
   wire n_8_0_1497;
   wire n_8_0_1498;
   wire n_8_0_1499;
   wire n_8_0_1500;
   wire n_8_0_1501;
   wire n_8_0_1502;
   wire n_8_0_1503;
   wire n_8_0_1504;
   wire n_8_0_1505;
   wire n_8_0_1506;
   wire n_8_0_1507;
   wire n_8_0_1508;
   wire n_8_0_1509;
   wire n_8_0_1510;
   wire n_8_0_1511;
   wire n_8_0_1512;
   wire n_8_0_1513;
   wire n_8_0_1514;
   wire n_8_0_1515;
   wire n_8_0_1516;
   wire n_8_0_1517;
   wire n_8_0_1518;
   wire n_8_0_1519;
   wire n_8_0_1520;
   wire n_8_0_1521;
   wire n_8_0_1522;
   wire n_8_0_1523;
   wire n_8_0_1524;
   wire n_8_0_1525;
   wire n_8_0_1526;
   wire n_8_0_1530;
   wire n_8_0_1531;
   wire n_8_0_1532;
   wire n_8_0_1533;
   wire n_8_0_1534;
   wire n_8_0_1535;
   wire n_8_0_1536;
   wire n_8_0_1537;
   wire n_8_0_1538;
   wire n_8_0_1539;
   wire n_8_0_1540;
   wire n_8_0_1541;
   wire n_8_0_1542;
   wire n_8_0_1543;
   wire n_8_0_1544;
   wire n_8_0_1545;
   wire n_8_0_1546;
   wire n_8_0_1547;
   wire n_8_0_1548;
   wire n_8_0_1549;
   wire n_8_0_1550;
   wire n_8_0_1551;
   wire n_8_0_1552;
   wire n_8_0_1553;
   wire n_8_0_1554;
   wire n_8_0_1555;
   wire n_8_0_1556;
   wire n_8_0_1557;
   wire n_8_0_1558;
   wire n_8_0_1559;
   wire n_8_0_1560;
   wire n_8_0_1561;
   wire n_8_0_1562;
   wire n_8_0_1563;
   wire n_8_0_1564;
   wire n_8_0_1565;
   wire n_8_0_1566;
   wire n_8_0_1567;
   wire n_8_0_1568;
   wire n_8_0_1569;
   wire n_8_0_1570;
   wire n_8_0_1571;
   wire n_8_0_1572;
   wire n_8_0_1573;
   wire n_8_0_1574;
   wire n_8_0_1575;
   wire n_8_0_1576;
   wire n_8_0_1577;
   wire n_8_0_1578;
   wire n_8_0_1579;
   wire n_8_0_1580;
   wire n_8_0_1581;
   wire n_8_0_1582;
   wire n_8_0_1583;
   wire n_8_0_1584;
   wire n_8_0_1585;
   wire n_8_0_1586;
   wire n_8_0_1587;
   wire n_8_0_1588;
   wire n_8_0_1591;
   wire n_8_0_1592;
   wire n_8_0_1593;
   wire n_8_0_1594;
   wire n_8_0_1595;
   wire n_8_0_1596;
   wire n_8_0_1597;
   wire n_8_0_1598;
   wire n_8_0_1601;
   wire n_8_0_1602;
   wire n_8_0_1603;
   wire n_8_0_1604;
   wire n_8_0_1605;
   wire n_8_0_1606;
   wire n_8_0_1608;
   wire n_8_0_1609;
   wire n_8_0_1610;
   wire n_8_0_1611;
   wire n_8_0_1612;
   wire n_8_0_1613;
   wire n_8_0_1614;
   wire n_8_0_1615;
   wire n_8_0_1618;
   wire n_8_0_1619;
   wire n_8_0_1620;
   wire n_8_0_1621;
   wire n_8_0_1622;
   wire n_8_0_1623;
   wire n_8_0_1624;
   wire n_8_0_1625;
   wire n_8_0_1626;
   wire n_8_0_1627;
   wire n_8_0_1628;
   wire n_8_0_1629;
   wire n_8_0_1630;
   wire n_8_0_1631;
   wire n_8_0_1632;
   wire n_8_0_1633;
   wire n_8_0_1634;
   wire n_8_0_1635;
   wire n_8_0_1636;
   wire n_8_0_1637;
   wire n_8_0_1638;
   wire n_8_0_1639;
   wire n_8_0_1640;
   wire n_8_0_1641;
   wire n_8_0_1642;
   wire n_8_0_1643;
   wire n_8_0_1644;
   wire n_8_0_1645;
   wire n_8_0_1646;
   wire n_8_0_1647;
   wire n_8_0_1648;
   wire n_8_0_1649;
   wire n_8_0_1650;
   wire n_8_0_1651;
   wire n_8_0_1652;
   wire n_8_0_1653;
   wire n_8_0_1654;
   wire n_8_0_1655;
   wire n_8_0_1658;
   wire n_8_0_1659;
   wire n_8_0_1660;
   wire n_8_0_1661;
   wire n_8_0_1662;
   wire n_8_0_1663;
   wire n_8_0_1664;
   wire n_8_0_1665;
   wire n_8_0_1666;
   wire n_8_0_1667;
   wire n_8_0_1668;
   wire n_8_0_1669;
   wire n_8_0_1670;
   wire n_8_0_1671;
   wire n_8_0_1672;
   wire n_8_0_1673;
   wire n_8_0_1674;
   wire n_8_0_1675;
   wire n_8_0_1676;
   wire n_8_0_1677;
   wire n_8_0_1678;
   wire n_8_0_1679;
   wire n_8_0_1680;
   wire n_8_0_1681;
   wire n_8_0_1682;
   wire n_8_0_1683;
   wire n_8_0_1684;
   wire n_8_0_1685;
   wire n_8_0_1686;
   wire n_8_0_1687;
   wire n_8_0_1688;
   wire n_8_0_1689;
   wire n_8_0_1690;
   wire n_8_0_1691;
   wire n_8_0_1692;
   wire n_8_0_1693;
   wire n_8_0_1694;
   wire n_8_0_1695;
   wire n_8_0_1696;
   wire n_8_0_1697;
   wire n_8_0_1698;
   wire n_8_0_1699;
   wire n_8_0_1700;
   wire n_8_0_1701;
   wire n_8_0_1702;
   wire n_8_0_1703;
   wire n_8_0_1704;
   wire n_8_0_1705;
   wire n_8_0_1706;
   wire n_8_0_1707;
   wire n_8_0_1708;
   wire n_8_0_1709;
   wire n_8_0_1710;
   wire n_8_0_1711;
   wire n_8_0_1712;
   wire n_8_0_1713;
   wire n_8_0_1714;
   wire n_8_0_1715;
   wire n_8_0_1716;
   wire n_8_0_1717;
   wire n_8_0_1718;
   wire n_8_0_1719;
   wire n_8_0_1720;
   wire n_8_0_1721;
   wire n_8_0_1722;
   wire n_8_0_1723;
   wire n_8_0_1724;
   wire n_8_0_1725;
   wire n_8_0_1726;
   wire n_8_0_1727;
   wire n_8_0_1728;
   wire n_8_0_1729;
   wire n_8_0_1730;
   wire n_8_0_1731;
   wire n_8_0_1732;
   wire n_8_0_1733;
   wire n_8_0_1738;
   wire n_8_0_1739;
   wire n_8_0_1740;
   wire n_8_0_1741;
   wire n_8_0_1742;
   wire n_8_0_1743;
   wire n_8_0_1744;
   wire n_8_0_1745;
   wire n_8_0_1746;
   wire n_8_0_1747;
   wire n_8_0_1748;
   wire n_8_0_1749;
   wire n_8_0_1750;
   wire n_8_0_1751;
   wire n_8_0_1752;
   wire n_8_0_1756;
   wire n_8_0_1757;
   wire n_8_0_1758;
   wire n_8_0_1759;
   wire n_8_0_1760;
   wire n_8_0_1761;
   wire n_8_0_1762;
   wire n_8_0_1763;
   wire n_8_0_1764;
   wire n_8_0_1765;
   wire n_8_0_1766;
   wire n_8_0_1767;
   wire n_8_0_1768;
   wire n_8_0_1769;
   wire n_8_0_1770;
   wire n_8_0_1771;
   wire n_8_0_1772;
   wire n_8_0_1773;
   wire n_8_0_1775;
   wire n_8_0_1776;
   wire n_8_0_1777;
   wire n_8_0_1778;
   wire n_8_0_1779;
   wire n_8_0_1780;
   wire n_8_0_1781;
   wire n_8_0_1784;
   wire n_8_0_1785;
   wire n_8_0_1786;
   wire n_8_0_1787;
   wire n_8_0_1788;
   wire n_8_0_1789;
   wire n_8_0_1790;
   wire n_8_0_1791;
   wire n_8_0_1792;
   wire n_8_0_1793;
   wire n_8_0_1794;
   wire n_8_0_1795;
   wire n_8_0_1796;
   wire n_8_0_1797;
   wire n_8_0_1798;
   wire n_8_0_1799;
   wire n_8_0_1800;
   wire n_8_0_1801;
   wire n_8_0_1802;
   wire n_8_0_1803;
   wire n_8_0_1804;
   wire n_8_0_1805;
   wire n_8_0_1806;
   wire n_8_0_1807;
   wire n_8_0_1808;
   wire n_8_0_1809;
   wire n_8_0_1810;
   wire n_8_0_1811;
   wire n_8_0_1812;
   wire n_8_0_1813;
   wire n_8_0_1814;
   wire n_8_0_1815;
   wire n_8_0_1816;
   wire n_8_0_1817;
   wire n_8_0_1818;
   wire n_8_0_1819;
   wire n_8_0_1820;
   wire n_8_0_1821;
   wire n_8_0_1822;
   wire n_8_0_1823;
   wire n_8_0_1824;
   wire n_8_0_1825;
   wire n_8_0_1826;
   wire n_8_0_1827;
   wire n_8_0_1828;
   wire n_8_0_1829;
   wire n_8_0_1830;
   wire n_8_0_1831;
   wire n_8_0_1832;
   wire n_8_0_1833;
   wire n_8_0_1834;
   wire n_8_0_1835;
   wire n_8_0_1836;
   wire n_8_0_1837;
   wire n_8_0_1838;
   wire n_8_0_1839;
   wire n_8_0_1840;
   wire n_8_0_1841;
   wire n_8_0_1842;
   wire n_8_0_1843;
   wire n_8_0_1844;
   wire n_8_0_1845;
   wire n_8_0_1846;
   wire n_8_0_1847;
   wire n_8_0_1848;
   wire n_8_0_1849;
   wire n_8_0_1850;
   wire n_8_0_1851;
   wire n_8_0_1852;
   wire n_8_0_1853;
   wire n_8_0_1854;
   wire n_8_0_1855;
   wire n_8_0_1856;
   wire n_8_0_1857;
   wire n_8_0_1858;
   wire n_8_0_1859;
   wire n_8_0_1860;
   wire n_8_0_1861;
   wire n_8_0_1862;
   wire n_8_0_1863;
   wire n_8_0_1864;
   wire n_8_0_1865;
   wire n_8_0_1866;
   wire n_8_0_1867;
   wire n_8_0_1868;
   wire n_8_0_1869;
   wire n_8_0_1870;
   wire n_8_0_1871;
   wire n_8_0_1872;
   wire n_8_0_1874;
   wire n_8_0_1875;
   wire n_8_0_1876;
   wire n_8_0_1877;
   wire n_8_0_1878;
   wire n_8_0_1879;
   wire n_8_0_1880;
   wire n_8_0_1881;
   wire n_8_0_1882;
   wire n_8_0_1885;
   wire n_8_0_1886;
   wire n_8_0_1887;
   wire n_8_0_1888;
   wire n_8_0_1889;
   wire n_8_0_1890;
   wire n_8_0_1891;
   wire n_8_0_1892;
   wire n_8_0_1893;
   wire n_8_0_1894;
   wire n_8_0_1895;
   wire n_8_0_1896;
   wire n_8_0_1897;
   wire n_8_0_1898;
   wire n_8_0_1899;
   wire n_8_0_1900;
   wire n_8_0_1901;
   wire n_8_0_1902;
   wire n_8_0_1903;
   wire n_8_0_1906;
   wire n_8_0_1907;
   wire n_8_0_1908;
   wire n_8_0_1909;
   wire n_8_0_1910;
   wire n_8_0_1911;
   wire n_8_0_1912;
   wire n_8_0_1913;
   wire n_8_0_1914;
   wire n_8_0_1915;
   wire n_8_0_1916;
   wire n_8_0_1917;
   wire n_8_0_1918;
   wire n_8_0_1919;
   wire n_8_0_1920;
   wire n_8_0_1921;
   wire n_8_0_1922;
   wire n_8_0_1923;
   wire n_8_0_1924;
   wire n_8_0_1925;
   wire n_8_0_1926;
   wire n_8_0_1927;
   wire n_8_0_1928;
   wire n_8_0_1929;
   wire n_8_0_1930;
   wire n_8_0_1931;
   wire n_8_0_1932;
   wire n_8_0_1933;
   wire n_8_0_1934;
   wire n_8_0_1935;
   wire n_8_0_1936;
   wire n_8_0_1937;
   wire n_8_0_1938;
   wire n_8_0_1939;
   wire n_8_0_1940;
   wire n_8_0_1941;
   wire n_8_0_1942;
   wire n_8_0_1943;
   wire n_8_0_1947;
   wire n_8_0_1948;
   wire n_8_0_1949;
   wire n_8_0_1950;
   wire n_8_0_1951;
   wire n_8_0_1952;
   wire n_8_0_1953;
   wire n_8_0_1954;
   wire n_8_0_1955;
   wire n_8_0_1956;
   wire n_8_0_1957;
   wire n_8_0_1958;
   wire n_8_0_1959;
   wire n_8_0_1960;
   wire n_8_0_1961;
   wire n_8_0_1962;
   wire n_8_0_1963;
   wire n_8_0_1964;
   wire n_8_0_1965;
   wire n_8_0_1966;
   wire n_8_0_1967;
   wire n_8_0_1968;
   wire n_8_0_1969;
   wire n_8_0_1970;
   wire n_8_0_1971;
   wire n_8_0_1974;
   wire n_8_0_1975;
   wire n_8_0_1976;
   wire n_8_0_1977;
   wire n_8_0_1978;
   wire n_8_0_1979;
   wire n_8_0_1980;
   wire n_8_0_1981;
   wire n_8_0_1982;
   wire n_8_0_1983;
   wire n_8_0_1984;
   wire n_8_0_1985;
   wire n_8_0_1986;
   wire n_8_0_1987;
   wire n_8_0_1988;
   wire n_8_0_1989;
   wire n_8_0_1990;
   wire n_8_0_1991;
   wire n_8_0_1992;
   wire n_8_0_1993;
   wire n_8_0_1994;
   wire n_8_0_1995;
   wire n_8_0_1996;
   wire n_8_0_1997;
   wire n_8_0_1998;
   wire n_8_0_1999;
   wire n_8_0_2000;
   wire n_8_0_2001;
   wire n_8_0_2002;
   wire n_8_0_2003;
   wire n_8_0_2004;
   wire n_8_0_2005;
   wire n_8_0_2006;
   wire n_8_0_2007;
   wire n_8_0_2008;
   wire n_8_0_2009;
   wire n_8_0_2010;
   wire n_8_0_2011;
   wire n_8_0_2012;
   wire n_8_0_2013;
   wire n_8_0_2014;
   wire n_8_0_2015;
   wire n_8_0_2016;
   wire n_8_0_2017;
   wire n_8_0_2018;
   wire n_8_0_2019;
   wire n_8_0_2020;
   wire n_8_0_2021;
   wire n_8_0_2022;
   wire n_8_0_2023;
   wire n_8_0_2024;
   wire n_8_0_2025;
   wire n_8_0_2026;
   wire n_8_0_2027;
   wire n_8_0_2028;
   wire n_8_0_2029;
   wire n_8_0_2030;
   wire n_8_0_2031;
   wire n_8_0_2032;
   wire n_8_0_2033;
   wire n_8_0_2034;
   wire n_8_0_2035;
   wire n_8_0_2036;
   wire n_8_0_2037;
   wire n_8_0_2038;
   wire n_8_0_2039;
   wire n_8_0_2040;
   wire n_8_0_2041;
   wire n_8_0_2042;
   wire n_8_0_2043;
   wire n_8_0_2044;
   wire n_8_0_2045;
   wire n_8_0_2046;
   wire n_8_0_2047;
   wire n_8_0_2048;
   wire n_8_0_2049;
   wire n_8_0_2050;
   wire n_8_0_2051;
   wire n_8_0_2052;
   wire n_8_0_2053;
   wire n_8_0_2054;
   wire n_8_0_2055;
   wire n_8_0_2056;
   wire n_8_0_2057;
   wire n_8_0_2058;
   wire n_8_0_2059;
   wire n_8_0_2060;
   wire n_8_0_2061;
   wire n_8_0_2062;
   wire n_8_0_2063;
   wire n_8_0_2064;
   wire n_8_0_2065;
   wire n_8_0_2066;
   wire n_8_0_2067;
   wire n_8_0_2068;
   wire n_8_0_2069;
   wire n_8_0_2070;
   wire n_8_0_2071;
   wire n_8_0_2072;
   wire n_8_0_2073;
   wire n_8_0_2074;
   wire n_8_0_2075;
   wire n_8_0_2076;
   wire n_8_0_2077;
   wire n_8_0_2078;
   wire n_8_0_2079;
   wire n_8_0_2080;
   wire n_8_0_2081;
   wire n_8_0_2082;
   wire n_8_0_2083;
   wire n_8_0_2084;
   wire n_8_0_2085;
   wire n_8_0_2086;
   wire n_8_0_2087;
   wire n_8_0_2088;
   wire n_8_0_2089;
   wire n_8_0_2090;
   wire n_8_0_2091;
   wire n_8_0_2092;
   wire n_8_0_2093;
   wire n_8_0_2094;
   wire n_8_0_2095;
   wire n_8_0_2096;
   wire n_8_0_2097;
   wire n_8_0_2098;
   wire n_8_0_2099;
   wire n_8_0_2100;
   wire n_8_0_2101;
   wire n_8_0_2102;
   wire n_8_0_2103;
   wire n_8_0_2104;
   wire n_8_0_2105;
   wire n_8_0_2106;
   wire n_8_0_2107;
   wire n_8_0_2108;
   wire n_8_0_2109;
   wire n_8_0_2110;
   wire n_8_0_2111;
   wire n_8_0_2112;
   wire n_8_0_2113;
   wire n_8_0_2114;
   wire n_8_0_2115;
   wire n_8_0_2116;
   wire n_8_0_2117;
   wire n_8_0_2118;
   wire n_8_0_2119;
   wire n_8_0_2120;
   wire n_8_0_2121;
   wire n_8_0_2122;
   wire n_8_0_2123;
   wire n_8_0_2124;
   wire n_8_0_2125;
   wire n_8_0_2126;
   wire n_8_0_2127;
   wire n_8_0_2128;
   wire n_8_0_2129;
   wire n_8_0_2130;
   wire n_8_0_2131;
   wire n_8_0_2132;
   wire n_8_0_2133;
   wire n_8_0_2134;
   wire n_8_0_2135;
   wire n_8_0_2136;
   wire n_8_0_2137;
   wire n_8_0_2138;
   wire n_8_0_2139;
   wire n_8_0_2140;
   wire n_8_0_2141;
   wire n_8_0_2142;
   wire n_8_0_2143;
   wire n_8_0_2144;
   wire n_8_0_2145;
   wire n_8_0_2146;
   wire n_8_0_2147;
   wire n_8_0_2148;
   wire n_8_0_2149;
   wire n_8_0_2150;
   wire n_8_0_2151;
   wire n_8_0_2152;
   wire n_8_0_2153;
   wire n_8_0_2154;
   wire n_8_0_2155;
   wire n_8_0_2156;
   wire n_8_0_2157;
   wire n_8_0_2158;
   wire n_8_0_2159;
   wire n_8_0_2160;
   wire n_8_0_2161;
   wire n_8_0_2162;
   wire n_8_0_2163;
   wire n_8_0_2164;
   wire n_8_0_2165;
   wire n_8_0_2166;
   wire n_8_0_2167;
   wire n_8_0_2168;
   wire n_8_0_2169;
   wire n_8_0_2170;
   wire n_8_0_2171;
   wire n_8_0_2172;
   wire n_8_0_2173;
   wire n_8_0_2174;
   wire n_8_0_2175;
   wire n_8_0_2176;
   wire n_8_0_2177;
   wire n_8_0_2178;
   wire n_8_0_2179;
   wire n_8_0_2180;
   wire n_8_0_2181;
   wire n_8_0_2182;
   wire n_8_0_2183;
   wire n_8_0_2184;
   wire n_8_0_2185;
   wire n_8_0_2186;
   wire n_8_0_2187;
   wire n_8_0_2188;
   wire n_8_0_2189;
   wire n_8_0_2190;
   wire n_8_0_2191;
   wire n_8_0_2192;
   wire n_8_0_2193;
   wire n_8_0_2194;
   wire n_8_0_2195;
   wire n_8_0_2196;
   wire n_8_0_2197;
   wire n_8_0_2198;
   wire n_8_0_2199;
   wire n_8_0_2200;
   wire n_8_0_2201;
   wire n_8_0_2202;
   wire n_8_0_2203;
   wire n_8_0_2204;
   wire n_8_0_2205;
   wire n_8_0_2206;
   wire n_8_0_2207;
   wire n_8_0_2208;
   wire n_8_0_2209;
   wire n_8_0_2210;
   wire n_8_0_2211;
   wire n_8_0_2212;
   wire n_8_0_2213;
   wire n_8_0_2214;
   wire n_8_0_2215;
   wire n_8_0_2216;
   wire n_8_0_2217;
   wire n_8_0_2218;
   wire n_8_0_2219;
   wire n_8_0_2220;
   wire n_8_0_2221;
   wire n_8_0_2222;
   wire n_8_0_2223;
   wire n_8_0_2224;
   wire n_8_0_2225;
   wire n_8_0_2226;
   wire n_8_0_2227;
   wire n_8_0_2228;
   wire n_8_0_2229;
   wire n_8_0_2230;
   wire n_8_0_2231;
   wire n_8_0_2232;
   wire n_8_0_2233;
   wire n_8_0_2234;
   wire n_8_0_2235;
   wire n_8_0_2236;
   wire n_8_0_2237;
   wire n_8_0_2238;
   wire n_8_0_2239;
   wire n_8_0_2240;
   wire n_8_0_2241;
   wire n_8_0_2242;
   wire n_8_0_2243;
   wire n_8_0_2244;
   wire n_8_0_2245;
   wire n_8_0_2246;
   wire n_8_0_2247;
   wire n_8_0_2248;
   wire n_8_0_2249;
   wire n_8_0_2250;
   wire n_8_0_2251;
   wire n_8_0_2252;
   wire n_8_0_2253;
   wire n_8_0_2254;
   wire n_8_0_2255;
   wire n_8_0_2256;
   wire n_8_0_2257;
   wire n_8_0_2258;
   wire n_8_0_2259;
   wire n_8_0_2260;
   wire n_8_0_2261;
   wire n_8_0_2262;
   wire n_8_0_2263;
   wire n_8_0_2264;
   wire n_8_0_2265;
   wire n_8_0_2266;
   wire n_8_0_2267;
   wire n_8_0_2268;
   wire n_8_0_2269;
   wire n_8_0_2270;
   wire n_8_0_2271;
   wire n_8_0_2272;
   wire n_8_0_2273;
   wire n_8_0_2274;
   wire n_8_0_2275;
   wire n_8_0_2276;
   wire n_8_0_2277;
   wire n_8_0_2278;
   wire n_8_0_2279;
   wire n_8_0_2280;
   wire n_8_0_2281;
   wire n_8_0_2282;
   wire n_8_0_2283;
   wire n_8_0_2284;
   wire n_8_0_2285;
   wire n_8_0_2286;
   wire n_8_0_2287;
   wire n_8_0_2288;
   wire n_8_0_2289;
   wire n_8_0_2290;
   wire n_8_0_2291;
   wire n_8_0_2292;
   wire n_8_0_2293;
   wire n_8_0_2294;
   wire n_8_0_2295;
   wire n_8_0_2296;
   wire n_8_0_2297;
   wire n_8_0_2298;
   wire n_8_0_2299;
   wire n_8_0_2300;
   wire n_8_0_2301;
   wire n_8_0_2302;
   wire n_8_0_2303;
   wire n_8_0_2304;
   wire n_8_0_2305;
   wire n_8_0_2306;
   wire n_8_0_2307;
   wire n_8_0_2308;
   wire n_8_0_2309;
   wire n_8_0_2310;
   wire n_8_0_2311;
   wire n_8_0_2312;
   wire n_8_0_2313;
   wire n_8_0_2314;
   wire n_8_0_2315;
   wire n_8_0_2316;
   wire n_8_0_2317;
   wire n_8_0_2318;
   wire n_8_0_2319;
   wire n_8_0_2320;
   wire n_8_0_2321;
   wire n_8_0_2322;
   wire n_8_0_2323;
   wire n_8_0_2324;
   wire n_8_0_2325;
   wire n_8_0_2326;
   wire n_8_0_2327;
   wire n_8_0_2328;
   wire n_8_0_2329;
   wire n_8_0_2330;
   wire n_8_0_2331;
   wire n_8_0_2332;
   wire n_8_0_2333;
   wire n_8_0_2334;
   wire n_8_0_2335;
   wire n_8_0_2336;
   wire n_8_0_2337;
   wire n_8_0_2338;
   wire n_8_0_2339;
   wire n_8_0_2340;
   wire n_8_0_2341;
   wire n_8_0_2342;
   wire n_8_0_2343;
   wire n_8_0_2344;
   wire n_8_0_2345;
   wire n_8_0_2346;
   wire n_8_0_2347;
   wire n_8_0_2348;
   wire n_8_0_2349;
   wire n_8_0_2350;
   wire n_8_0_2351;
   wire n_8_0_2352;
   wire n_8_0_2353;
   wire n_8_0_2354;
   wire n_8_0_2355;
   wire n_8_0_2356;
   wire n_8_0_2357;
   wire n_8_0_2358;
   wire n_8_0_2359;
   wire n_8_0_2360;
   wire n_8_0_2361;
   wire n_8_0_2362;
   wire n_8_0_2363;
   wire n_8_0_2364;
   wire n_8_0_2365;
   wire n_8_0_2366;
   wire n_8_0_2367;
   wire n_8_0_2368;
   wire n_8_0_2369;
   wire n_8_0_2370;
   wire n_8_0_2371;
   wire n_8_0_2372;
   wire n_8_0_2373;
   wire n_8_0_2374;
   wire n_8_0_2375;
   wire n_8_0_2376;
   wire n_8_0_2377;
   wire n_8_0_2378;
   wire n_8_0_2379;
   wire n_8_0_2380;
   wire n_8_0_2381;
   wire n_8_0_2382;
   wire n_8_0_2383;
   wire n_8_0_2384;
   wire n_8_0_2385;
   wire n_8_0_2386;
   wire n_8_0_2387;
   wire n_8_0_2388;
   wire n_8_0_2389;
   wire n_8_0_2390;
   wire n_8_0_2391;
   wire n_8_0_2392;
   wire n_8_0_2393;
   wire n_8_0_2394;
   wire n_8_0_2395;
   wire n_8_0_2396;
   wire n_8_0_2397;
   wire n_8_0_2398;
   wire n_8_0_2399;
   wire n_8_0_2400;
   wire n_8_0_2401;
   wire n_8_0_2402;
   wire n_8_0_2403;
   wire n_8_0_2404;
   wire n_8_0_2405;
   wire n_8_0_2406;
   wire n_8_0_2407;
   wire n_8_0_2408;
   wire n_8_0_2409;
   wire n_8_0_2410;
   wire n_8_0_2411;
   wire n_8_0_2412;
   wire n_8_0_2413;
   wire n_8_0_2414;
   wire n_8_0_2415;
   wire n_8_0_2416;
   wire n_8_0_2417;
   wire n_8_0_2418;
   wire n_8_0_2419;
   wire n_8_0_2420;
   wire n_8_0_2421;
   wire n_8_0_2422;
   wire n_8_0_2423;
   wire n_8_0_2424;
   wire n_8_0_2425;
   wire n_8_0_2426;
   wire n_8_0_2427;
   wire n_8_0_2428;
   wire n_8_0_2429;
   wire n_8_0_2430;
   wire n_8_0_2431;
   wire n_8_0_2432;
   wire n_8_0_2433;
   wire n_8_0_2434;
   wire n_8_0_2435;
   wire n_8_0_2436;
   wire n_8_0_2437;
   wire n_8_0_2438;
   wire n_8_0_2439;
   wire n_8_0_2440;
   wire n_8_0_2441;
   wire n_8_0_2442;
   wire n_8_0_2443;
   wire n_8_0_2444;
   wire n_8_0_2445;
   wire n_8_0_2446;
   wire n_8_0_2447;
   wire n_8_0_2448;
   wire n_8_0_2449;
   wire n_8_0_2450;
   wire n_8_0_2451;
   wire n_8_0_2452;
   wire n_8_0_2453;
   wire n_8_0_2454;
   wire n_8_0_2455;
   wire n_8_0_2456;
   wire n_8_0_2457;
   wire n_8_0_2458;
   wire n_8_0_2459;
   wire n_8_0_2460;
   wire n_8_0_2461;
   wire n_8_0_2462;
   wire n_8_0_2463;
   wire n_8_0_2464;
   wire n_8_0_2465;
   wire n_8_0_2466;
   wire n_8_0_2467;
   wire n_8_0_2468;
   wire n_8_0_2469;
   wire n_8_0_2470;
   wire n_8_0_2471;
   wire n_8_0_2472;
   wire n_8_0_2473;
   wire n_8_0_2474;
   wire n_8_0_2475;
   wire n_8_0_2476;
   wire n_8_0_2477;
   wire n_8_0_2478;
   wire n_8_0_2479;
   wire n_8_0_2480;
   wire n_8_0_2481;
   wire n_8_0_2482;
   wire n_8_0_2483;
   wire n_8_0_2484;
   wire n_8_0_2485;
   wire n_8_0_2486;
   wire n_8_0_2487;
   wire n_8_0_2488;
   wire n_8_0_2489;
   wire n_8_0_2490;
   wire n_8_0_2491;
   wire n_8_0_2492;
   wire n_8_0_2493;
   wire n_8_0_2494;
   wire n_8_0_2495;
   wire n_8_0_2496;
   wire n_8_0_2497;
   wire n_8_0_2498;
   wire n_8_0_2499;
   wire n_8_0_2500;
   wire n_8_0_2501;
   wire n_8_0_2502;
   wire n_8_0_2503;
   wire n_8_0_2504;
   wire n_8_0_2505;
   wire n_8_0_2506;
   wire n_8_0_2507;
   wire n_8_0_2508;
   wire n_8_0_2509;
   wire n_8_0_2510;
   wire n_8_0_2511;
   wire n_8_0_2512;
   wire n_8_0_2513;
   wire n_8_0_2514;
   wire n_8_0_2515;
   wire n_8_0_2516;
   wire n_8_0_2517;
   wire n_8_0_2518;
   wire n_8_0_2519;
   wire n_8_0_2520;
   wire n_8_0_2521;
   wire n_8_0_2522;
   wire n_8_0_2523;
   wire n_8_0_2524;
   wire n_8_0_2525;
   wire n_8_0_2526;
   wire n_8_0_2527;
   wire n_8_0_2528;
   wire n_8_0_2529;
   wire n_8_0_2530;
   wire n_8_0_2531;
   wire n_8_0_2532;
   wire n_8_0_2533;
   wire n_8_0_2534;
   wire n_8_0_2535;
   wire n_8_0_2536;
   wire n_8_0_2537;
   wire n_8_0_2538;
   wire n_8_0_2539;
   wire n_8_0_2540;
   wire n_8_0_2543;
   wire n_8_0_2546;
   wire n_8_0_2547;
   wire n_8_0_2548;
   wire n_8_0_2549;
   wire n_8_0_2550;
   wire n_8_0_2551;
   wire n_8_0_2552;
   wire n_8_0_2553;
   wire n_8_0_2554;
   wire n_8_0_2555;
   wire n_8_0_2556;
   wire n_8_0_2557;
   wire n_8_0_2558;
   wire n_8_0_2559;
   wire n_8_0_2560;
   wire n_8_0_2561;
   wire n_8_0_2562;
   wire n_8_0_2563;
   wire n_8_0_2564;
   wire n_8_0_2565;
   wire n_8_0_2566;
   wire n_8_0_2567;
   wire n_8_0_2568;
   wire n_8_0_2569;
   wire n_8_0_2570;
   wire n_8_0_2571;
   wire n_8_0_2572;
   wire n_8_0_2573;
   wire n_8_0_2574;
   wire n_8_0_2575;
   wire n_8_0_2576;
   wire n_8_0_2577;
   wire n_8_0_2578;
   wire n_8_0_2579;
   wire n_8_0_2580;
   wire n_8_0_2581;
   wire n_8_0_2582;
   wire n_8_0_2583;
   wire n_8_0_2584;
   wire n_8_0_2585;
   wire n_8_0_2586;
   wire n_8_0_2587;
   wire n_8_0_2588;
   wire n_8_0_2589;
   wire n_8_0_2590;
   wire n_8_0_2591;
   wire n_8_0_2592;
   wire n_8_0_2593;
   wire n_8_0_2594;
   wire n_8_0_2595;
   wire n_8_0_2596;
   wire n_8_0_2597;
   wire n_8_0_2598;
   wire n_8_0_2599;
   wire n_8_0_2600;
   wire n_8_0_2601;
   wire n_8_0_2602;
   wire n_8_0_2603;
   wire n_8_0_2604;
   wire n_8_0_2605;
   wire n_8_0_2606;
   wire n_8_0_2607;
   wire n_8_0_2608;
   wire n_8_0_2609;
   wire n_8_0_2610;
   wire n_8_0_2611;
   wire n_8_0_2612;
   wire n_8_0_2613;
   wire n_8_0_2614;
   wire n_8_0_2615;
   wire n_8_0_2616;
   wire n_8_0_2617;
   wire n_8_0_2618;
   wire n_8_0_2619;
   wire n_8_0_2620;
   wire n_8_0_2621;
   wire n_8_0_2622;
   wire n_8_0_2623;
   wire n_8_0_2624;
   wire n_8_0_2625;
   wire n_8_0_2626;
   wire n_8_0_2627;
   wire n_8_0_2628;
   wire n_8_0_2629;
   wire n_8_0_2630;
   wire n_8_0_2631;
   wire n_8_0_2632;
   wire n_8_0_2633;
   wire n_8_0_2634;
   wire n_8_0_2635;
   wire n_8_0_2636;
   wire n_8_0_2637;
   wire n_8_0_2638;
   wire n_8_0_2639;
   wire n_8_0_2640;
   wire n_8_0_2641;
   wire n_8_0_2642;
   wire n_8_0_2643;
   wire n_8_0_2644;
   wire n_8_0_2645;
   wire n_8_0_2646;
   wire n_8_0_2647;
   wire n_8_0_2648;
   wire n_8_0_2649;
   wire n_8_0_2650;
   wire n_8_0_2651;
   wire n_8_0_2652;
   wire n_8_0_2653;
   wire n_8_0_2654;
   wire n_8_0_2655;
   wire n_8_0_2656;
   wire n_8_0_2657;
   wire n_8_0_2658;
   wire n_8_0_2659;
   wire n_8_0_2660;
   wire n_8_0_2661;
   wire n_8_0_2662;
   wire n_8_0_2663;
   wire n_8_0_2664;
   wire n_8_0_2665;
   wire n_8_0_2666;
   wire n_8_0_2667;
   wire n_8_0_2668;
   wire n_8_0_2669;
   wire n_8_0_2670;
   wire n_8_0_2671;
   wire n_8_0_2672;
   wire n_8_0_2673;
   wire n_8_0_2674;
   wire n_8_0_2675;
   wire n_8_0_2676;
   wire n_8_0_2677;
   wire n_8_0_2678;
   wire n_8_0_2679;
   wire n_8_0_2680;
   wire n_8_0_2681;
   wire n_8_0_2682;
   wire n_8_0_2683;
   wire n_8_0_2684;
   wire n_8_0_2685;
   wire n_8_0_2686;
   wire n_8_0_2687;
   wire n_8_0_2688;
   wire n_8_0_2689;
   wire n_8_0_2690;
   wire n_8_0_2691;
   wire n_8_0_2692;
   wire n_8_0_2693;
   wire n_8_0_2694;
   wire n_8_0_2695;
   wire n_8_0_2696;
   wire n_8_0_2697;
   wire n_8_0_2698;
   wire n_8_0_2699;
   wire n_8_0_2700;
   wire n_8_0_2701;
   wire n_8_0_2702;
   wire n_8_0_2703;
   wire n_8_0_2704;
   wire n_8_0_2705;
   wire n_8_0_2706;
   wire n_8_0_2707;
   wire n_8_0_2708;
   wire n_8_0_2709;
   wire n_8_0_2710;
   wire n_8_0_2711;
   wire n_8_0_2712;
   wire n_8_0_2713;
   wire n_8_0_2714;
   wire n_8_0_2715;
   wire n_8_0_2716;
   wire n_8_0_2717;
   wire n_8_0_2718;
   wire n_8_0_2719;
   wire n_8_0_2720;
   wire n_8_0_2721;
   wire n_8_0_2722;
   wire n_8_0_2723;
   wire n_8_0_2724;
   wire n_8_0_1167;
   wire n_8_0_1168;
   wire n_8_0_2725;
   wire n_8_0_2726;
   wire n_8_0_1169;
   wire n_8_0_1170;
   wire n_8_0_2727;
   wire n_8_0_1171;
   wire n_8_0_2728;
   wire n_8_0_2729;
   wire n_8_0_1172;
   wire n_8_0_1173;
   wire n_8_0_2730;
   wire n_8_0_1174;
   wire n_8_0_1175;
   wire n_8_0_1176;
   wire n_8_0_2731;
   wire n_8_0_1177;
   wire n_8_0_1178;
   wire n_8_0_2732;
   wire n_8_0_1179;
   wire n_8_0_2733;
   wire n_8_0_1180;
   wire n_8_0_1181;
   wire n_8_0_2734;
   wire n_8_0_2735;
   wire n_8_0_1182;
   wire n_8_0_2736;
   wire n_8_0_1183;
   wire n_8_0_2738;
   wire n_8_0_2739;
   wire n_8_0_2740;
   wire n_8_0_1184;
   wire n_8_0_1185;
   wire n_8_0_2741;
   wire n_8_0_2742;
   wire n_8_0_2743;
   wire n_8_0_1186;
   wire n_8_0_1187;
   wire n_8_0_2744;
   wire n_8_0_2745;
   wire n_8_0_2746;
   wire n_8_0_1188;
   wire n_8_0_2747;
   wire n_8_0_2748;
   wire n_8_0_2749;
   wire n_8_0_2750;
   wire n_8_0_1189;
   wire n_8_0_1190;
   wire n_8_0_1191;
   wire n_8_0_2751;
   wire n_8_0_1192;
   wire n_8_0_1193;
   wire n_8_0_2757;
   wire n_8_0_2759;
   wire n_8_0_1194;
   wire n_8_0_1195;
   wire n_8_0_2760;
   wire n_8_0_2762;
   wire n_8_0_2763;
   wire n_8_0_1196;
   wire n_8_0_1197;
   wire n_8_0_2764;
   wire n_8_0_2766;
   wire n_8_0_1198;
   wire n_8_0_2767;
   wire n_8_0_2768;
   wire n_8_0_1199;
   wire n_8_0_1200;
   wire n_8_0_1201;
   wire n_8_0_2769;
   wire n_8_0_2770;
   wire n_8_0_2771;
   wire n_8_0_2772;
   wire n_8_0_2773;
   wire n_8_0_2774;
   wire n_8_0_1202;
   wire n_8_0_1203;
   wire n_8_0_2775;
   wire n_8_0_2776;
   wire n_8_0_2777;
   wire n_8_0_2778;
   wire n_8_0_1204;
   wire n_8_0_2779;
   wire n_8_0_2780;
   wire n_8_0_2781;
   wire n_8_0_2782;
   wire n_8_0_2783;
   wire n_8_0_1205;
   wire n_8_0_1206;
   wire n_8_0_2784;
   wire n_8_0_2785;
   wire n_8_0_2786;
   wire n_8_0_1207;
   wire n_8_0_1208;
   wire n_8_0_2787;
   wire n_8_0_2788;
   wire n_8_0_2789;
   wire n_8_0_2790;
   wire n_8_0_1209;
   wire n_8_0_1210;
   wire n_8_0_2791;
   wire n_8_0_2792;
   wire n_8_0_2793;
   wire n_8_0_2794;
   wire n_8_0_2795;
   wire n_8_0_1211;
   wire n_8_0_1212;
   wire n_8_0_2796;
   wire n_8_0_2797;
   wire n_8_0_2798;
   wire n_8_0_2799;
   wire n_8_0_2800;
   wire n_8_0_2801;
   wire n_8_0_2802;
   wire n_8_0_1213;
   wire n_8_0_2803;
   wire n_8_0_2804;
   wire n_8_0_2805;
   wire n_8_0_2806;
   wire n_8_0_2807;
   wire n_8_0_2808;
   wire n_8_0_2809;
   wire n_8_0_2810;
   wire n_8_0_2811;
   wire n_8_0_1214;
   wire n_8_0_2812;
   wire n_8_0_2813;
   wire n_8_0_2814;
   wire n_8_0_2815;
   wire n_8_0_1215;
   wire n_8_0_1216;
   wire n_8_0_2816;
   wire n_8_0_1217;
   wire n_8_0_1218;
   wire n_8_0_2817;
   wire n_8_0_2818;
   wire n_8_0_2819;
   wire n_8_0_2820;
   wire n_8_0_2821;
   wire n_8_0_2822;
   wire n_8_0_1219;
   wire n_8_0_1220;
   wire n_8_0_1221;
   wire n_8_0_2823;
   wire n_8_0_2824;
   wire n_8_0_2825;
   wire n_8_0_2826;
   wire n_8_0_2827;
   wire n_8_0_2828;
   wire n_8_0_1222;
   wire n_8_0_1223;
   wire n_8_0_1224;
   wire n_8_0_2829;
   wire n_8_0_2830;
   wire n_8_0_2831;
   wire n_8_0_2832;
   wire n_8_0_1225;
   wire n_8_0_1226;
   wire n_8_0_2833;
   wire n_8_0_2834;
   wire n_8_0_1227;
   wire n_8_0_2835;
   wire n_8_0_1228;
   wire n_8_0_2836;
   wire n_8_0_2837;
   wire n_8_0_2838;
   wire n_8_0_2839;
   wire n_8_0_2840;
   wire n_8_0_1229;
   wire n_8_0_1230;
   wire n_8_0_2841;
   wire n_8_0_1231;
   wire n_8_0_2842;
   wire n_8_0_2843;
   wire n_8_0_2844;
   wire n_8_0_1232;
   wire n_8_0_1233;
   wire n_8_0_2845;
   wire n_8_0_2846;
   wire n_8_0_2847;
   wire n_8_0_2848;
   wire n_8_0_2849;
   wire n_8_0_2850;
   wire n_8_0_1234;
   wire n_8_0_1235;
   wire n_8_0_1236;
   wire n_8_0_2851;
   wire n_8_0_2852;
   wire n_8_0_2853;
   wire n_8_0_1237;
   wire n_8_0_1238;
   wire n_8_0_2854;
   wire n_8_0_2855;
   wire n_8_0_2856;
   wire n_8_0_2857;
   wire n_8_0_2858;
   wire n_8_0_2859;
   wire n_8_0_1239;
   wire n_8_0_1240;
   wire n_8_0_2860;
   wire n_8_0_2861;
   wire n_8_0_1241;
   wire n_8_0_2862;
   wire n_8_0_2863;
   wire n_8_0_2864;
   wire n_8_0_2865;
   wire n_8_0_2866;
   wire n_8_0_2867;
   wire n_8_0_1242;
   wire n_8_0_2868;
   wire n_8_0_2869;
   wire n_8_0_1243;
   wire n_8_0_1244;
   wire n_8_0_2870;
   wire n_8_0_2871;
   wire n_8_0_2872;
   wire n_8_0_2873;
   wire n_8_0_1245;
   wire n_8_0_1246;
   wire n_8_0_1247;
   wire n_8_0_2874;
   wire n_8_0_2875;
   wire n_8_0_2876;
   wire n_8_0_2877;
   wire n_8_0_1248;
   wire n_8_0_1249;
   wire n_8_0_1250;
   wire n_8_0_2878;
   wire n_8_0_2879;
   wire n_8_0_2880;
   wire n_8_0_2881;
   wire n_8_0_2882;
   wire n_8_0_2883;
   wire n_8_0_2884;
   wire n_8_0_1251;
   wire n_8_0_2885;
   wire n_8_0_2886;
   wire n_8_0_2887;
   wire n_8_0_2888;
   wire n_8_0_2889;
   wire n_8_0_1252;
   wire n_8_0_2890;
   wire n_8_0_2891;
   wire n_8_0_2892;
   wire n_8_0_1253;
   wire n_8_0_1254;
   wire n_8_0_2893;
   wire n_8_0_1255;
   wire n_8_0_1256;
   wire n_8_0_2894;
   wire n_8_0_2895;
   wire n_8_0_2896;
   wire n_8_0_2897;
   wire n_8_0_2898;
   wire n_8_0_2899;
   wire n_8_0_1257;
   wire n_8_0_1258;
   wire n_8_0_2900;
   wire n_8_0_2901;
   wire n_8_0_2902;
   wire n_8_0_1259;
   wire n_8_0_2903;
   wire n_8_0_1260;
   wire n_8_0_1261;
   wire n_8_0_2904;
   wire n_8_0_2905;
   wire n_8_0_2906;
   wire n_8_0_2907;
   wire n_8_0_2908;
   wire n_8_0_1262;
   wire n_8_0_2909;
   wire n_8_0_2910;
   wire n_8_0_1263;
   wire n_8_0_1264;
   wire n_8_0_2911;
   wire n_8_0_2912;
   wire n_8_0_2913;
   wire n_8_0_2914;
   wire n_8_0_2915;
   wire n_8_0_2916;
   wire n_8_0_1265;
   wire n_8_0_1266;
   wire n_8_0_1267;
   wire n_8_0_2917;
   wire n_8_0_2921;
   wire n_8_0_2922;
   wire n_8_0_1268;
   wire n_8_0_1269;
   wire n_8_0_2923;
   wire n_8_0_2924;
   wire n_8_0_2925;
   wire n_8_0_2926;
   wire n_8_0_1270;
   wire n_8_0_1271;
   wire n_8_0_1272;
   wire n_8_0_1273;
   wire n_8_0_2927;
   wire n_8_0_2929;
   wire n_8_0_2930;
   wire n_8_0_2931;
   wire n_8_0_1274;
   wire n_8_0_1275;
   wire n_8_0_1276;
   wire n_8_0_2932;
   wire n_8_0_2933;
   wire n_8_0_1277;
   wire n_8_0_1278;
   wire n_8_0_2934;
   wire n_8_0_2936;
   wire n_8_0_2937;
   wire n_8_0_1279;
   wire n_8_0_1280;
   wire n_8_0_1281;
   wire n_8_0_2938;
   wire n_8_0_2940;
   wire n_8_0_2941;
   wire n_8_0_2942;
   wire n_8_0_1282;
   wire n_8_0_1283;
   wire n_8_0_1284;
   wire n_8_0_2945;
   wire n_8_0_1285;
   wire n_8_0_1286;
   wire n_8_0_2947;
   wire n_8_0_2948;
   wire n_8_0_2949;
   wire n_8_0_1287;
   wire n_8_0_1288;
   wire n_8_0_2950;
   wire n_8_0_2951;
   wire n_8_0_2952;
   wire n_8_0_2953;
   wire n_8_0_2954;
   wire n_8_0_2955;
   wire n_8_0_2956;
   wire n_8_0_2957;
   wire n_8_0_1289;
   wire n_8_0_2958;
   wire n_8_0_2959;
   wire n_8_0_2960;
   wire n_8_0_2961;
   wire n_8_0_2962;
   wire n_8_0_1290;
   wire n_8_0_2963;
   wire n_8_0_2964;
   wire n_8_0_2965;
   wire n_8_0_1291;
   wire n_8_0_2966;
   wire n_8_0_2967;
   wire n_8_0_2968;
   wire n_8_0_2969;
   wire n_8_0_1292;
   wire n_8_0_2970;
   wire n_8_0_2971;
   wire n_8_0_2972;
   wire n_8_0_2973;
   wire n_8_0_2974;
   wire n_8_0_2975;
   wire n_8_0_1293;
   wire n_8_0_2976;
   wire n_8_0_1294;
   wire n_8_0_2977;
   wire n_8_0_1295;
   wire n_8_0_2978;
   wire n_8_0_1296;
   wire n_8_0_2983;
   wire n_8_0_2984;
   wire n_8_0_2985;
   wire n_8_0_2986;
   wire n_8_0_2987;
   wire n_8_0_1297;
   wire n_8_0_2988;
   wire n_8_0_2993;
   wire n_8_0_1298;
   wire n_8_0_2995;
   wire n_8_0_2996;
   wire n_8_0_1299;
   wire n_8_0_2997;
   wire n_8_0_2999;
   wire n_8_0_1300;
   wire n_8_0_1301;
   wire n_8_0_3000;
   wire n_8_0_3001;
   wire n_8_0_1302;
   wire n_8_0_1303;
   wire n_8_0_3005;
   wire n_8_0_3006;
   wire n_8_0_1304;
   wire n_8_0_3010;
   wire n_8_0_1305;
   wire n_8_0_3012;
   wire n_8_0_1306;
   wire n_8_0_3013;
   wire n_8_0_3015;
   wire n_8_0_3016;
   wire n_8_0_3017;
   wire n_8_0_3018;
   wire n_8_0_1307;
   wire n_8_0_3019;
   wire n_8_0_3020;
   wire n_8_0_3021;
   wire n_8_0_3022;
   wire n_8_0_3023;
   wire n_8_0_3024;
   wire n_8_0_3025;
   wire n_8_0_3026;
   wire n_8_0_3027;
   wire n_8_0_1308;
   wire n_8_0_3028;
   wire n_8_0_3029;
   wire n_8_0_3030;
   wire n_8_0_1309;
   wire n_8_0_3031;
   wire n_8_0_3032;
   wire n_8_0_3033;
   wire n_8_0_3034;
   wire n_8_0_1310;
   wire n_8_0_3035;
   wire n_8_0_3036;
   wire n_8_0_1311;
   wire n_8_0_3037;
   wire n_8_0_3038;
   wire n_8_0_3039;
   wire n_8_0_3040;
   wire n_8_0_1312;
   wire n_8_0_3041;
   wire n_8_0_1313;
   wire n_8_0_3042;
   wire n_8_0_3043;
   wire n_8_0_1314;
   wire n_8_0_3044;
   wire n_8_0_3045;
   wire n_8_0_3046;
   wire n_8_0_3047;
   wire n_8_0_3048;
   wire n_8_0_3049;
   wire n_8_0_3050;
   wire n_8_0_3051;
   wire n_8_0_3052;
   wire n_8_0_1315;
   wire n_8_0_3053;
   wire n_8_0_1316;
   wire n_8_0_3054;
   wire n_8_0_3055;
   wire n_8_0_3056;
   wire n_8_0_3057;
   wire n_8_0_1317;
   wire n_8_0_3058;
   wire n_8_0_3059;
   wire n_8_0_3060;
   wire n_8_0_1318;
   wire n_8_0_3061;
   wire n_8_0_3062;
   wire n_8_0_3063;
   wire n_8_0_1319;
   wire n_8_0_3064;
   wire n_8_0_3065;
   wire n_8_0_3066;
   wire n_8_0_3067;
   wire n_8_0_1320;
   wire n_8_0_3068;
   wire n_8_0_3069;
   wire n_8_0_3070;
   wire n_8_0_3071;
   wire n_8_0_1321;
   wire n_8_0_3072;
   wire n_8_0_3073;
   wire n_8_0_3076;
   wire n_8_0_3077;
   wire n_8_0_3078;
   wire n_8_0_1322;
   wire n_8_0_1323;
   wire n_8_0_3082;
   wire n_8_0_3083;
   wire n_8_0_3084;
   wire n_8_0_1324;
   wire n_8_0_3086;
   wire n_8_0_1325;
   wire n_8_0_1326;
   wire n_8_0_3087;
   wire n_8_0_3088;
   wire n_8_0_3089;
   wire n_8_0_3091;
   wire n_8_0_3092;
   wire n_8_0_1327;
   wire n_8_0_1328;
   wire n_8_0_3093;
   wire n_8_0_3094;
   wire n_8_0_1329;
   wire n_8_0_3096;
   wire n_8_0_1330;
   wire n_8_0_3097;
   wire n_8_0_3101;
   wire n_8_0_1331;
   wire n_8_0_3103;
   wire n_8_0_3104;
   wire n_8_0_1332;
   wire n_8_0_3105;
   wire n_8_0_3106;
   wire n_8_0_3107;
   wire n_8_0_1333;
   wire n_8_0_3108;
   wire n_8_0_3109;
   wire n_8_0_3110;
   wire n_8_0_1334;
   wire n_8_0_3111;
   wire n_8_0_3112;
   wire n_8_0_1335;
   wire n_8_0_3113;
   wire n_8_0_1336;
   wire n_8_0_3118;
   wire n_8_0_3119;
   wire n_8_0_1337;
   wire n_8_0_3120;
   wire n_8_0_3121;
   wire n_8_0_3122;
   wire n_8_0_3125;
   wire n_8_0_3126;
   wire n_8_0_3127;
   wire n_8_0_3129;
   wire n_8_0_3130;
   wire n_8_0_1338;
   wire n_8_0_3131;
   wire n_8_0_3132;
   wire n_8_0_3133;
   wire n_8_0_1339;
   wire n_8_0_3134;
   wire n_8_0_3135;
   wire n_8_0_3136;
   wire n_8_0_1340;
   wire n_8_0_3137;
   wire n_8_0_3138;
   wire n_8_0_1341;
   wire n_8_0_1342;
   wire n_8_0_1343;
   wire n_8_0_3143;
   wire n_8_0_3144;
   wire n_8_0_1344;
   wire n_8_0_3146;
   wire n_8_0_3147;
   wire n_8_0_3148;
   wire n_8_0_3149;
   wire n_8_0_3150;
   wire n_8_0_3151;
   wire n_8_0_3152;
   wire n_8_0_3153;
   wire n_8_0_3154;
   wire n_8_0_1345;
   wire n_8_0_3155;
   wire n_8_0_3156;
   wire n_8_0_3157;
   wire n_8_0_3158;
   wire n_8_0_1346;
   wire n_8_0_3159;
   wire n_8_0_3160;
   wire n_8_0_1347;
   wire n_8_0_3161;
   wire n_8_0_3162;
   wire n_8_0_3163;
   wire n_8_0_3164;
   wire n_8_0_1348;
   wire n_8_0_3165;
   wire n_8_0_3166;
   wire n_8_0_3167;
   wire n_8_0_1349;
   wire n_8_0_1350;
   wire n_8_0_3168;
   wire n_8_0_3169;
   wire n_8_0_3170;
   wire n_8_0_1351;
   wire n_8_0_3171;
   wire n_8_0_3172;
   wire n_8_0_3173;
   wire n_8_0_1352;
   wire n_8_0_3178;
   wire n_8_0_3179;
   wire n_8_0_3180;
   wire n_8_0_3181;
   wire n_8_0_1353;
   wire n_8_0_3182;
   wire n_8_0_3183;
   wire n_8_0_3184;
   wire n_8_0_3185;
   wire n_8_0_3186;
   wire n_8_0_1354;
   wire n_8_0_3188;
   wire n_8_0_3189;
   wire n_8_0_3190;
   wire n_8_0_1355;
   wire n_8_0_3191;
   wire n_8_0_3192;
   wire n_8_0_3193;
   wire n_8_0_3194;
   wire n_8_0_3195;
   wire n_8_0_1356;
   wire n_8_0_3197;
   wire n_8_0_3198;
   wire n_8_0_3199;
   wire n_8_0_1357;
   wire n_8_0_3201;
   wire n_8_0_3202;
   wire n_8_0_3203;
   wire n_8_0_1358;
   wire n_8_0_3204;
   wire n_8_0_3206;
   wire n_8_0_3207;
   wire n_8_0_1359;
   wire n_8_0_3208;
   wire n_8_0_1360;
   wire n_8_0_3216;
   wire n_8_0_3217;
   wire n_8_0_3218;
   wire n_8_0_1361;
   wire n_8_0_3220;
   wire n_8_0_1362;
   wire n_8_0_3221;
   wire n_8_0_3222;
   wire n_8_0_3223;
   wire n_8_0_3224;
   wire n_8_0_3225;
   wire n_8_0_3226;
   wire n_8_0_3227;
   wire n_8_0_3229;
   wire n_8_0_3230;
   wire n_8_0_1363;
   wire n_8_0_3232;
   wire n_8_0_3233;
   wire n_8_0_3234;
   wire n_8_0_1364;
   wire n_8_0_3236;
   wire n_8_0_3237;
   wire n_8_0_1365;
   wire n_8_0_3240;
   wire n_8_0_1366;
   wire n_8_0_3245;
   wire n_8_0_3246;
   wire n_8_0_3247;
   wire n_8_0_3248;
   wire n_8_0_3249;
   wire n_8_0_3250;
   wire n_8_0_3251;
   wire n_8_0_3252;
   wire n_8_0_3253;
   wire n_8_0_3254;
   wire n_8_0_3255;
   wire n_8_0_3256;
   wire n_8_0_3257;
   wire n_8_0_3258;
   wire n_8_0_1367;
   wire n_8_0_1368;
   wire n_8_0_3259;
   wire n_8_0_3260;
   wire n_8_0_3261;
   wire n_8_0_1369;
   wire n_8_0_3262;
   wire n_8_0_3263;
   wire n_8_0_3264;
   wire n_8_0_3265;
   wire n_8_0_1370;
   wire n_8_0_3266;
   wire n_8_0_3267;
   wire n_8_0_3268;
   wire n_8_0_3269;
   wire n_8_0_3270;
   wire n_8_0_3271;
   wire n_8_0_3272;
   wire n_8_0_3273;
   wire n_8_0_3274;
   wire n_8_0_3275;
   wire n_8_0_1371;
   wire n_8_0_3281;
   wire n_8_0_3283;
   wire n_8_0_3284;
   wire n_8_0_3286;
   wire n_8_0_3287;
   wire n_8_0_1372;
   wire n_8_0_3288;
   wire n_8_0_3289;
   wire n_8_0_3290;
   wire n_8_0_3291;
   wire n_8_0_1373;
   wire n_8_0_3292;
   wire n_8_0_3293;
   wire n_8_0_3294;
   wire n_8_0_3295;
   wire n_8_0_1374;
   wire n_8_0_3297;
   wire n_8_0_3299;
   wire n_8_0_3300;
   wire n_8_0_3301;
   wire n_8_0_3304;
   wire n_8_0_3305;
   wire n_8_0_3306;
   wire n_8_0_3307;
   wire n_8_0_3308;
   wire n_8_0_3310;
   wire n_8_0_3311;
   wire n_8_0_3312;
   wire n_8_0_1375;
   wire n_8_0_3313;
   wire n_8_0_3314;
   wire n_8_0_3315;
   wire n_8_0_3316;
   wire n_8_0_3317;
   wire n_8_0_3318;
   wire n_8_0_1376;
   wire n_8_0_1377;
   wire n_8_0_3319;
   wire n_8_0_3320;
   wire n_8_0_3321;
   wire n_8_0_3322;
   wire n_8_0_3323;
   wire n_8_0_3324;
   wire n_8_0_3325;
   wire n_8_0_3326;
   wire n_8_0_3327;
   wire n_8_0_3329;
   wire n_8_0_3331;
   wire n_8_0_3332;
   wire n_8_0_3333;
   wire n_8_0_3334;
   wire n_8_0_3335;
   wire n_8_0_3338;
   wire n_8_0_3339;
   wire n_8_0_3340;
   wire n_8_0_3341;
   wire n_8_0_3342;
   wire n_8_0_3343;
   wire n_8_0_3344;
   wire n_8_0_3345;
   wire n_8_0_1378;
   wire n_8_0_3346;
   wire n_8_0_3347;
   wire n_8_0_3348;
   wire n_8_0_1379;
   wire n_8_0_3349;
   wire n_8_0_3350;
   wire n_8_0_3351;
   wire n_8_0_3353;
   wire n_8_0_3356;
   wire n_8_0_3358;
   wire n_8_0_3359;
   wire n_8_0_3360;
   wire n_8_0_3361;
   wire n_8_0_1380;
   wire n_8_0_3362;
   wire n_8_0_3363;
   wire n_8_0_3364;
   wire n_8_0_3366;
   wire n_8_0_3367;
   wire n_8_0_3368;
   wire n_8_0_3369;
   wire n_8_0_3370;
   wire n_8_0_3371;
   wire n_8_0_3373;
   wire n_8_0_3374;
   wire n_8_0_3378;
   wire n_8_0_3379;
   wire n_8_0_3380;
   wire n_8_0_3381;
   wire n_8_0_3382;
   wire n_8_0_3383;
   wire n_8_0_3384;
   wire n_8_0_3385;
   wire n_8_0_3386;
   wire n_8_0_3387;
   wire n_8_0_1381;
   wire n_8_0_3388;
   wire n_8_0_3389;
   wire n_8_0_3390;
   wire n_8_0_3391;
   wire n_8_0_3392;
   wire n_8_0_3393;
   wire n_8_0_1382;
   wire n_8_0_3394;
   wire n_8_0_3395;
   wire n_8_0_1383;
   wire n_8_0_3396;
   wire n_8_0_3397;
   wire n_8_0_3398;
   wire n_8_0_1384;
   wire n_8_0_3399;
   wire n_8_0_3400;
   wire n_8_0_3401;
   wire n_8_0_3402;
   wire n_8_0_3403;
   wire n_8_0_3404;
   wire n_8_0_3405;
   wire n_8_0_3406;
   wire n_8_0_3407;
   wire n_8_0_3408;
   wire n_8_0_3409;
   wire n_8_0_3410;
   wire n_8_0_3411;
   wire n_8_0_3412;
   wire n_8_0_3413;
   wire n_8_0_3414;
   wire n_8_0_3415;
   wire n_8_0_3416;
   wire n_8_0_3417;
   wire n_8_0_3418;
   wire n_8_0_3419;
   wire n_8_0_3420;
   wire n_8_0_3421;
   wire n_8_0_3422;
   wire n_8_0_3423;
   wire n_8_0_3424;
   wire n_8_0_3425;
   wire n_8_0_3426;
   wire n_8_0_3427;
   wire n_8_0_1385;
   wire n_8_0_3428;
   wire n_8_0_3429;
   wire n_8_0_1386;
   wire n_8_0_3430;
   wire n_8_0_3431;
   wire n_8_0_3432;
   wire n_8_0_1387;
   wire n_8_0_3433;
   wire n_8_0_3434;
   wire n_8_0_3435;
   wire n_8_0_3436;
   wire n_8_0_3437;
   wire n_8_0_3438;
   wire n_8_0_1388;
   wire n_8_0_3439;
   wire n_8_0_3440;
   wire n_8_0_3441;
   wire n_8_0_1389;
   wire n_8_0_3442;
   wire n_8_0_3443;
   wire n_8_0_3444;
   wire n_8_0_1390;
   wire n_8_0_3445;
   wire n_8_0_3446;
   wire n_8_0_3447;
   wire n_8_0_3448;
   wire n_8_0_3449;
   wire n_8_0_3450;
   wire n_8_0_3451;
   wire n_8_0_3452;
   wire n_8_0_3453;
   wire n_8_0_3454;
   wire n_8_0_3455;
   wire n_8_0_3456;
   wire n_8_0_3457;
   wire n_8_0_3458;
   wire n_8_0_1391;
   wire n_8_0_3459;
   wire n_8_0_3462;
   wire n_8_0_3463;
   wire n_8_0_3464;
   wire n_8_0_3465;
   wire n_8_0_3466;
   wire n_8_0_3467;
   wire n_8_0_3469;
   wire n_8_0_3470;
   wire n_8_0_3471;
   wire n_8_0_3472;
   wire n_8_0_3473;
   wire n_8_0_3479;
   wire n_8_0_3480;
   wire n_8_0_3481;
   wire n_8_0_3482;
   wire n_8_0_3483;
   wire n_8_0_1392;
   wire n_8_0_3485;
   wire n_8_0_1393;
   wire n_8_0_3486;
   wire n_8_0_3487;
   wire n_8_0_3488;
   wire n_8_0_3489;
   wire n_8_0_3490;
   wire n_8_0_3491;
   wire n_8_0_3492;
   wire n_8_0_3493;
   wire n_8_0_3494;
   wire n_8_0_3495;
   wire n_8_0_3496;
   wire n_8_0_3497;
   wire n_8_0_3498;
   wire n_8_0_3499;
   wire n_8_0_1394;
   wire n_8_0_3500;
   wire n_8_0_3501;
   wire n_8_0_3502;
   wire n_8_0_3503;
   wire n_8_0_3504;
   wire n_8_0_1395;
   wire n_8_0_3505;
   wire n_8_0_3506;
   wire n_8_0_3507;
   wire n_8_0_3508;
   wire n_8_0_3509;
   wire n_8_0_3510;
   wire n_8_0_1396;
   wire n_8_0_3511;
   wire n_8_0_3512;
   wire n_8_0_1397;
   wire n_8_0_3513;
   wire n_8_0_3514;
   wire n_8_0_3515;
   wire n_8_0_3516;
   wire n_8_0_3517;
   wire n_8_0_3518;
   wire n_8_0_3519;
   wire n_8_0_3520;
   wire n_8_0_3521;
   wire n_8_0_3522;
   wire n_8_0_1398;
   wire n_8_0_3523;
   wire n_8_0_3524;
   wire n_8_0_3525;
   wire n_8_0_3526;
   wire n_8_0_3527;
   wire n_8_0_3528;
   wire n_8_0_3529;
   wire n_8_0_1399;
   wire n_8_0_3530;
   wire n_8_0_3531;
   wire n_8_0_3532;
   wire n_8_0_3533;
   wire n_8_0_1400;
   wire n_8_0_3534;
   wire n_8_0_3535;
   wire n_8_0_3536;
   wire n_8_0_3537;
   wire n_8_0_3538;
   wire n_8_0_1401;
   wire n_8_0_3539;
   wire n_8_0_3540;
   wire n_8_0_3541;
   wire n_8_0_3542;
   wire n_8_0_3543;
   wire n_8_0_3547;
   wire n_8_0_3549;
   wire n_8_0_1402;
   wire n_8_0_3550;
   wire n_8_0_3551;
   wire n_8_0_3552;
   wire n_8_0_3553;
   wire n_8_0_1403;
   wire n_8_0_1404;
   wire n_8_0_3559;
   wire n_8_0_1405;
   wire n_8_0_3560;
   wire n_8_0_3562;
   wire n_8_0_3563;
   wire n_8_0_3564;
   wire n_8_0_3565;
   wire n_8_0_1406;
   wire n_8_0_3567;
   wire n_8_0_3568;
   wire n_8_0_1407;
   wire n_8_0_3571;
   wire n_8_0_3572;
   wire n_8_0_3575;
   wire n_8_0_1408;
   wire n_8_0_3576;
   wire n_8_0_3578;
   wire n_8_0_3579;
   wire n_8_0_1409;
   wire n_8_0_3583;
   wire n_8_0_3584;
   wire n_8_0_3585;
   wire n_8_0_3586;
   wire n_8_0_3588;
   wire n_8_0_3589;
   wire n_8_0_3590;
   wire n_8_0_3592;
   wire n_8_0_3593;
   wire n_8_0_1410;
   wire n_8_0_3595;
   wire n_8_0_3596;
   wire n_8_0_3597;
   wire n_8_0_3598;
   wire n_8_0_1411;
   wire n_8_0_3606;
   wire n_8_0_3607;
   wire n_8_0_3608;
   wire n_8_0_1412;
   wire n_8_0_3609;
   wire n_8_0_3610;
   wire n_8_0_3611;
   wire n_8_0_3612;
   wire n_8_0_3613;
   wire n_8_0_3614;
   wire n_8_0_1413;
   wire n_8_0_3616;
   wire n_8_0_3617;
   wire n_8_0_3618;
   wire n_8_0_3619;
   wire n_8_0_3620;
   wire n_8_0_3621;
   wire n_8_0_3622;
   wire n_8_0_3623;
   wire n_8_0_3625;
   wire n_8_0_3626;
   wire n_8_0_3627;
   wire n_8_0_3628;
   wire n_8_0_3629;
   wire n_8_0_1414;
   wire n_8_0_3630;
   wire n_8_0_3631;
   wire n_8_0_3632;
   wire n_8_0_1415;
   wire n_8_0_3633;
   wire n_8_0_3634;
   wire n_8_0_3635;
   wire n_8_0_3636;
   wire n_8_0_3637;
   wire n_8_0_3638;
   wire n_8_0_3639;
   wire n_8_0_3640;
   wire n_8_0_3641;
   wire n_8_0_3642;
   wire n_8_0_3643;
   wire n_8_0_3644;
   wire n_8_0_3645;
   wire n_8_0_3646;
   wire n_8_0_3647;
   wire n_8_0_3648;
   wire n_8_0_3649;
   wire n_8_0_3650;
   wire n_8_0_3651;
   wire n_8_0_3652;
   wire n_8_0_3653;
   wire n_8_0_3654;
   wire n_8_0_3655;
   wire n_8_0_3656;
   wire n_8_0_3660;
   wire n_8_0_3661;
   wire n_8_0_3662;
   wire n_8_0_3663;
   wire n_8_0_3664;
   wire n_8_0_3665;
   wire n_8_0_3666;
   wire n_8_0_3667;
   wire n_8_0_3668;
   wire n_8_0_3669;
   wire n_8_0_3670;
   wire n_8_0_3671;
   wire n_8_0_3672;
   wire n_8_0_3673;
   wire n_8_0_3674;
   wire n_8_0_3675;
   wire n_8_0_3676;
   wire n_8_0_3677;
   wire n_8_0_3683;
   wire n_8_0_3684;
   wire n_8_0_3685;
   wire n_8_0_3686;
   wire n_8_0_3688;
   wire n_8_0_3693;
   wire n_8_0_3695;
   wire n_8_0_3696;
   wire n_8_0_3697;
   wire n_8_0_3700;
   wire n_8_0_3701;
   wire n_8_0_3703;
   wire n_8_0_3704;
   wire n_8_0_3706;
   wire n_8_0_3707;
   wire n_8_0_3712;
   wire n_8_0_3713;
   wire n_8_0_3714;
   wire n_8_0_3715;
   wire n_8_0_3716;
   wire n_8_0_3717;
   wire n_8_0_3718;
   wire n_8_0_3719;
   wire n_8_0_3720;
   wire n_8_0_3721;
   wire n_8_0_3722;
   wire n_8_0_3723;
   wire n_8_0_3724;
   wire n_8_0_3725;
   wire n_8_0_3726;
   wire n_8_0_3727;
   wire n_8_0_3728;
   wire n_8_0_3729;
   wire n_8_0_3730;
   wire n_8_0_3731;
   wire n_8_0_3732;
   wire n_8_0_3733;
   wire n_8_0_3734;
   wire n_8_0_3735;
   wire n_8_0_3736;
   wire n_8_0_3737;
   wire n_8_0_3738;
   wire n_8_0_3739;
   wire n_8_0_3740;
   wire n_8_0_3741;
   wire n_8_0_3742;
   wire n_8_0_3743;
   wire n_8_0_3744;
   wire n_8_0_3745;
   wire n_8_0_3746;
   wire n_8_0_3747;
   wire n_8_0_3748;
   wire n_8_0_3749;
   wire n_8_0_3750;
   wire n_8_0_3753;
   wire n_8_0_3754;
   wire n_8_0_3760;
   wire n_8_0_3761;
   wire n_8_0_3763;
   wire n_8_0_3764;
   wire n_8_0_3765;
   wire n_8_0_3766;
   wire n_8_0_3767;
   wire n_8_0_3768;
   wire n_8_0_3769;
   wire n_8_0_3770;
   wire n_8_0_3771;
   wire n_8_0_3772;
   wire n_8_0_3773;
   wire n_8_0_3774;
   wire n_8_0_3775;
   wire n_8_0_3776;
   wire n_8_0_3777;
   wire n_8_0_3778;
   wire n_8_0_3779;
   wire n_8_0_3780;
   wire n_8_0_3781;
   wire n_8_0_3782;
   wire n_8_0_3783;
   wire n_8_0_3784;
   wire n_8_0_3785;
   wire n_8_0_3786;
   wire n_8_0_3787;
   wire n_8_0_3788;
   wire n_8_0_3789;
   wire n_8_0_3790;
   wire n_8_0_3791;
   wire n_8_0_3792;
   wire n_8_0_3793;
   wire n_8_0_3794;
   wire n_8_0_3795;
   wire n_8_0_3796;
   wire n_8_0_3797;
   wire n_8_0_3798;
   wire n_8_0_3799;
   wire n_8_0_3800;
   wire n_8_0_3801;
   wire n_8_0_3802;
   wire n_8_0_3803;
   wire n_8_0_3804;
   wire n_8_0_3805;
   wire n_8_0_3806;
   wire n_8_0_3807;
   wire n_8_0_3808;
   wire n_8_0_3809;
   wire n_8_0_3813;
   wire n_8_0_3814;
   wire n_8_0_3815;
   wire n_8_0_3816;
   wire n_8_0_3817;
   wire n_8_0_3818;
   wire n_8_0_3822;
   wire n_8_0_3823;
   wire n_8_0_3824;
   wire n_8_0_3825;
   wire n_8_0_3826;
   wire n_8_0_3827;
   wire n_8_0_3828;
   wire n_8_0_3829;
   wire n_8_0_3830;
   wire n_8_0_3831;
   wire n_8_0_3832;
   wire n_8_0_3833;
   wire n_8_0_3834;
   wire n_8_0_3836;
   wire n_8_0_3837;
   wire n_8_0_3838;
   wire n_8_0_3841;
   wire n_8_0_3842;
   wire n_8_0_3843;
   wire n_8_0_3844;
   wire n_8_0_3845;
   wire n_8_0_3846;
   wire n_8_0_3847;
   wire n_8_0_3848;
   wire n_8_0_3849;
   wire n_8_0_3850;
   wire n_8_0_3851;
   wire n_8_0_3852;
   wire n_8_0_3856;
   wire n_8_0_3857;
   wire n_8_0_3858;
   wire n_8_0_3859;
   wire n_8_0_3860;
   wire n_8_0_3861;
   wire n_8_0_3862;
   wire n_8_0_3864;
   wire n_8_0_3865;
   wire n_8_0_3867;
   wire n_8_0_3868;
   wire n_8_0_3869;
   wire n_8_0_3870;
   wire n_8_0_3871;
   wire n_8_0_3872;
   wire n_8_0_3873;
   wire n_8_0_3874;
   wire n_8_0_3875;
   wire n_8_0_3879;
   wire n_8_0_3880;
   wire n_8_0_3888;
   wire n_8_0_3890;
   wire n_8_0_3891;
   wire n_8_0_3894;
   wire n_8_0_3896;
   wire n_8_0_3897;
   wire n_8_0_3898;
   wire n_8_0_3900;
   wire n_8_0_3901;
   wire n_8_0_3902;
   wire n_8_0_3908;
   wire n_8_0_3909;
   wire n_8_0_3910;
   wire n_8_0_3911;
   wire n_8_0_3912;
   wire n_8_0_3913;
   wire n_8_0_3914;
   wire n_8_0_3915;
   wire n_8_0_3916;
   wire n_8_0_3920;
   wire n_8_0_3921;
   wire n_8_0_3922;
   wire n_8_0_3924;
   wire n_8_0_3925;
   wire n_8_0_3926;
   wire n_8_0_3927;
   wire n_8_0_3929;
   wire n_8_0_3930;
   wire n_8_0_3931;
   wire n_8_0_3932;
   wire n_8_0_3933;
   wire n_8_0_3935;
   wire n_8_0_3936;
   wire n_8_0_3937;
   wire n_8_0_3938;
   wire n_8_0_3942;
   wire n_8_0_3943;
   wire n_8_0_3944;
   wire n_8_0_3945;
   wire n_8_0_3946;
   wire n_8_0_3947;
   wire n_8_0_3948;
   wire n_8_0_3949;
   wire n_8_0_3950;
   wire n_8_0_3951;
   wire n_8_0_3952;
   wire n_8_0_3953;
   wire n_8_0_3954;
   wire n_8_0_3955;
   wire n_8_0_3956;
   wire n_8_0_3957;
   wire n_8_0_3958;
   wire n_8_0_3959;
   wire n_8_0_3960;
   wire n_8_0_3961;
   wire n_8_0_3962;
   wire n_8_0_3963;
   wire n_8_0_3964;
   wire n_8_0_3965;
   wire n_8_0_3966;
   wire n_8_0_3967;
   wire n_8_0_3968;
   wire n_8_0_3969;
   wire n_8_0_3970;
   wire n_8_0_3971;
   wire n_8_0_3972;
   wire n_8_0_3973;
   wire n_8_0_3974;
   wire n_8_0_3975;
   wire n_8_0_3976;
   wire n_8_0_3977;
   wire n_8_0_3978;
   wire n_8_0_3979;
   wire n_8_0_3980;
   wire n_8_0_3981;
   wire n_8_0_3982;
   wire n_8_0_3983;
   wire n_8_0_3984;
   wire n_8_0_3985;
   wire n_8_0_3986;
   wire n_8_0_3987;
   wire n_8_0_3988;
   wire n_8_0_3989;
   wire n_8_0_3990;
   wire n_8_0_3991;
   wire n_8_0_3992;
   wire n_8_0_3993;
   wire n_8_0_3994;
   wire n_8_0_3997;
   wire n_8_0_3999;
   wire n_8_0_4000;
   wire n_8_0_4004;
   wire n_8_0_4005;
   wire n_8_0_4006;
   wire n_8_0_4007;
   wire n_8_0_4008;
   wire n_8_0_4009;
   wire n_8_0_4010;
   wire n_8_0_4011;
   wire n_8_0_4012;
   wire n_8_0_4014;
   wire n_8_0_4015;
   wire n_8_0_4016;
   wire n_8_0_4017;
   wire n_8_0_4018;
   wire n_8_0_4019;
   wire n_8_0_4026;
   wire n_8_0_4027;
   wire n_8_0_4028;
   wire n_8_0_4029;
   wire n_8_0_4030;
   wire n_8_0_4031;
   wire n_8_0_4032;
   wire n_8_0_4034;
   wire n_8_0_4036;
   wire n_8_0_4038;
   wire n_8_0_4039;
   wire n_8_0_4041;
   wire n_8_0_4042;
   wire n_8_0_4044;
   wire n_8_0_4045;
   wire n_8_0_4049;
   wire n_8_0_4054;
   wire n_8_0_4055;
   wire n_8_0_4057;
   wire n_8_0_4058;
   wire n_8_0_4059;
   wire n_8_0_4060;
   wire n_8_0_4061;
   wire n_8_0_4062;
   wire n_8_0_4063;
   wire n_8_0_4064;
   wire n_8_0_4066;
   wire n_8_0_4067;
   wire n_8_0_4068;
   wire n_8_0_4069;
   wire n_8_0_4070;
   wire n_8_0_4071;
   wire n_8_0_4072;
   wire n_8_0_4073;
   wire n_8_0_4074;
   wire n_8_0_4078;
   wire n_8_0_4082;
   wire n_8_0_4084;
   wire n_8_0_4085;
   wire n_8_0_4086;
   wire n_8_0_4087;
   wire n_8_0_4088;
   wire n_8_0_4089;
   wire n_8_0_4091;
   wire n_8_0_4092;
   wire n_8_0_4093;
   wire n_8_0_4094;
   wire n_8_0_4095;
   wire n_8_0_4097;
   wire n_8_0_4098;
   wire n_8_0_4099;
   wire n_8_0_4101;
   wire n_8_0_4102;
   wire n_8_0_4103;
   wire n_8_0_4104;
   wire n_8_0_4105;
   wire n_8_0_4106;
   wire n_8_0_4107;
   wire n_8_0_4108;
   wire n_8_0_4109;
   wire n_8_0_4110;
   wire n_8_0_4111;
   wire n_8_0_4112;
   wire n_8_0_4113;
   wire n_8_0_4114;
   wire n_8_0_4117;
   wire n_8_0_4118;
   wire n_8_0_4119;
   wire n_8_0_4120;
   wire n_8_0_4121;
   wire n_8_0_4122;
   wire n_8_0_4123;
   wire n_8_0_4124;
   wire n_8_0_4125;
   wire n_8_0_4126;
   wire n_8_0_4127;
   wire n_8_0_4128;
   wire n_8_0_4129;
   wire n_8_0_4130;
   wire n_8_0_4131;
   wire n_8_0_4132;
   wire n_8_0_4133;
   wire n_8_0_4134;
   wire n_8_0_4135;
   wire n_8_0_4138;
   wire n_8_0_4139;
   wire n_8_0_4140;
   wire n_8_0_4141;
   wire n_8_0_4142;
   wire n_8_0_4143;
   wire n_8_0_4144;
   wire n_8_0_4145;
   wire n_8_0_4146;
   wire n_8_0_4147;
   wire n_8_0_4148;
   wire n_8_0_4149;
   wire n_8_0_4150;
   wire n_8_0_4151;
   wire n_8_0_4152;
   wire n_8_0_4153;
   wire n_8_0_4154;
   wire n_8_0_4155;
   wire n_8_0_4157;
   wire n_8_0_4158;
   wire n_8_0_4159;
   wire n_8_0_4165;
   wire n_8_0_4166;
   wire n_8_0_4167;
   wire n_8_0_4168;
   wire n_8_0_4169;
   wire n_8_0_4170;
   wire n_8_0_4171;
   wire n_8_0_4172;
   wire n_8_0_4173;
   wire n_8_0_4174;
   wire n_8_0_4175;
   wire n_8_0_4176;
   wire n_8_0_4177;
   wire n_8_0_4179;
   wire n_8_0_4180;
   wire n_8_0_4182;
   wire n_8_0_4183;
   wire n_8_0_4186;
   wire n_8_0_4188;
   wire n_8_0_4189;
   wire n_8_0_4191;
   wire n_8_0_4192;
   wire n_8_0_4193;
   wire n_8_0_4194;
   wire n_8_0_4195;
   wire n_8_0_4196;
   wire n_8_0_4197;
   wire n_8_0_4198;
   wire n_8_0_4199;
   wire n_8_0_4200;
   wire n_8_0_4201;
   wire n_8_0_4202;
   wire n_8_0_4203;
   wire n_8_0_4204;
   wire n_8_0_4205;
   wire n_8_0_4208;
   wire n_8_0_4209;
   wire n_8_0_4210;
   wire n_8_0_4212;
   wire n_8_0_4213;
   wire n_8_0_4214;
   wire n_8_0_4215;
   wire n_8_0_4216;
   wire n_8_0_4217;
   wire n_8_0_4218;
   wire n_8_0_4219;
   wire n_8_0_4220;
   wire n_8_0_4221;
   wire n_8_0_4222;
   wire n_8_0_4223;
   wire n_8_0_4224;
   wire n_8_0_4225;
   wire n_8_0_4226;
   wire n_8_0_4227;
   wire n_8_0_4228;
   wire n_8_0_4229;
   wire n_8_0_4230;
   wire n_8_0_4231;
   wire n_8_0_4232;
   wire n_8_0_4233;
   wire n_8_0_4234;
   wire n_8_0_4235;
   wire n_8_0_4236;
   wire n_8_0_4237;
   wire n_8_0_4238;
   wire n_8_0_4239;
   wire n_8_0_4240;
   wire n_8_0_4241;
   wire n_8_0_4242;
   wire n_8_0_4243;
   wire n_8_0_4244;
   wire n_8_0_4245;
   wire n_8_0_4248;
   wire n_8_0_4249;
   wire n_8_0_4251;
   wire n_8_0_4253;
   wire n_8_0_4254;
   wire n_8_0_4255;
   wire n_8_0_4259;
   wire n_8_0_4261;
   wire n_8_0_4262;
   wire n_8_0_4263;
   wire n_8_0_4264;
   wire n_8_0_4265;
   wire n_8_0_4267;
   wire n_8_0_4268;
   wire n_8_0_4269;
   wire n_8_0_4270;
   wire n_8_0_4271;
   wire n_8_0_4273;
   wire n_8_0_4274;
   wire n_8_0_4278;
   wire n_8_0_4279;
   wire n_8_0_4280;
   wire n_8_0_4281;
   wire n_8_0_4282;
   wire n_8_0_4283;
   wire n_8_0_4284;
   wire n_8_0_4285;
   wire n_8_0_4286;
   wire n_8_0_4287;
   wire n_8_0_4288;
   wire n_8_0_4289;
   wire n_8_0_4293;
   wire n_8_0_4295;
   wire n_8_0_4296;
   wire n_8_0_4297;
   wire n_8_0_4298;
   wire n_8_0_4299;
   wire n_8_0_4300;
   wire n_8_0_4304;
   wire n_8_0_4305;
   wire n_8_0_4306;
   wire n_8_0_4307;
   wire n_8_0_4308;
   wire n_8_0_4309;
   wire n_8_0_4310;
   wire n_8_0_4311;
   wire n_8_0_4313;
   wire n_8_0_4315;
   wire n_8_0_4316;
   wire n_8_0_4317;
   wire n_8_0_4319;
   wire n_8_0_4320;
   wire n_8_0_4321;
   wire n_8_0_4322;
   wire n_8_0_4323;
   wire n_8_0_4324;
   wire n_8_0_4325;
   wire n_8_0_4326;
   wire n_8_0_4327;
   wire n_8_0_4329;
   wire n_8_0_4331;
   wire n_8_0_4335;
   wire n_8_0_4336;
   wire n_8_0_4337;
   wire n_8_0_4338;
   wire n_8_0_4339;
   wire n_8_0_4340;
   wire n_8_0_4341;
   wire n_8_0_4342;
   wire n_8_0_4343;
   wire n_8_0_4344;
   wire n_8_0_4345;
   wire n_8_0_4346;
   wire n_8_0_4347;
   wire n_8_0_4348;
   wire n_8_0_4349;
   wire n_8_0_4350;
   wire n_8_0_4351;
   wire n_8_0_4352;
   wire n_8_0_4353;
   wire n_8_0_4354;
   wire n_8_0_4357;
   wire n_8_0_4358;
   wire n_8_0_4359;
   wire n_8_0_4360;
   wire n_8_0_4361;
   wire n_8_0_4362;
   wire n_8_0_4364;
   wire n_8_0_4365;
   wire n_8_0_4366;
   wire n_8_0_4367;
   wire n_8_0_4368;
   wire n_8_0_4369;
   wire n_8_0_4373;
   wire n_8_0_4374;
   wire n_8_0_4376;
   wire n_8_0_4377;
   wire n_8_0_4378;
   wire n_8_0_4380;
   wire n_8_0_4381;
   wire n_8_0_4382;
   wire n_8_0_4383;
   wire n_8_0_4384;
   wire n_8_0_4385;
   wire n_8_0_4386;
   wire n_8_0_4387;
   wire n_8_0_4389;
   wire n_8_0_4390;
   wire n_8_0_4391;
   wire n_8_0_4392;
   wire n_8_0_4393;
   wire n_8_0_4394;
   wire n_8_0_4395;
   wire n_8_0_4396;
   wire n_8_0_4397;
   wire n_8_0_4398;
   wire n_8_0_4399;
   wire n_8_0_4400;
   wire n_8_0_4401;
   wire n_8_0_4402;
   wire n_8_0_4403;
   wire n_8_0_4405;
   wire n_8_0_4406;
   wire n_8_0_4407;
   wire n_8_0_4411;
   wire n_8_0_4412;
   wire n_8_0_4413;
   wire n_8_0_4414;
   wire n_8_0_4415;
   wire n_8_0_4416;
   wire n_8_0_4417;
   wire n_8_0_4418;
   wire n_8_0_4419;
   wire n_8_0_4420;
   wire n_8_0_4421;
   wire n_8_0_4425;
   wire n_8_0_4426;
   wire n_8_0_4427;
   wire n_8_0_4428;
   wire n_8_0_4429;
   wire n_8_0_4430;
   wire n_8_0_4431;
   wire n_8_0_4432;
   wire n_8_0_4433;
   wire n_8_0_4434;
   wire n_8_0_4435;
   wire n_8_0_4436;
   wire n_8_0_4437;
   wire n_8_0_4438;
   wire n_8_0_4439;
   wire n_8_0_4440;
   wire n_8_0_4441;
   wire n_8_0_4442;
   wire n_8_0_4443;
   wire n_8_0_4445;
   wire n_8_0_4446;
   wire n_8_0_4447;
   wire n_8_0_4448;
   wire n_8_0_4449;
   wire n_8_0_4450;
   wire n_8_0_4451;
   wire n_8_0_4452;
   wire n_8_0_4453;
   wire n_8_0_4454;
   wire n_8_0_4455;
   wire n_8_0_4456;
   wire n_8_0_4457;
   wire n_8_0_4458;
   wire n_8_0_4461;
   wire n_8_0_4462;
   wire n_8_0_4463;
   wire n_8_0_4464;
   wire n_8_0_4466;
   wire n_8_0_4467;
   wire n_8_0_4472;
   wire n_8_0_4473;
   wire n_8_0_4477;
   wire n_8_0_4478;
   wire n_8_0_4479;
   wire n_8_0_4480;
   wire n_8_0_4481;
   wire n_8_0_4482;
   wire n_8_0_4483;
   wire n_8_0_4484;
   wire n_8_0_4485;
   wire n_8_0_4486;
   wire n_8_0_4487;
   wire n_8_0_4488;
   wire n_8_0_4489;
   wire n_8_0_4490;
   wire n_8_0_4491;
   wire n_8_0_4492;
   wire n_8_0_4493;
   wire n_8_0_4494;
   wire n_8_0_4495;
   wire n_8_0_4496;
   wire n_8_0_4497;
   wire n_8_0_4498;
   wire n_8_0_4499;
   wire n_8_0_4505;
   wire n_8_0_4506;
   wire n_8_0_4507;
   wire n_8_0_4508;
   wire n_8_0_4509;
   wire n_8_0_4510;
   wire n_8_0_4511;
   wire n_8_0_4512;
   wire n_8_0_4513;
   wire n_8_0_4515;
   wire n_8_0_4516;
   wire n_8_0_4517;
   wire n_8_0_4518;
   wire n_8_0_4519;
   wire n_8_0_4520;
   wire n_8_0_4521;
   wire n_8_0_4522;
   wire n_8_0_4523;
   wire n_8_0_4524;
   wire n_8_0_4525;
   wire n_8_0_4526;
   wire n_8_0_4527;
   wire n_8_0_4528;
   wire n_8_0_4529;
   wire n_8_0_4530;
   wire n_8_0_4533;
   wire n_8_0_4534;
   wire n_8_0_4535;
   wire n_8_0_4536;
   wire n_8_0_4537;
   wire n_8_0_4538;
   wire n_8_0_4539;
   wire n_8_0_4540;
   wire n_8_0_4541;
   wire n_8_0_4542;
   wire n_8_0_4543;
   wire n_8_0_4544;
   wire n_8_0_4545;
   wire n_8_0_4546;
   wire n_8_0_4547;
   wire n_8_0_4548;
   wire n_8_0_4549;
   wire n_8_0_4550;
   wire n_8_0_4551;
   wire n_8_0_4552;
   wire n_8_0_4553;
   wire n_8_0_4554;
   wire n_8_0_4555;
   wire n_8_0_4556;
   wire n_8_0_4557;
   wire n_8_0_4558;
   wire n_8_0_4559;
   wire n_8_0_4560;
   wire n_8_0_4561;
   wire n_8_0_4562;
   wire n_8_0_4563;
   wire n_8_0_4564;
   wire n_8_0_4565;
   wire n_8_0_4570;
   wire n_8_0_4571;
   wire n_8_0_4572;
   wire n_8_0_4573;
   wire n_8_0_4574;
   wire n_8_0_4575;
   wire n_8_0_4576;
   wire n_8_0_4577;
   wire n_8_0_4578;
   wire n_8_0_4579;
   wire n_8_0_4580;
   wire n_8_0_4581;
   wire n_8_0_4582;
   wire n_8_0_4584;
   wire n_8_0_4585;
   wire n_8_0_4586;
   wire n_8_0_4587;
   wire n_8_0_4588;
   wire n_8_0_4590;
   wire n_8_0_4591;
   wire n_8_0_4592;
   wire n_8_0_4593;
   wire n_8_0_4601;
   wire n_8_0_4602;
   wire n_8_0_4603;
   wire n_8_0_4604;
   wire n_8_0_4605;
   wire n_8_0_4606;
   wire n_8_0_4607;
   wire n_8_0_4608;
   wire n_8_0_4609;
   wire n_8_0_4610;
   wire n_8_0_4611;
   wire n_8_0_4612;
   wire n_8_0_4620;
   wire n_8_0_4621;
   wire n_8_0_4622;
   wire n_8_0_4626;
   wire n_8_0_4627;
   wire n_8_0_4628;
   wire n_8_0_4629;
   wire n_8_0_4630;
   wire n_8_0_4631;
   wire n_8_0_4632;
   wire n_8_0_4633;
   wire n_8_0_4634;
   wire n_8_0_4635;
   wire n_8_0_4636;
   wire n_8_0_4637;
   wire n_8_0_4638;
   wire n_8_0_4639;
   wire n_8_0_4640;
   wire n_8_0_4641;
   wire n_8_0_4642;
   wire n_8_0_4643;
   wire n_8_0_4644;
   wire n_8_0_4645;
   wire n_8_0_4646;
   wire n_8_0_4647;
   wire n_8_0_4648;
   wire n_8_0_4649;
   wire n_8_0_4650;
   wire n_8_0_4651;
   wire n_8_0_4652;
   wire n_8_0_4653;
   wire n_8_0_4654;
   wire n_8_0_4655;
   wire n_8_0_4656;
   wire n_8_0_4657;
   wire n_8_0_4658;
   wire n_8_0_4659;
   wire n_8_0_4660;
   wire n_8_0_4661;
   wire n_8_0_4662;
   wire n_8_0_4663;
   wire n_8_0_4664;
   wire n_8_0_4665;
   wire n_8_0_4666;
   wire n_8_0_4667;
   wire n_8_0_4668;
   wire n_8_0_4669;
   wire n_8_0_4670;
   wire n_8_0_4671;
   wire n_8_0_4672;
   wire n_8_0_4673;
   wire n_8_0_4674;
   wire n_8_0_4675;
   wire n_8_0_4676;
   wire n_8_0_4677;
   wire n_8_0_4678;
   wire n_8_0_4679;
   wire n_8_0_4680;
   wire n_8_0_4681;
   wire n_8_0_4682;
   wire n_8_0_4683;
   wire n_8_0_4684;
   wire n_8_0_4685;
   wire n_8_0_4686;
   wire n_8_0_4687;
   wire n_8_0_4688;
   wire n_8_0_4689;
   wire n_8_0_4690;
   wire n_8_0_4691;
   wire n_8_0_4692;
   wire n_8_0_4693;
   wire n_8_0_4694;
   wire n_8_0_4695;
   wire n_8_0_4696;
   wire n_8_0_4697;
   wire n_8_0_4698;
   wire n_8_0_4699;
   wire n_8_0_4700;
   wire n_8_0_4701;
   wire n_8_0_4702;
   wire n_8_0_4703;
   wire n_8_0_4704;
   wire n_8_0_4705;
   wire n_8_0_4706;
   wire n_8_0_4707;
   wire n_8_0_4708;
   wire n_8_0_4709;
   wire n_8_0_4710;
   wire n_8_0_4711;
   wire n_8_0_4712;
   wire n_8_0_4713;
   wire n_8_0_4714;
   wire n_8_0_4715;
   wire n_8_0_4716;
   wire n_8_0_4717;
   wire n_8_0_4718;
   wire n_8_0_4719;
   wire n_8_0_4720;
   wire n_8_0_4721;
   wire n_8_0_4722;
   wire n_8_0_4723;
   wire n_8_0_4724;
   wire n_8_0_4725;
   wire n_8_0_4726;
   wire n_8_0_4727;
   wire n_8_0_4728;
   wire n_8_0_4729;
   wire n_8_0_4730;
   wire n_8_0_4731;
   wire n_8_0_4732;
   wire n_8_0_4733;
   wire n_8_0_4734;
   wire n_8_0_4735;
   wire n_8_0_4736;
   wire n_8_0_4737;
   wire n_8_0_4738;
   wire n_8_0_4739;
   wire n_8_0_4740;
   wire n_8_0_4741;
   wire n_8_0_4742;
   wire n_8_0_4743;
   wire n_8_0_4744;
   wire n_8_0_4745;
   wire n_8_0_4746;
   wire n_8_0_4747;
   wire n_8_0_4748;
   wire n_8_0_4749;
   wire n_8_0_4750;
   wire n_8_0_4751;
   wire n_8_0_4752;
   wire n_8_0_4753;
   wire n_8_0_4754;
   wire n_8_0_4755;
   wire n_8_0_4756;
   wire n_8_0_4757;
   wire n_8_0_4758;
   wire n_8_0_4759;
   wire n_8_0_4760;
   wire n_8_0_4761;
   wire n_8_0_4762;
   wire n_8_0_4763;
   wire n_8_0_4764;
   wire n_8_0_4765;
   wire n_8_0_4766;
   wire n_8_0_4767;
   wire n_8_0_4768;
   wire n_8_0_4769;
   wire n_8_0_4770;
   wire n_8_0_4771;
   wire n_8_0_4772;
   wire n_8_0_4773;
   wire n_8_0_4774;
   wire n_8_0_4775;
   wire n_8_0_4776;
   wire n_8_0_4777;
   wire n_8_0_4778;
   wire n_8_0_4779;
   wire n_8_0_4780;
   wire n_8_0_4781;
   wire n_8_0_4782;
   wire n_8_0_4783;
   wire n_8_0_4784;
   wire n_8_0_4785;
   wire n_8_0_4786;
   wire n_8_0_4787;
   wire n_8_0_4788;
   wire n_8_0_4789;
   wire n_8_0_4790;
   wire n_8_0_4791;
   wire n_8_0_4792;
   wire n_8_0_4793;
   wire n_8_0_4794;
   wire n_8_0_4795;
   wire n_8_0_4796;
   wire n_8_0_4797;
   wire n_8_0_4798;
   wire n_8_0_4799;
   wire n_8_0_4800;
   wire n_8_0_4801;
   wire n_8_0_4802;
   wire n_8_0_4803;
   wire n_8_0_4804;
   wire n_8_0_4805;
   wire n_8_0_4806;
   wire n_8_0_4807;
   wire n_8_0_4808;
   wire n_8_0_4809;
   wire n_8_0_4810;
   wire n_8_0_4811;
   wire n_8_0_4812;
   wire n_8_0_4813;
   wire n_8_0_4817;
   wire n_8_0_4818;
   wire n_8_0_4819;
   wire n_8_0_4825;
   wire n_8_0_4826;
   wire n_8_0_4828;
   wire n_8_0_4829;
   wire n_8_0_4831;
   wire n_8_0_4832;
   wire n_8_0_4833;
   wire n_8_0_4834;
   wire n_8_0_4835;
   wire n_8_0_4836;
   wire n_8_0_4837;
   wire n_8_0_4838;
   wire n_8_0_4839;
   wire n_8_0_4840;
   wire n_8_0_4841;
   wire n_8_0_4842;
   wire n_8_0_4843;
   wire n_8_0_4852;
   wire n_8_0_4853;
   wire n_8_0_4854;
   wire n_8_0_4855;
   wire n_8_0_4856;
   wire n_8_0_4857;
   wire n_8_0_4858;
   wire n_8_0_4859;
   wire n_8_0_4860;
   wire n_8_0_4862;
   wire n_8_0_4863;
   wire n_8_0_4865;
   wire n_8_0_4866;
   wire n_8_0_4868;
   wire n_8_0_4869;
   wire n_8_0_4870;
   wire n_8_0_4871;
   wire n_8_0_4872;
   wire n_8_0_4873;
   wire n_8_0_4874;
   wire n_8_0_4875;
   wire n_8_0_4876;
   wire n_8_0_4877;
   wire n_8_0_4878;
   wire n_8_0_4879;
   wire n_8_0_4880;
   wire n_8_0_4881;
   wire n_8_0_4882;
   wire n_8_0_4883;
   wire n_8_0_4884;
   wire n_8_0_4885;
   wire n_8_0_4886;
   wire n_8_0_4887;
   wire n_8_0_4888;
   wire n_8_0_4889;
   wire n_8_0_4890;
   wire n_8_0_4891;
   wire n_8_0_4892;
   wire n_8_0_4893;
   wire n_8_0_4894;
   wire n_8_0_4895;
   wire n_8_0_4896;
   wire n_8_0_4897;
   wire n_8_0_4898;
   wire n_8_0_4899;
   wire n_8_0_4900;
   wire n_8_0_4901;
   wire n_8_0_4902;
   wire n_8_0_4903;
   wire n_8_0_4904;
   wire n_8_0_4905;
   wire n_8_0_4906;
   wire n_8_0_4907;
   wire n_8_0_4908;
   wire n_8_0_4909;
   wire n_8_0_4910;
   wire n_8_0_4911;
   wire n_8_0_4912;
   wire n_8_0_4913;
   wire n_8_0_4914;
   wire n_8_0_4915;
   wire n_8_0_4916;
   wire n_8_0_4917;
   wire n_8_0_4918;
   wire n_8_0_4919;
   wire n_8_0_4920;
   wire n_8_0_4921;
   wire n_8_0_4922;
   wire n_8_0_4923;
   wire n_8_0_4924;
   wire n_8_0_4925;
   wire n_8_0_4926;
   wire n_8_0_4927;
   wire n_8_0_4928;
   wire n_8_0_4929;
   wire n_8_0_4930;
   wire n_8_0_4931;
   wire n_8_0_4932;
   wire n_8_0_4933;
   wire n_8_0_4934;
   wire n_8_0_4935;
   wire n_8_0_4936;
   wire n_8_0_4937;
   wire n_8_0_4938;
   wire n_8_0_4939;
   wire n_8_0_4940;
   wire n_8_0_4941;
   wire n_8_0_4942;
   wire n_8_0_4943;
   wire n_8_0_4944;
   wire n_8_0_4945;
   wire n_8_0_4946;
   wire n_8_0_4947;
   wire n_8_0_4948;
   wire n_8_0_4949;
   wire n_8_0_4950;
   wire n_8_0_4951;
   wire n_8_0_4952;
   wire n_8_0_4953;
   wire n_8_0_4954;
   wire n_8_0_4955;
   wire n_8_0_4956;
   wire n_8_0_4957;
   wire n_8_0_4958;
   wire n_8_0_4959;
   wire n_8_0_4960;
   wire n_8_0_4961;
   wire n_8_0_4962;
   wire n_8_0_4963;
   wire n_8_0_4964;
   wire n_8_0_4965;
   wire n_8_0_4966;
   wire n_8_0_4967;
   wire n_8_0_4968;
   wire n_8_0_4969;
   wire n_8_0_4970;
   wire n_8_0_4971;
   wire n_8_0_4972;
   wire n_8_0_4973;
   wire n_8_0_4974;
   wire n_8_0_4975;
   wire n_8_0_4976;
   wire n_8_0_4977;
   wire n_8_0_4978;
   wire n_8_0_4979;
   wire n_8_0_4980;
   wire n_8_0_4981;
   wire n_8_0_4982;
   wire n_8_0_4983;
   wire n_8_0_4984;
   wire n_8_0_4985;
   wire n_8_0_4986;
   wire n_8_0_4987;
   wire n_8_0_4988;
   wire n_8_0_4989;
   wire n_8_0_4990;
   wire n_8_0_4991;
   wire n_8_0_4992;
   wire n_8_0_4993;
   wire n_8_0_4994;
   wire n_8_0_4995;
   wire n_8_0_4996;
   wire n_8_0_4997;
   wire n_8_0_4998;
   wire n_8_0_4999;
   wire n_8_0_5000;
   wire n_8_0_5001;
   wire n_8_0_5002;
   wire n_8_0_5003;
   wire n_8_0_5004;
   wire n_8_0_5005;
   wire n_8_0_5006;
   wire n_8_0_5007;
   wire n_8_0_5008;
   wire n_8_0_5009;
   wire n_8_0_5010;
   wire n_8_0_5011;
   wire n_8_0_5012;
   wire n_8_0_5013;
   wire n_8_0_5014;
   wire n_8_0_5015;
   wire n_8_0_5016;
   wire n_8_0_5017;
   wire n_8_0_5018;
   wire n_8_0_5019;
   wire n_8_0_5020;
   wire n_8_0_5021;
   wire n_8_0_5022;
   wire n_8_0_5023;
   wire n_8_0_5024;
   wire n_8_0_5025;
   wire n_8_0_5026;
   wire n_8_0_5027;
   wire n_8_0_5028;
   wire n_8_0_5029;
   wire n_8_0_5030;
   wire n_8_0_5031;
   wire n_8_0_5032;
   wire n_8_0_5033;
   wire n_8_0_5034;
   wire n_8_0_5035;
   wire n_8_0_5036;
   wire n_8_0_5037;
   wire n_8_0_5038;
   wire n_8_0_5039;
   wire n_8_0_5040;
   wire n_8_0_5041;
   wire n_8_0_5042;
   wire n_8_0_5043;
   wire n_8_0_5044;
   wire n_8_0_5045;
   wire n_8_0_5046;
   wire n_8_0_5047;
   wire n_8_0_5048;
   wire n_8_0_5049;
   wire n_8_0_5050;
   wire n_8_0_5051;
   wire n_8_0_5052;
   wire n_8_0_5053;
   wire n_8_0_5054;
   wire n_8_0_5055;
   wire n_8_0_5057;
   wire n_8_0_5058;
   wire n_8_0_5066;
   wire n_8_0_5067;
   wire n_8_0_5069;
   wire n_8_0_5070;
   wire n_8_0_5072;
   wire n_8_0_5073;
   wire n_8_0_5075;
   wire n_8_0_5076;
   wire n_8_0_5078;
   wire n_8_0_5079;
   wire n_8_0_5080;
   wire n_8_0_5083;
   wire n_8_0_5084;
   wire n_8_0_5085;
   wire n_8_0_5086;
   wire n_8_0_5087;
   wire n_8_0_5088;
   wire n_8_0_5089;
   wire n_8_0_5090;
   wire n_8_0_5091;
   wire n_8_0_5092;
   wire n_8_0_5093;
   wire n_8_0_5094;
   wire n_8_0_5095;
   wire n_8_0_5096;
   wire n_8_0_5097;
   wire n_8_0_5098;
   wire n_8_0_5099;
   wire n_8_0_5100;
   wire n_8_0_5101;
   wire n_8_0_5102;
   wire n_8_0_5103;
   wire n_8_0_5104;
   wire n_8_0_5105;
   wire n_8_0_5106;
   wire n_8_0_5107;
   wire n_8_0_5108;
   wire n_8_0_5109;
   wire n_8_0_5110;
   wire n_8_0_5111;
   wire n_8_0_5112;
   wire n_8_0_5113;
   wire n_8_0_5114;
   wire n_8_0_5115;
   wire n_8_0_5116;
   wire n_8_0_5117;
   wire n_8_0_5118;
   wire n_8_0_5119;
   wire n_8_0_5120;
   wire n_8_0_5121;
   wire n_8_0_5122;
   wire n_8_0_5123;
   wire n_8_0_5124;
   wire n_8_0_5125;
   wire n_8_0_5126;
   wire n_8_0_5127;
   wire n_8_0_5128;
   wire n_8_0_5129;
   wire n_8_0_5130;
   wire n_8_0_5131;
   wire n_8_0_5132;
   wire n_8_0_5133;
   wire n_8_0_5134;
   wire n_8_0_5135;
   wire n_8_0_5136;
   wire n_8_0_5137;
   wire n_8_0_5138;
   wire n_8_0_5139;
   wire n_8_0_5140;
   wire n_8_0_5141;
   wire n_8_0_5142;
   wire n_8_0_5143;
   wire n_8_0_5144;
   wire n_8_0_5145;
   wire n_8_0_5146;
   wire n_8_0_5147;
   wire n_8_0_5148;
   wire n_8_0_5149;
   wire n_8_0_5150;
   wire n_8_0_5151;
   wire n_8_0_5152;
   wire n_8_0_5153;
   wire n_8_0_5154;
   wire n_8_0_5155;
   wire n_8_0_5156;
   wire n_8_0_5157;
   wire n_8_0_5158;
   wire n_8_0_5159;
   wire n_8_0_5160;
   wire n_8_0_5161;
   wire n_8_0_5162;
   wire n_8_0_5163;
   wire n_8_0_5164;
   wire n_8_0_5165;
   wire n_8_0_5166;
   wire n_8_0_5167;
   wire n_8_0_5168;
   wire n_8_0_5169;
   wire n_8_0_5170;
   wire n_8_0_5177;
   wire n_8_0_5179;
   wire n_8_0_5180;
   wire n_8_0_5181;
   wire n_8_0_5183;
   wire n_8_0_5184;
   wire n_8_0_5185;
   wire n_8_0_5187;
   wire n_8_0_5189;
   wire n_8_0_5190;
   wire n_8_0_5191;
   wire n_8_0_5194;
   wire n_8_0_5196;
   wire n_8_0_5197;
   wire n_8_0_5198;
   wire n_8_0_5199;
   wire n_8_0_5200;
   wire n_8_0_5201;
   wire n_8_0_5202;
   wire n_8_0_5203;
   wire n_8_0_5204;
   wire n_8_0_5205;
   wire n_8_0_5206;
   wire n_8_0_5207;
   wire n_8_0_5208;
   wire n_8_0_5209;
   wire n_8_0_5210;
   wire n_8_0_5211;
   wire n_8_0_5212;
   wire n_8_0_5213;
   wire n_8_0_5214;
   wire n_8_0_5215;
   wire n_8_0_5216;
   wire n_8_0_5217;
   wire n_8_0_5218;
   wire n_8_0_5219;
   wire n_8_0_5220;
   wire n_8_0_5221;
   wire n_8_0_5222;
   wire n_8_0_5223;
   wire n_8_0_5224;
   wire n_8_0_5225;
   wire n_8_0_5226;
   wire n_8_0_5227;
   wire n_8_0_5228;
   wire n_8_0_5229;
   wire n_8_0_5230;
   wire n_8_0_5231;
   wire n_8_0_5232;
   wire n_8_0_5233;
   wire n_8_0_5234;
   wire n_8_0_5235;
   wire n_8_0_5236;
   wire n_8_0_5237;
   wire n_8_0_5238;
   wire n_8_0_5239;
   wire n_8_0_5240;
   wire n_8_0_5241;
   wire n_8_0_5242;
   wire n_8_0_5243;
   wire n_8_0_5244;
   wire n_8_0_5245;
   wire n_8_0_5246;
   wire n_8_0_5247;
   wire n_8_0_5248;
   wire n_8_0_5249;
   wire n_8_0_5250;
   wire n_8_0_5251;
   wire n_8_0_5252;
   wire n_8_0_5253;
   wire n_8_0_5254;
   wire n_8_0_5255;
   wire n_8_0_5256;
   wire n_8_0_5257;
   wire n_8_0_5258;
   wire n_8_0_5259;
   wire n_8_0_5260;
   wire n_8_0_5261;
   wire n_8_0_5262;
   wire n_8_0_5263;
   wire n_8_0_5264;
   wire n_8_0_5265;
   wire n_8_0_5266;
   wire n_8_0_5267;
   wire n_8_0_5268;
   wire n_8_0_5269;
   wire n_8_0_5270;
   wire n_8_0_5271;
   wire n_8_0_5272;
   wire n_8_0_5273;
   wire n_8_0_5274;
   wire n_8_0_5275;
   wire n_8_0_5276;
   wire n_8_0_5277;
   wire n_8_0_5278;
   wire n_8_0_5279;
   wire n_8_0_5280;
   wire n_8_0_5281;
   wire n_8_0_5282;
   wire n_8_0_5283;
   wire n_8_0_5284;
   wire n_8_0_5285;
   wire n_8_0_5286;
   wire n_8_0_5287;
   wire n_8_0_5288;
   wire n_8_0_5289;
   wire n_8_0_5290;
   wire n_8_0_5291;
   wire n_8_0_5292;
   wire n_8_0_5293;
   wire n_8_0_5294;
   wire n_8_0_5295;
   wire n_8_0_5296;
   wire n_8_0_5297;
   wire n_8_0_5298;
   wire n_8_0_5299;
   wire n_8_0_5300;
   wire n_8_0_5301;
   wire n_8_0_5302;
   wire n_8_0_5303;
   wire n_8_0_5304;
   wire n_8_0_5305;
   wire n_8_0_5306;
   wire n_8_0_5307;
   wire n_8_0_5308;
   wire n_8_0_5309;
   wire n_8_0_5310;
   wire n_8_0_5311;
   wire n_8_0_5312;
   wire n_8_0_5313;
   wire n_8_0_5314;
   wire n_8_0_5315;
   wire n_8_0_5316;
   wire n_8_0_5317;
   wire n_8_0_5318;
   wire n_8_0_5319;
   wire n_8_0_5320;
   wire n_8_0_5321;
   wire n_8_0_5322;
   wire n_8_0_5323;
   wire n_8_0_5324;
   wire n_8_0_5325;
   wire n_8_0_5326;
   wire n_8_0_5327;
   wire n_8_0_5328;
   wire n_8_0_5329;
   wire n_8_0_5330;
   wire n_8_0_5331;
   wire n_8_0_5332;
   wire n_8_0_5333;
   wire n_8_0_5334;
   wire n_8_0_5335;
   wire n_8_0_5336;
   wire n_8_0_5337;
   wire n_8_0_5338;
   wire n_8_0_5339;
   wire n_8_0_5340;
   wire n_8_0_5341;
   wire n_8_0_5342;
   wire n_8_0_5343;
   wire n_8_0_5344;
   wire n_8_0_5345;
   wire n_8_0_5346;
   wire n_8_0_5347;
   wire n_8_0_5348;
   wire n_8_0_5349;
   wire n_8_0_5350;
   wire n_8_0_5351;
   wire n_8_0_5352;
   wire n_8_0_5353;
   wire n_8_0_5354;
   wire n_8_0_5355;
   wire n_8_0_5360;
   wire n_8_0_5363;
   wire n_8_0_5364;
   wire n_8_0_5366;
   wire n_8_0_5367;
   wire n_8_0_5368;
   wire n_8_0_5369;
   wire n_8_0_5370;
   wire n_8_0_5372;
   wire n_8_0_5373;
   wire n_8_0_5375;
   wire n_8_0_5376;
   wire n_8_0_5378;
   wire n_8_0_5379;
   wire n_8_0_5382;
   wire n_8_0_5383;
   wire n_8_0_5384;
   wire n_8_0_5385;
   wire n_8_0_5386;
   wire n_8_0_5387;
   wire n_8_0_5389;
   wire n_8_0_5390;
   wire n_8_0_5393;
   wire n_8_0_5394;
   wire n_8_0_5395;
   wire n_8_0_5396;
   wire n_8_0_5397;
   wire n_8_0_5399;
   wire n_8_0_5400;
   wire n_8_0_5406;
   wire n_8_0_5408;
   wire n_8_0_5409;
   wire n_8_0_5415;
   wire n_8_0_5417;
   wire n_8_0_5418;
   wire n_8_0_5419;
   wire n_8_0_5421;
   wire n_8_0_5422;
   wire n_8_0_5424;
   wire n_8_0_5425;
   wire n_8_0_5426;
   wire n_8_0_5427;
   wire n_8_0_5428;
   wire n_8_0_5429;
   wire n_8_0_5431;
   wire n_8_0_5432;
   wire n_8_0_5433;
   wire n_8_0_5434;
   wire n_8_0_5435;
   wire n_8_0_5439;
   wire n_8_0_5440;
   wire n_8_0_5441;
   wire n_8_0_5442;
   wire n_8_0_5443;
   wire n_8_0_5444;
   wire n_8_0_5445;
   wire n_8_0_5446;
   wire n_8_0_5447;
   wire n_8_0_5448;
   wire n_8_0_5449;
   wire n_8_0_5450;
   wire n_8_0_5451;
   wire n_8_0_5452;
   wire n_8_0_5453;
   wire n_8_0_5454;
   wire n_8_0_5455;
   wire n_8_0_5456;
   wire n_8_0_5457;
   wire n_8_0_5458;
   wire n_8_0_5459;
   wire n_8_0_5460;
   wire n_8_0_5461;
   wire n_8_0_5462;
   wire n_8_0_5463;
   wire n_8_0_5464;
   wire n_8_0_5465;
   wire n_8_0_5466;
   wire n_8_0_5467;
   wire n_8_0_5468;
   wire n_8_0_5469;
   wire n_8_0_5470;
   wire n_8_0_5471;
   wire n_8_0_5472;
   wire n_8_0_5473;
   wire n_8_0_5474;
   wire n_8_0_5475;
   wire n_8_0_5476;
   wire n_8_0_5477;
   wire n_8_0_5478;
   wire n_8_0_5479;
   wire n_8_0_5481;
   wire n_8_0_5482;
   wire n_8_0_5483;
   wire n_8_0_5484;
   wire n_8_0_5485;
   wire n_8_0_5486;
   wire n_8_0_5487;
   wire n_8_0_5488;
   wire n_8_0_5489;
   wire n_8_0_5490;
   wire n_8_0_5491;
   wire n_8_0_5492;
   wire n_8_0_5493;
   wire n_8_0_5494;
   wire n_8_0_5495;
   wire n_8_0_5496;
   wire n_8_0_5497;
   wire n_8_0_5498;
   wire n_8_0_5499;
   wire n_8_0_5500;
   wire n_8_0_5501;
   wire n_8_0_5502;
   wire n_8_0_5503;
   wire n_8_0_5504;
   wire n_8_0_5505;
   wire n_8_0_5506;
   wire n_8_0_5507;
   wire n_8_0_5508;
   wire n_8_0_5509;
   wire n_8_0_5510;
   wire n_8_0_5511;
   wire n_8_0_5512;
   wire n_8_0_5513;
   wire n_8_0_5514;
   wire n_8_0_5515;
   wire n_8_0_5516;
   wire n_8_0_5517;
   wire n_8_0_5518;
   wire n_8_0_5519;
   wire n_8_0_5520;
   wire n_8_0_5521;
   wire n_8_0_5522;
   wire n_8_0_5523;
   wire n_8_0_5524;
   wire n_8_0_5525;
   wire n_8_0_5526;
   wire n_8_0_5527;
   wire n_8_0_5528;
   wire n_8_0_5529;
   wire n_8_0_5530;
   wire n_8_0_5531;
   wire n_8_0_5532;
   wire n_8_0_5533;
   wire n_8_0_5534;
   wire n_8_0_5535;
   wire n_8_0_5536;
   wire n_8_0_5537;
   wire n_8_0_5538;
   wire n_8_0_5539;
   wire n_8_0_5540;
   wire n_8_0_5541;
   wire n_8_0_5542;
   wire n_8_0_5543;
   wire n_8_0_5544;
   wire n_8_0_5545;
   wire n_8_0_5546;
   wire n_8_0_5547;
   wire n_8_0_5548;
   wire n_8_0_5549;
   wire n_8_0_5550;
   wire n_8_0_5551;
   wire n_8_0_5552;
   wire n_8_0_5553;
   wire n_8_0_5554;
   wire n_8_0_5555;
   wire n_8_0_5556;
   wire n_8_0_5557;
   wire n_8_0_5558;
   wire n_8_0_5559;
   wire n_8_0_5560;
   wire n_8_0_5561;
   wire n_8_0_5562;
   wire n_8_0_5563;
   wire n_8_0_5564;
   wire n_8_0_5565;
   wire n_8_0_5566;
   wire n_8_0_5567;
   wire n_8_0_5568;
   wire n_8_0_5569;
   wire n_8_0_5570;
   wire n_8_0_5571;
   wire n_8_0_5572;
   wire n_8_0_5573;
   wire n_8_0_5574;
   wire n_8_0_5575;
   wire n_8_0_5576;
   wire n_8_0_5577;
   wire n_8_0_5578;
   wire n_8_0_5579;
   wire n_8_0_5580;
   wire n_8_0_5581;
   wire n_8_0_5582;
   wire n_8_0_5583;
   wire n_8_0_5584;
   wire n_8_0_5585;
   wire n_8_0_5586;
   wire n_8_0_5587;
   wire n_8_0_5588;
   wire n_8_0_5589;
   wire n_8_0_5590;
   wire n_8_0_5591;
   wire n_8_0_5592;
   wire n_8_0_5593;
   wire n_8_0_5595;
   wire n_8_0_5596;
   wire n_8_0_5597;
   wire n_8_0_5598;
   wire n_8_0_5599;
   wire n_8_0_5600;
   wire n_8_0_5601;
   wire n_8_0_5602;
   wire n_8_0_5603;
   wire n_8_0_5604;
   wire n_8_0_5605;
   wire n_8_0_5606;
   wire n_8_0_5607;
   wire n_8_0_5608;
   wire n_8_0_5609;
   wire n_8_0_5610;
   wire n_8_0_5611;
   wire n_8_0_5612;
   wire n_8_0_5613;
   wire n_8_0_5614;
   wire n_8_0_5615;
   wire n_8_0_5616;
   wire n_8_0_5617;
   wire n_8_0_5618;
   wire n_8_0_5619;
   wire n_8_0_5620;
   wire n_8_0_5621;
   wire n_8_0_5622;
   wire n_8_0_5623;
   wire n_8_0_5624;
   wire n_8_0_5625;
   wire n_8_0_5626;
   wire n_8_0_5627;
   wire n_8_0_5628;
   wire n_8_0_5629;
   wire n_8_0_5630;
   wire n_8_0_5631;
   wire n_8_0_5632;
   wire n_8_0_5633;
   wire n_8_0_5634;
   wire n_8_0_5635;
   wire n_8_0_5636;
   wire n_8_0_5637;
   wire n_8_0_5638;
   wire n_8_0_5639;
   wire n_8_0_5640;
   wire n_8_0_5641;
   wire n_8_0_5642;
   wire n_8_0_5643;
   wire n_8_0_5644;
   wire n_8_0_5645;
   wire n_8_0_5646;
   wire n_8_0_5647;
   wire n_8_0_5648;
   wire n_8_0_5649;
   wire n_8_0_5650;
   wire n_8_0_5651;
   wire n_8_0_5653;
   wire n_8_0_5654;
   wire n_8_0_5655;
   wire n_8_0_5656;
   wire n_8_0_5657;
   wire n_8_0_5658;
   wire n_8_0_5659;
   wire n_8_0_5660;
   wire n_8_0_5661;
   wire n_8_0_5662;
   wire n_8_0_5663;
   wire n_8_0_5664;
   wire n_8_0_5665;
   wire n_8_0_5666;
   wire n_8_0_5667;
   wire n_8_0_5668;
   wire n_8_0_5669;
   wire n_8_0_5670;
   wire n_8_0_5671;
   wire n_8_0_5672;
   wire n_8_0_5673;
   wire n_8_0_5675;
   wire n_8_0_5676;
   wire n_8_0_5677;
   wire n_8_0_5678;
   wire n_8_0_5679;
   wire n_8_0_5680;
   wire n_8_0_5681;
   wire n_8_0_5682;
   wire n_8_0_5683;
   wire n_8_0_5684;
   wire n_8_0_5685;
   wire n_8_0_5686;
   wire n_8_0_5687;
   wire n_8_0_5688;
   wire n_8_0_5689;
   wire n_8_0_5690;
   wire n_8_0_5691;
   wire n_8_0_5692;
   wire n_8_0_5693;
   wire n_8_0_5694;
   wire n_8_0_5695;
   wire n_8_0_5696;
   wire n_8_0_5697;
   wire n_8_0_5698;
   wire n_8_0_5699;
   wire n_8_0_5700;
   wire n_8_0_5701;
   wire n_8_0_5702;
   wire n_8_0_5703;
   wire n_8_0_5704;
   wire n_8_0_5705;
   wire n_8_0_5706;
   wire n_8_0_5707;
   wire n_8_0_5708;
   wire n_8_0_5709;
   wire n_8_0_5710;
   wire n_8_0_5711;
   wire n_8_0_5712;
   wire n_8_0_5713;
   wire n_8_0_5714;
   wire n_8_0_5715;
   wire n_8_0_5716;
   wire n_8_0_5717;
   wire n_8_0_5718;
   wire n_8_0_5719;
   wire n_8_0_5720;
   wire n_8_0_5721;
   wire n_8_0_5722;
   wire n_8_0_5723;
   wire n_8_0_5725;
   wire n_8_0_5726;
   wire n_8_0_5727;
   wire n_8_0_5728;
   wire n_8_0_5729;
   wire n_8_0_5730;
   wire n_8_0_5731;
   wire n_8_0_5732;
   wire n_8_0_5733;
   wire n_8_0_5734;
   wire n_8_0_5735;
   wire n_8_0_5736;
   wire n_8_0_5737;
   wire n_8_0_5738;
   wire n_8_0_5739;
   wire n_8_0_5740;
   wire n_8_0_5741;
   wire n_8_0_5742;
   wire n_8_0_5743;
   wire n_8_0_5744;
   wire n_8_0_5745;
   wire n_8_0_5746;
   wire n_8_0_5747;
   wire n_8_0_5748;
   wire n_8_0_5749;
   wire n_8_0_5750;
   wire n_8_0_5751;
   wire n_8_0_5752;
   wire n_8_0_5753;
   wire n_8_0_5754;
   wire n_8_0_5755;
   wire n_8_0_5756;
   wire n_8_0_5757;
   wire n_8_0_5758;
   wire n_8_0_5759;
   wire n_8_0_5760;
   wire n_8_0_5761;
   wire n_8_0_5762;
   wire n_8_0_5763;
   wire n_8_0_5764;
   wire n_8_0_5765;
   wire n_8_0_5766;
   wire n_8_0_5767;
   wire n_8_0_5768;
   wire n_8_0_5769;
   wire n_8_0_5770;
   wire n_8_0_5771;
   wire n_8_0_5772;
   wire n_8_0_5773;
   wire n_8_0_5774;
   wire n_8_0_5775;
   wire n_8_0_5776;
   wire n_8_0_5777;
   wire n_8_0_5778;
   wire n_8_0_5779;
   wire n_8_0_5780;
   wire n_8_0_5781;
   wire n_8_0_5782;
   wire n_8_0_5783;
   wire n_8_0_5784;
   wire n_8_0_5785;
   wire n_8_0_5786;
   wire n_8_0_5787;
   wire n_8_0_5788;
   wire n_8_0_5789;
   wire n_8_0_5790;
   wire n_8_0_5791;
   wire n_8_0_5792;
   wire n_8_0_5793;
   wire n_8_0_5794;
   wire n_8_0_5795;
   wire n_8_0_5796;
   wire n_8_0_5797;
   wire n_8_0_5798;
   wire n_8_0_5799;
   wire n_8_0_5800;
   wire n_8_0_5801;
   wire n_8_0_5802;
   wire n_8_0_5803;
   wire n_8_0_5804;
   wire n_8_0_5805;
   wire n_8_0_5806;
   wire n_8_0_5807;
   wire n_8_0_5808;
   wire n_8_0_5809;
   wire n_8_0_5810;
   wire n_8_0_5811;
   wire n_8_0_5812;
   wire n_8_0_5813;
   wire n_8_0_5814;
   wire n_8_0_5815;
   wire n_8_0_5816;
   wire n_8_0_5817;
   wire n_8_0_5818;
   wire n_8_0_5819;
   wire n_8_0_5820;
   wire n_8_0_5821;
   wire n_8_0_5822;
   wire n_8_0_5823;
   wire n_8_0_5824;
   wire n_8_0_5825;
   wire n_8_0_5826;
   wire n_8_0_5827;
   wire n_8_0_5828;
   wire n_8_0_5829;
   wire n_8_0_5830;
   wire n_8_0_5831;
   wire n_8_0_5832;
   wire n_8_0_5833;
   wire n_8_0_5834;
   wire n_8_0_5835;
   wire n_8_0_5836;
   wire n_8_0_5837;
   wire n_8_0_5838;
   wire n_8_0_5839;
   wire n_8_0_5840;
   wire n_8_0_5841;
   wire n_8_0_5843;
   wire n_8_0_5844;
   wire n_8_0_5845;
   wire n_8_0_5846;
   wire n_8_0_5847;
   wire n_8_0_5848;
   wire n_8_0_5849;
   wire n_8_0_5850;
   wire n_8_0_5851;
   wire n_8_0_5852;
   wire n_8_0_5853;
   wire n_8_0_5854;
   wire n_8_0_5855;
   wire n_8_0_5856;
   wire n_8_0_5857;
   wire n_8_0_5858;
   wire n_8_0_5859;
   wire n_8_0_5860;
   wire n_8_0_5861;
   wire n_8_0_5862;
   wire n_8_0_5863;
   wire n_8_0_5864;
   wire n_8_0_5865;
   wire n_8_0_5866;
   wire n_8_0_5867;
   wire n_8_0_5868;
   wire n_8_0_5869;
   wire n_8_0_5870;
   wire n_8_0_5871;
   wire n_8_0_5872;
   wire n_8_0_5873;
   wire n_8_0_5874;
   wire n_8_0_5875;
   wire n_8_0_5876;
   wire n_8_0_5877;
   wire n_8_0_5878;
   wire n_8_0_5879;
   wire n_8_0_5880;
   wire n_8_0_5881;
   wire n_8_0_5882;
   wire n_8_0_5883;
   wire n_8_0_5884;
   wire n_8_0_5885;
   wire n_8_0_5886;
   wire n_8_0_5887;
   wire n_8_0_5888;
   wire n_8_0_5889;
   wire n_8_0_5890;
   wire n_8_0_5891;
   wire n_8_0_5892;
   wire n_8_0_5893;
   wire n_8_0_5894;
   wire n_8_0_5895;
   wire n_8_0_5896;
   wire n_8_0_5897;
   wire n_8_0_5898;
   wire n_8_0_5899;
   wire n_8_0_5900;
   wire n_8_0_5901;
   wire n_8_0_5902;
   wire n_8_0_5903;
   wire n_8_0_5904;
   wire n_8_0_5905;
   wire n_8_0_5906;
   wire n_8_0_5907;
   wire n_8_0_5908;
   wire n_8_0_5909;
   wire n_8_0_5910;
   wire n_8_0_5911;
   wire n_8_0_5912;
   wire n_8_0_5913;
   wire n_8_0_5915;
   wire n_8_0_5916;
   wire n_8_0_5917;
   wire n_8_0_5918;
   wire n_8_0_5919;
   wire n_8_0_5920;
   wire n_8_0_5921;
   wire n_8_0_5922;
   wire n_8_0_5923;
   wire n_8_0_5924;
   wire n_8_0_5925;
   wire n_8_0_5926;
   wire n_8_0_5927;
   wire n_8_0_5928;
   wire n_8_0_5929;
   wire n_8_0_5930;
   wire n_8_0_5931;
   wire n_8_0_5932;
   wire n_8_0_5933;
   wire n_8_0_5934;
   wire n_8_0_5935;
   wire n_8_0_5936;
   wire n_8_0_5937;
   wire n_8_0_5938;
   wire n_8_0_5939;
   wire n_8_0_5940;
   wire n_8_0_5941;
   wire n_8_0_5942;
   wire n_8_0_5943;
   wire n_8_0_5944;
   wire n_8_0_5945;
   wire n_8_0_5946;
   wire n_8_0_5947;
   wire n_8_0_5948;
   wire n_8_0_5949;
   wire n_8_0_5950;
   wire n_8_0_5951;
   wire n_8_0_5953;
   wire n_8_0_5955;
   wire n_8_0_5956;
   wire n_8_0_5957;
   wire n_8_0_5958;
   wire n_8_0_5959;
   wire n_8_0_5960;
   wire n_8_0_5961;
   wire n_8_0_5965;
   wire n_8_0_5966;
   wire n_8_0_5969;
   wire n_8_0_5970;
   wire n_8_0_5977;
   wire n_8_0_5978;
   wire n_8_0_5979;
   wire n_8_0_5980;
   wire n_8_0_5981;
   wire n_8_0_5982;
   wire n_8_0_5983;
   wire n_8_0_5984;
   wire n_8_0_5986;
   wire n_8_0_5987;
   wire n_8_0_5988;
   wire n_8_0_5989;
   wire n_8_0_5990;
   wire n_8_0_5991;
   wire n_8_0_5992;
   wire n_8_0_5994;
   wire n_8_0_5995;
   wire n_8_0_5996;
   wire n_8_0_5997;
   wire n_8_0_5998;
   wire n_8_0_5999;
   wire n_8_0_6000;
   wire n_8_0_6001;
   wire n_8_0_6002;
   wire n_8_0_6003;
   wire n_8_0_6004;
   wire n_8_0_6005;
   wire n_8_0_6006;
   wire n_8_0_6007;
   wire n_8_0_6008;
   wire n_8_0_6009;
   wire n_8_0_6010;
   wire n_8_0_6011;
   wire n_8_0_6012;
   wire n_8_0_6013;
   wire n_8_0_6014;
   wire n_8_0_6015;
   wire n_8_0_6016;
   wire n_8_0_6017;
   wire n_8_0_6018;
   wire n_8_0_6019;
   wire n_8_0_6020;
   wire n_8_0_6021;
   wire n_8_0_6022;
   wire n_8_0_6023;
   wire n_8_0_6024;
   wire n_8_0_6025;
   wire n_8_0_6026;
   wire n_8_0_6027;
   wire n_8_0_6028;
   wire n_8_0_6029;
   wire n_8_0_6030;
   wire n_8_0_6031;
   wire n_8_0_6032;
   wire n_8_0_6033;
   wire n_8_0_6034;
   wire n_8_0_6035;
   wire n_8_0_6036;
   wire n_8_0_6037;
   wire n_8_0_6038;
   wire n_8_0_6039;
   wire n_8_0_6040;
   wire n_8_0_6043;
   wire n_8_0_6044;
   wire n_8_0_6045;
   wire n_8_0_6046;
   wire n_8_0_6047;
   wire n_8_0_6048;
   wire n_8_0_6049;
   wire n_8_0_6050;
   wire n_8_0_6051;
   wire n_8_0_6052;
   wire n_8_0_6053;
   wire n_8_0_6055;
   wire n_8_0_6056;
   wire n_8_0_6057;
   wire n_8_0_6058;
   wire n_8_0_6059;
   wire n_8_0_6060;
   wire n_8_0_6061;
   wire n_8_0_6062;
   wire n_8_0_6063;
   wire n_8_0_6064;
   wire n_8_0_6065;
   wire n_8_0_6066;
   wire n_8_0_6067;
   wire n_8_0_6068;
   wire n_8_0_6069;
   wire n_8_0_6070;
   wire n_8_0_6071;
   wire n_8_0_6072;
   wire n_8_0_6073;
   wire n_8_0_6074;
   wire n_8_0_6075;
   wire n_8_0_6076;
   wire n_8_0_6077;
   wire n_8_0_6078;
   wire n_8_0_6079;
   wire n_8_0_6081;
   wire n_8_0_6082;
   wire n_8_0_6083;
   wire n_8_0_6084;
   wire n_8_0_6085;
   wire n_8_0_6086;
   wire n_8_0_6087;
   wire n_8_0_6088;
   wire n_8_0_6089;
   wire n_8_0_6090;
   wire n_8_0_6091;
   wire n_8_0_6092;
   wire n_8_0_6093;
   wire n_8_0_6094;
   wire n_8_0_6095;
   wire n_8_0_6096;
   wire n_8_0_6097;
   wire n_8_0_6098;
   wire n_8_0_6099;
   wire n_8_0_6100;
   wire n_8_0_6101;
   wire n_8_0_6106;
   wire n_8_0_6107;
   wire n_8_0_6108;
   wire n_8_0_6109;
   wire n_8_0_6111;
   wire n_8_0_6112;
   wire n_8_0_6113;
   wire n_8_0_6114;
   wire n_8_0_6120;
   wire n_8_0_6121;
   wire n_8_0_6122;
   wire n_8_0_6123;
   wire n_8_0_6125;
   wire n_8_0_6126;
   wire n_8_0_6127;
   wire n_8_0_6128;
   wire n_8_0_6130;
   wire n_8_0_6131;
   wire n_8_0_6132;
   wire n_8_0_6133;
   wire n_8_0_6134;
   wire n_8_0_6135;
   wire n_8_0_6136;
   wire n_8_0_6138;
   wire n_8_0_6139;
   wire n_8_0_6140;
   wire n_8_0_6141;
   wire n_8_0_6142;
   wire n_8_0_6143;
   wire n_8_0_6144;
   wire n_8_0_6145;
   wire n_8_0_6146;
   wire n_8_0_6147;
   wire n_8_0_6148;
   wire n_8_0_6149;
   wire n_8_0_6150;
   wire n_8_0_6151;
   wire n_8_0_6152;
   wire n_8_0_6153;
   wire n_8_0_6154;
   wire n_8_0_6155;
   wire n_8_0_6156;
   wire n_8_0_6158;
   wire n_8_0_6159;
   wire n_8_0_6160;
   wire n_8_0_6161;
   wire n_8_0_6162;
   wire n_8_0_6163;
   wire n_8_0_6164;
   wire n_8_0_6165;
   wire n_8_0_6166;
   wire n_8_0_6167;
   wire n_8_0_6168;
   wire n_8_0_6169;
   wire n_8_0_6170;
   wire n_8_0_6171;
   wire n_8_0_6172;
   wire n_8_0_6173;
   wire n_8_0_6174;
   wire n_8_0_6175;
   wire n_8_0_6180;
   wire n_8_0_6181;
   wire n_8_0_6182;
   wire n_8_0_6183;
   wire n_8_0_6184;
   wire n_8_0_6185;
   wire n_8_0_6187;
   wire n_8_0_6188;
   wire n_8_0_6189;
   wire n_8_0_6190;
   wire n_8_0_6191;
   wire n_8_0_6192;
   wire n_8_0_6194;
   wire n_8_0_6195;
   wire n_8_0_6196;
   wire n_8_0_6197;
   wire n_8_0_6198;
   wire n_8_0_6204;
   wire n_8_0_6205;
   wire n_8_0_6206;
   wire n_8_0_6208;
   wire n_8_0_6209;
   wire n_8_0_6210;
   wire n_8_0_6211;
   wire n_8_0_6213;
   wire n_8_0_6214;
   wire n_8_0_6215;
   wire n_8_0_6216;
   wire n_8_0_6217;
   wire n_8_0_6218;
   wire n_8_0_6219;
   wire n_8_0_6220;
   wire n_8_0_6221;
   wire n_8_0_6222;
   wire n_8_0_6223;
   wire n_8_0_6224;
   wire n_8_0_6225;
   wire n_8_0_6226;
   wire n_8_0_6227;
   wire n_8_0_6228;
   wire n_8_0_6229;
   wire n_8_0_6230;
   wire n_8_0_6231;
   wire n_8_0_6234;
   wire n_8_0_6235;
   wire n_8_0_6236;
   wire n_8_0_6239;
   wire n_8_0_6240;
   wire n_8_0_6241;
   wire n_8_0_6242;
   wire n_8_0_6243;
   wire n_8_0_6244;
   wire n_8_0_6245;
   wire n_8_0_6246;
   wire n_8_0_6248;
   wire n_8_0_6250;
   wire n_8_0_6251;
   wire n_8_0_6252;
   wire n_8_0_6253;
   wire n_8_0_6254;
   wire n_8_0_6255;
   wire n_8_0_6256;
   wire n_8_0_6261;
   wire n_8_0_6262;
   wire n_8_0_6263;
   wire n_8_0_6264;
   wire n_8_0_6265;
   wire n_8_0_6266;
   wire n_8_0_6267;
   wire n_8_0_6268;
   wire n_8_0_6269;
   wire n_8_0_6270;
   wire n_8_0_6271;
   wire n_8_0_6273;
   wire n_8_0_6274;
   wire n_8_0_6275;
   wire n_8_0_6281;
   wire n_8_0_6282;
   wire n_8_0_6283;
   wire n_8_0_6284;
   wire n_8_0_6285;
   wire n_8_0_6286;
   wire n_8_0_6287;
   wire n_8_0_6288;
   wire n_8_0_6290;
   wire n_8_0_6291;
   wire n_8_0_6292;
   wire n_8_0_6293;
   wire n_8_0_6294;
   wire n_8_0_6295;
   wire n_8_0_6297;
   wire n_8_0_6298;
   wire n_8_0_6299;
   wire n_8_0_6300;
   wire n_8_0_6301;
   wire n_8_0_6303;
   wire n_8_0_6304;
   wire n_8_0_6305;
   wire n_8_0_6306;
   wire n_8_0_6307;
   wire n_8_0_6308;
   wire n_8_0_6309;
   wire n_8_0_6310;
   wire n_8_0_6311;
   wire n_8_0_6312;
   wire n_8_0_6313;
   wire n_8_0_6314;
   wire n_8_0_6315;
   wire n_8_0_6316;
   wire n_8_0_6317;
   wire n_8_0_6318;
   wire n_8_0_6319;
   wire n_8_0_6320;
   wire n_8_0_6321;
   wire n_8_0_6322;
   wire n_8_0_6323;
   wire n_8_0_6324;
   wire n_8_0_6325;
   wire n_8_0_6326;
   wire n_8_0_6327;
   wire n_8_0_6328;
   wire n_8_0_6329;
   wire n_8_0_6330;
   wire n_8_0_6331;
   wire n_8_0_6332;
   wire n_8_0_6333;
   wire n_8_0_6334;
   wire n_8_0_6335;
   wire n_8_0_6336;
   wire n_8_0_6337;
   wire n_8_0_6338;
   wire n_8_0_6339;
   wire n_8_0_6340;
   wire n_8_0_6341;
   wire n_8_0_6342;
   wire n_8_0_6343;
   wire n_8_0_6344;
   wire n_8_0_6345;
   wire n_8_0_6346;
   wire n_8_0_6347;
   wire n_8_0_6348;
   wire n_8_0_6349;
   wire n_8_0_6350;
   wire n_8_0_6351;
   wire n_8_0_6352;
   wire n_8_0_6353;
   wire n_8_0_6354;
   wire n_8_0_6355;
   wire n_8_0_6356;
   wire n_8_0_6357;
   wire n_8_0_6358;
   wire n_8_0_6359;
   wire n_8_0_6360;
   wire n_8_0_6363;
   wire n_8_0_6364;
   wire n_8_0_6365;
   wire n_8_0_6366;
   wire n_8_0_6367;
   wire n_8_0_6368;
   wire n_8_0_6369;
   wire n_8_0_6370;
   wire n_8_0_6371;
   wire n_8_0_6372;
   wire n_8_0_6373;
   wire n_8_0_6374;
   wire n_8_0_6375;
   wire n_8_0_6376;
   wire n_8_0_6379;
   wire n_8_0_6380;
   wire n_8_0_6381;
   wire n_8_0_6382;
   wire n_8_0_6384;
   wire n_8_0_6385;
   wire n_8_0_6386;
   wire n_8_0_6387;
   wire n_8_0_6390;
   wire n_8_0_6391;
   wire n_8_0_6392;
   wire n_8_0_6393;
   wire n_8_0_6394;
   wire n_8_0_6395;
   wire n_8_0_6397;
   wire n_8_0_6398;
   wire n_8_0_6399;
   wire n_8_0_6400;
   wire n_8_0_6405;
   wire n_8_0_6407;
   wire n_8_0_6408;
   wire n_8_0_6409;
   wire n_8_0_6411;
   wire n_8_0_6412;
   wire n_8_0_6413;
   wire n_8_0_6414;
   wire n_8_0_6416;
   wire n_8_0_6417;
   wire n_8_0_6418;
   wire n_8_0_6419;
   wire n_8_0_6420;
   wire n_8_0_6421;
   wire n_8_0_6422;
   wire n_8_0_6423;
   wire n_8_0_6424;
   wire n_8_0_6425;
   wire n_8_0_6426;
   wire n_8_0_6427;
   wire n_8_0_6428;
   wire n_8_0_6429;
   wire n_8_0_6430;
   wire n_8_0_6431;
   wire n_8_0_6432;
   wire n_8_0_6433;
   wire n_8_0_6434;
   wire n_8_0_6435;
   wire n_8_0_6436;
   wire n_8_0_6437;
   wire n_8_0_6438;
   wire n_8_0_6439;
   wire n_8_0_6440;
   wire n_8_0_6441;
   wire n_8_0_6442;
   wire n_8_0_6443;
   wire n_8_0_6444;
   wire n_8_0_6445;
   wire n_8_0_6446;
   wire n_8_0_6447;
   wire n_8_0_6448;
   wire n_8_0_6449;
   wire n_8_0_6450;
   wire n_8_0_6451;
   wire n_8_0_6452;
   wire n_8_0_6453;
   wire n_8_0_6454;
   wire n_8_0_6455;
   wire n_8_0_6456;
   wire n_8_0_6457;
   wire n_8_0_6458;
   wire n_8_0_6459;
   wire n_8_0_6460;
   wire n_8_0_6461;
   wire n_8_0_6462;
   wire n_8_0_6463;
   wire n_8_0_6464;
   wire n_8_0_6472;
   wire n_8_0_6473;
   wire n_8_0_6474;
   wire n_8_0_6475;
   wire n_8_0_6476;
   wire n_8_0_6477;
   wire n_8_0_6478;
   wire n_8_0_6479;
   wire n_8_0_6480;
   wire n_8_0_6481;
   wire n_8_0_6482;
   wire n_8_0_6483;
   wire n_8_0_6484;
   wire n_8_0_6485;
   wire n_8_0_6486;
   wire n_8_0_6487;
   wire n_8_0_6488;
   wire n_8_0_6489;
   wire n_8_0_6490;
   wire n_8_0_6491;
   wire n_8_0_6492;
   wire n_8_0_6493;
   wire n_8_0_6494;
   wire n_8_0_6495;
   wire n_8_0_6496;
   wire n_8_0_6497;
   wire n_8_0_6498;
   wire n_8_0_6499;
   wire n_8_0_6500;
   wire n_8_0_6501;
   wire n_8_0_6502;
   wire n_8_0_6503;
   wire n_8_0_6504;
   wire n_8_0_6505;
   wire n_8_0_6506;
   wire n_8_0_6507;
   wire n_8_0_6508;
   wire n_8_0_6509;
   wire n_8_0_6510;
   wire n_8_0_6511;
   wire n_8_0_6512;
   wire n_8_0_6513;
   wire n_8_0_6514;
   wire n_8_0_6515;
   wire n_8_0_6516;
   wire n_8_0_6517;
   wire n_8_0_6518;
   wire n_8_0_6519;
   wire n_8_0_6521;
   wire n_8_0_6522;
   wire n_8_0_6523;
   wire n_8_0_6524;
   wire n_8_0_6525;
   wire n_8_0_6526;
   wire n_8_0_6527;
   wire n_8_0_6528;
   wire n_8_0_6529;
   wire n_8_0_6530;
   wire n_8_0_6531;
   wire n_8_0_6532;
   wire n_8_0_6533;
   wire n_8_0_6534;
   wire n_8_0_6535;
   wire n_8_0_6536;
   wire n_8_0_6537;
   wire n_8_0_6538;
   wire n_8_0_6539;
   wire n_8_0_6542;
   wire n_8_0_6543;
   wire n_8_0_6544;
   wire n_8_0_6545;
   wire n_8_0_6546;
   wire n_8_0_6547;
   wire n_8_0_6548;
   wire n_8_0_6549;
   wire n_8_0_6550;
   wire n_8_0_6551;
   wire n_8_0_6552;
   wire n_8_0_6553;
   wire n_8_0_6554;
   wire n_8_0_6555;
   wire n_8_0_6556;
   wire n_8_0_6557;
   wire n_8_0_6558;
   wire n_8_0_6559;
   wire n_8_0_6560;
   wire n_8_0_6561;
   wire n_8_0_6562;
   wire n_8_0_6563;
   wire n_8_0_6564;
   wire n_8_0_6565;
   wire n_8_0_6566;
   wire n_8_0_6569;
   wire n_8_0_6570;
   wire n_8_0_6571;
   wire n_8_0_6572;
   wire n_8_0_6573;
   wire n_8_0_6574;
   wire n_8_0_6575;
   wire n_8_0_6576;
   wire n_8_0_6577;
   wire n_8_0_6578;
   wire n_8_0_6579;
   wire n_8_0_6580;
   wire n_8_0_6581;
   wire n_8_0_6583;
   wire n_8_0_6584;
   wire n_8_0_6585;
   wire n_8_0_6586;
   wire n_8_0_6587;
   wire n_8_0_6588;
   wire n_8_0_6589;
   wire n_8_0_6590;
   wire n_8_0_6591;
   wire n_8_0_6592;
   wire n_8_0_6594;
   wire n_8_0_6596;
   wire n_8_0_6598;
   wire n_8_0_6599;
   wire n_8_0_6600;
   wire n_8_0_6601;
   wire n_8_0_6603;
   wire n_8_0_6604;
   wire n_8_0_6605;
   wire n_8_0_6606;
   wire n_8_0_6607;
   wire n_8_0_6608;
   wire n_8_0_6609;
   wire n_8_0_6610;
   wire n_8_0_6611;
   wire n_8_0_6612;
   wire n_8_0_6613;
   wire n_8_0_6617;
   wire n_8_0_6618;
   wire n_8_0_6619;
   wire n_8_0_6620;
   wire n_8_0_6621;
   wire n_8_0_6622;
   wire n_8_0_6623;
   wire n_8_0_6624;
   wire n_8_0_6625;
   wire n_8_0_6626;
   wire n_8_0_6627;
   wire n_8_0_6628;
   wire n_8_0_6629;
   wire n_8_0_6630;
   wire n_8_0_6631;
   wire n_8_0_6632;
   wire n_8_0_6633;
   wire n_8_0_6634;
   wire n_8_0_6635;
   wire n_8_0_6636;
   wire n_8_0_6637;
   wire n_8_0_6638;
   wire n_8_0_6639;
   wire n_8_0_6640;
   wire n_8_0_6641;
   wire n_8_0_6642;
   wire n_8_0_6643;
   wire n_8_0_6644;
   wire n_8_0_6645;
   wire n_8_0_6646;
   wire n_8_0_6647;
   wire n_8_0_6648;
   wire n_8_0_6649;
   wire n_8_0_6650;
   wire n_8_0_6651;
   wire n_8_0_6652;
   wire n_8_0_6653;
   wire n_8_0_6654;
   wire n_8_0_6655;
   wire n_8_0_6656;
   wire n_8_0_6657;
   wire n_8_0_6658;
   wire n_8_0_6659;
   wire n_8_0_6660;
   wire n_8_0_6661;
   wire n_8_0_6662;
   wire n_8_0_6663;
   wire n_8_0_6664;
   wire n_8_0_6665;
   wire n_8_0_6666;
   wire n_8_0_6667;
   wire n_8_0_6668;
   wire n_8_0_6669;
   wire n_8_0_6670;
   wire n_8_0_6671;
   wire n_8_0_6672;
   wire n_8_0_6673;
   wire n_8_0_6674;
   wire n_8_0_6675;
   wire n_8_0_6676;
   wire n_8_0_6677;
   wire n_8_0_6678;
   wire n_8_0_6679;
   wire n_8_0_6680;
   wire n_8_0_6681;
   wire n_8_0_6682;
   wire n_8_0_6683;
   wire n_8_0_6684;
   wire n_8_0_6685;
   wire n_8_0_6686;
   wire n_8_0_6687;
   wire n_8_0_6688;
   wire n_8_0_6689;
   wire n_8_0_6690;
   wire n_8_0_6691;
   wire n_8_0_6692;
   wire n_8_0_6693;
   wire n_8_0_6694;
   wire n_8_0_6695;
   wire n_8_0_6696;
   wire n_8_0_6697;
   wire n_8_0_6698;
   wire n_8_0_6699;
   wire n_8_0_6700;
   wire n_8_0_6701;
   wire n_8_0_6702;
   wire n_8_0_6703;
   wire n_8_0_6704;
   wire n_8_0_6705;
   wire n_8_0_6706;
   wire n_8_0_6707;
   wire n_8_0_6708;
   wire n_8_0_6709;
   wire n_8_0_6710;
   wire n_8_0_6711;
   wire n_8_0_6712;
   wire n_8_0_6713;
   wire n_8_0_6716;
   wire n_8_0_6717;
   wire n_8_0_6718;
   wire n_8_0_6722;
   wire n_8_0_6723;
   wire n_8_0_6725;
   wire n_8_0_6726;
   wire n_8_0_6728;
   wire n_8_0_6739;
   wire n_8_0_6740;
   wire n_8_0_6741;
   wire n_8_0_6742;
   wire n_8_0_6743;
   wire n_8_0_6744;
   wire n_8_0_6745;
   wire n_8_0_6746;
   wire n_8_0_6747;
   wire n_8_0_6748;
   wire n_8_0_6749;
   wire n_8_0_6750;
   wire n_8_0_6751;
   wire n_8_0_6753;
   wire n_8_0_6754;
   wire n_8_0_6756;
   wire n_8_0_6757;
   wire n_8_0_6758;
   wire n_8_0_6759;
   wire n_8_0_6760;
   wire n_8_0_6761;
   wire n_8_0_6762;
   wire n_8_0_6763;
   wire n_8_0_6764;
   wire n_8_0_6765;
   wire n_8_0_6766;
   wire n_8_0_6767;
   wire n_8_0_6768;
   wire n_8_0_6769;
   wire n_8_0_6770;
   wire n_8_0_6771;
   wire n_8_0_6772;
   wire n_8_0_6773;
   wire n_8_0_6774;
   wire n_8_0_6775;
   wire n_8_0_6776;
   wire n_8_0_6777;
   wire n_8_0_6778;
   wire n_8_0_6779;
   wire n_8_0_6780;
   wire n_8_0_6781;
   wire n_8_0_6782;
   wire n_8_0_6783;
   wire n_8_0_6784;
   wire n_8_0_6785;
   wire n_8_0_6786;
   wire n_8_0_6787;
   wire n_8_0_6788;
   wire n_8_0_6789;
   wire n_8_0_6790;
   wire n_8_0_6791;
   wire n_8_0_6792;
   wire n_8_0_6793;
   wire n_8_0_6794;
   wire n_8_0_6795;
   wire n_8_0_6796;
   wire n_8_0_6797;
   wire n_8_0_6798;
   wire n_8_0_6799;
   wire n_8_0_6800;
   wire n_8_0_6801;
   wire n_8_0_6802;
   wire n_8_0_6803;
   wire n_8_0_6804;
   wire n_8_0_6805;
   wire n_8_0_6806;
   wire n_8_0_6807;
   wire n_8_0_6808;
   wire n_8_0_6809;
   wire n_8_0_6810;
   wire n_8_0_6812;
   wire n_8_0_6813;
   wire n_8_0_6814;
   wire n_8_0_6815;
   wire n_8_0_6816;
   wire n_8_0_6817;
   wire n_8_0_6818;
   wire n_8_0_6819;
   wire n_8_0_6820;
   wire n_8_0_6821;
   wire n_8_0_6822;
   wire n_8_0_6823;
   wire n_8_0_6824;
   wire n_8_0_6825;
   wire n_8_0_6826;
   wire n_8_0_6827;
   wire n_8_0_6828;
   wire n_8_0_6829;
   wire n_8_0_6830;
   wire n_8_0_6831;
   wire n_8_0_6832;
   wire n_8_0_6833;
   wire n_8_0_6834;
   wire n_8_0_6835;
   wire n_8_0_6836;
   wire n_8_0_6837;
   wire n_8_0_6838;
   wire n_8_0_6839;
   wire n_8_0_6840;
   wire n_8_0_6841;
   wire n_8_0_6842;
   wire n_8_0_6843;
   wire n_8_0_6844;
   wire n_8_0_6845;
   wire n_8_0_6846;
   wire n_8_0_6847;
   wire n_8_0_6848;
   wire n_8_0_6849;
   wire n_8_0_6850;
   wire n_8_0_6851;
   wire n_8_0_6852;
   wire n_8_0_6855;
   wire n_8_0_6856;
   wire n_8_0_6857;
   wire n_8_0_6858;
   wire n_8_0_6860;
   wire n_8_0_6861;
   wire n_8_0_6862;
   wire n_8_0_6863;
   wire n_8_0_6864;
   wire n_8_0_6865;
   wire n_8_0_6867;
   wire n_8_0_6869;
   wire n_8_0_6873;
   wire n_8_0_6874;
   wire n_8_0_6875;
   wire n_8_0_6876;
   wire n_8_0_6877;
   wire n_8_0_6878;
   wire n_8_0_6879;
   wire n_8_0_6880;
   wire n_8_0_6881;
   wire n_8_0_6882;
   wire n_8_0_6883;
   wire n_8_0_6884;
   wire n_8_0_6885;
   wire n_8_0_6886;
   wire n_8_0_6887;
   wire n_8_0_6888;
   wire n_8_0_6889;
   wire n_8_0_6890;
   wire n_8_0_6891;
   wire n_8_0_6892;
   wire n_8_0_6893;
   wire n_8_0_6894;
   wire n_8_0_6895;
   wire n_8_0_6896;
   wire n_8_0_6897;
   wire n_8_0_6898;
   wire n_8_0_6899;
   wire n_8_0_6900;
   wire n_8_0_6901;
   wire n_8_0_6902;
   wire n_8_0_6903;
   wire n_8_0_6904;
   wire n_8_0_6905;
   wire n_8_0_6906;
   wire n_8_0_6907;
   wire n_8_0_6908;
   wire n_8_0_6909;
   wire n_8_0_6910;
   wire n_8_0_6911;
   wire n_8_0_6912;
   wire n_8_0_6913;
   wire n_8_0_6914;
   wire n_8_0_6915;
   wire n_8_0_6916;
   wire n_8_0_6917;
   wire n_8_0_6918;
   wire n_8_0_6919;
   wire n_8_0_6920;
   wire n_8_0_6921;
   wire n_8_0_6922;
   wire n_8_0_6923;
   wire n_8_0_6924;
   wire n_8_0_6925;
   wire n_8_0_6926;
   wire n_8_0_6927;
   wire n_8_0_6928;
   wire n_8_0_6929;
   wire n_8_0_6930;
   wire n_8_0_6931;
   wire n_8_0_6932;
   wire n_8_0_6933;
   wire n_8_0_6934;
   wire n_8_0_6935;
   wire n_8_0_6936;
   wire n_8_0_6937;
   wire n_8_0_6938;
   wire n_8_0_6939;
   wire n_8_0_6940;
   wire n_8_0_6941;
   wire n_8_0_6942;
   wire n_8_0_6943;
   wire n_8_0_6944;
   wire n_8_0_6945;
   wire n_8_0_6946;
   wire n_8_0_6947;
   wire n_8_0_6948;
   wire n_8_0_6949;
   wire n_8_0_6950;
   wire n_8_0_6951;
   wire n_8_0_6952;
   wire n_8_0_6953;
   wire n_8_0_6954;
   wire n_8_0_6955;
   wire n_8_0_6956;
   wire n_8_0_6957;
   wire n_8_0_6958;
   wire n_8_0_6959;
   wire n_8_0_6960;
   wire n_8_0_6961;
   wire n_8_0_6962;
   wire n_8_0_6963;
   wire n_8_0_6964;
   wire n_8_0_6965;
   wire n_8_0_6966;
   wire n_8_0_6967;
   wire n_8_0_6968;
   wire n_8_0_6969;
   wire n_8_0_6970;
   wire n_8_0_6971;
   wire n_8_0_6972;
   wire n_8_0_6973;
   wire n_8_0_6974;
   wire n_8_0_6975;
   wire n_8_0_6976;
   wire n_8_0_6977;
   wire n_8_0_6978;
   wire n_8_0_6979;
   wire n_8_0_6980;
   wire n_8_0_6981;
   wire n_8_0_6982;
   wire n_8_0_6983;
   wire n_8_0_6984;
   wire n_8_0_6985;
   wire n_8_0_6986;
   wire n_8_0_6990;
   wire n_8_0_6991;
   wire n_8_0_6992;
   wire n_8_0_6993;
   wire n_8_0_6994;
   wire n_8_0_6995;
   wire n_8_0_7002;
   wire n_8_0_7006;
   wire n_8_0_7007;
   wire n_8_0_7008;
   wire n_8_0_7009;
   wire n_8_0_7010;
   wire n_8_0_7011;
   wire n_8_0_7012;
   wire n_8_0_7013;
   wire n_8_0_7014;
   wire n_8_0_7015;
   wire n_8_0_7016;
   wire n_8_0_7017;
   wire n_8_0_7018;
   wire n_8_0_7019;
   wire n_8_0_7020;
   wire n_8_0_7021;
   wire n_8_0_7022;
   wire n_8_0_7023;
   wire n_8_0_7024;
   wire n_8_0_7025;
   wire n_8_0_7026;
   wire n_8_0_7027;
   wire n_8_0_7028;
   wire n_8_0_7029;
   wire n_8_0_7030;
   wire n_8_0_7031;
   wire n_8_0_7032;
   wire n_8_0_7033;
   wire n_8_0_7034;
   wire n_8_0_7035;
   wire n_8_0_7036;
   wire n_8_0_7037;
   wire n_8_0_7038;
   wire n_8_0_7039;
   wire n_8_0_7040;
   wire n_8_0_7041;
   wire n_8_0_7042;
   wire n_8_0_7043;
   wire n_8_0_7044;
   wire n_8_0_7045;
   wire n_8_0_7046;
   wire n_8_0_7047;
   wire n_8_0_7048;
   wire n_8_0_7049;
   wire n_8_0_7050;
   wire n_8_0_7051;
   wire n_8_0_7052;
   wire n_8_0_7053;
   wire n_8_0_7054;
   wire n_8_0_7055;
   wire n_8_0_7056;
   wire n_8_0_7057;
   wire n_8_0_7058;
   wire n_8_0_7059;
   wire n_8_0_7060;
   wire n_8_0_7061;
   wire n_8_0_7062;
   wire n_8_0_7063;
   wire n_8_0_7064;
   wire n_8_0_7065;
   wire n_8_0_7066;
   wire n_8_0_7067;
   wire n_8_0_7068;
   wire n_8_0_7069;
   wire n_8_0_7070;
   wire n_8_0_7071;
   wire n_8_0_7072;
   wire n_8_0_7073;
   wire n_8_0_7074;
   wire n_8_0_7075;
   wire n_8_0_7076;
   wire n_8_0_7077;
   wire n_8_0_7078;
   wire n_8_0_7079;
   wire n_8_0_7080;
   wire n_8_0_7081;
   wire n_8_0_7082;
   wire n_8_0_7083;
   wire n_8_0_7084;
   wire n_8_0_7085;
   wire n_8_0_7086;
   wire n_8_0_7087;
   wire n_8_0_7088;
   wire n_8_0_7089;
   wire n_8_0_4314;
   wire n_8_0_1484;
   wire n_8_0_1527;
   wire n_8_0_1528;
   wire n_8_0_1529;
   wire n_8_0_1589;
   wire n_8_0_1590;
   wire n_8_0_1599;
   wire n_8_0_1600;
   wire n_8_0_4330;
   wire n_8_0_4303;
   wire n_8_0_4328;
   wire n_8_0_1607;
   wire n_8_0_1616;
   wire n_8_0_1617;
   wire n_8_0_1656;
   wire n_8_0_4600;
   wire n_8_0_1657;
   wire n_8_0_4531;
   wire n_8_0_4597;
   wire n_8_0_4501;
   wire n_8_0_4292;
   wire n_8_0_4290;
   wire n_8_0_4257;
   wire n_8_0_4050;
   wire n_8_0_4022;
   wire n_8_0_3939;
   wire n_8_0_1734;
   wire n_8_0_3008;
   wire n_8_0_3004;
   wire n_8_0_1735;
   wire n_8_0_1736;
   wire n_8_0_1737;
   wire n_8_0_1753;
   wire n_8_0_1754;
   wire n_8_0_1755;
   wire n_8_0_1774;
   wire n_8_0_1782;
   wire n_8_0_1783;
   wire n_8_0_1873;
   wire n_8_0_4312;
   wire n_8_0_1883;
   wire n_8_0_1884;
   wire n_8_0_6278;
   wire n_8_0_1904;
   wire n_8_0_1905;
   wire n_8_0_1944;
   wire n_8_0_1945;
   wire n_8_0_1946;
   wire n_8_0_1972;
   wire n_8_0_1973;
   wire n_8_0_3003;
   wire n_8_0_3011;
   wire n_8_0_2998;
   wire n_8_0_2541;
   wire n_8_0_2994;
   wire n_8_0_2992;
   wire n_8_0_3007;
   wire n_8_0_2542;
   wire n_8_0_2544;
   wire n_8_0_2545;
   wire n_8_0_2737;
   wire n_8_0_2752;
   wire n_8_0_3752;
   wire n_8_0_2754;
   wire n_8_0_2755;
   wire n_8_0_2756;
   wire n_8_0_5594;
   wire n_8_0_2918;
   wire n_8_0_2919;
   wire n_8_0_2920;
   wire n_8_0_2944;
   wire n_8_0_2946;
   wire n_8_0_5724;
   wire n_8_0_2980;
   wire n_8_0_3878;
   wire n_8_0_3887;
   wire n_8_0_3889;
   wire n_8_0_3883;
   wire n_8_0_2989;
   wire n_8_0_2990;
   wire n_8_0_2991;
   wire n_8_0_3002;
   wire n_8_0_3893;
   wire n_8_0_3895;
   wire n_8_0_3899;
   wire n_8_0_3009;
   wire n_8_0_3014;
   wire n_8_0_5976;
   wire n_8_0_3074;
   wire n_8_0_3075;
   wire n_8_0_3079;
   wire n_8_0_3080;
   wire n_8_0_3934;
   wire n_8_0_3923;
   wire n_8_0_3928;
   wire n_8_0_3081;
   wire n_8_0_3090;
   wire n_8_0_3098;
   wire n_8_0_3099;
   wire n_8_0_3100;
   wire n_8_0_3998;
   wire n_8_0_4013;
   wire n_8_0_3115;
   wire n_8_0_3116;
   wire n_8_0_3117;
   wire n_8_0_3123;
   wire n_8_0_3124;
   wire n_8_0_4035;
   wire n_8_0_4033;
   wire n_8_0_4025;
   wire n_8_0_3128;
   wire n_8_0_4040;
   wire n_8_0_4043;
   wire n_8_0_3140;
   wire n_8_0_3141;
   wire n_8_0_3174;
   wire n_8_0_3175;
   wire n_8_0_3176;
   wire n_8_0_3205;
   wire n_8_0_3210;
   wire n_8_0_3212;
   wire n_8_0_3213;
   wire n_8_0_4065;
   wire n_8_0_4053;
   wire n_8_0_4056;
   wire n_8_0_3214;
   wire n_8_0_3215;
   wire n_8_0_3238;
   wire n_8_0_3239;
   wire n_8_0_5952;
   wire n_8_0_3242;
   wire n_8_0_3276;
   wire n_8_0_3277;
   wire n_8_0_3278;
   wire n_8_0_3279;
   wire n_8_0_4260;
   wire n_8_0_4272;
   wire n_8_0_4247;
   wire n_8_0_4250;
   wire n_8_0_4252;
   wire n_8_0_3282;
   wire n_8_0_3303;
   wire n_8_0_3309;
   wire n_8_0_3328;
   wire n_8_0_3330;
   wire n_8_0_3336;
   wire n_8_0_3337;
   wire n_8_0_3354;
   wire n_8_0_3355;
   wire n_8_0_3357;
   wire n_8_0_3375;
   wire n_8_0_3376;
   wire n_8_0_3377;
   wire n_8_0_3460;
   wire n_8_0_3461;
   wire n_8_0_6237;
   wire n_8_0_3474;
   wire n_8_0_3475;
   wire n_8_0_3476;
   wire n_8_0_4596;
   wire n_8_0_3484;
   wire n_8_0_3544;
   wire n_8_0_3545;
   wire n_8_0_3546;
   wire n_8_0_3555;
   wire n_8_0_3556;
   wire n_8_0_6520;
   wire n_8_0_6597;
   wire n_8_0_3569;
   wire n_8_0_3570;
   wire n_8_0_4514;
   wire n_8_0_3573;
   wire n_8_0_3581;
   wire n_8_0_4504;
   wire n_8_0_3582;
   wire n_8_0_3599;
   wire n_8_0_3600;
   wire n_8_0_3602;
   wire n_8_0_3603;
   wire n_8_0_6541;
   wire n_8_0_3604;
   wire n_8_0_3605;
   wire n_8_0_3624;
   wire n_8_0_3678;
   wire n_8_0_3679;
   wire n_8_0_3680;
   wire n_8_0_3690;
   wire n_8_0_4583;
   wire n_8_0_3698;
   wire n_8_0_4589;
   wire n_8_0_4594;
   wire n_8_0_3708;
   wire n_8_0_3709;
   wire n_8_0_6719;
   wire n_8_0_3710;
   wire n_8_0_3711;
   wire n_8_0_3751;
   wire n_8_0_3755;
   wire n_8_0_3756;
   wire n_8_0_4184;
   wire n_8_0_6989;
   wire n_8_0_3757;
   wire n_8_0_3758;
   wire n_8_0_3759;
   wire n_8_0_3762;
   wire n_8_0_3810;
   wire n_8_0_3811;
   wire n_8_0_3812;
   wire n_8_0_3819;
   wire n_8_0_3820;
   wire n_8_0_3821;
   wire n_8_0_3839;
   wire n_8_0_3840;
   wire n_8_0_3853;
   wire n_8_0_3854;
   wire n_8_0_3863;
   wire n_8_0_3866;
   wire n_8_0_3876;
   wire n_8_0_3877;
   wire n_8_0_4181;
   wire n_8_0_4178;
   wire n_8_0_3881;
   wire n_8_0_4187;
   wire n_8_0_3882;
   wire n_8_0_3884;
   wire n_8_0_3885;
   wire n_8_0_6404;
   wire n_8_0_6361;
   wire n_8_0_6469;
   wire n_8_0_6721;
   wire n_8_0_6471;
   wire n_8_0_3657;
   wire n_8_0_5914;
   wire n_8_0_5842;
   wire n_8_0_5652;
   wire n_8_0_4423;
   wire n_8_0_6714;
   wire n_8_0_6410;
   wire n_8_0_6276;
   wire n_8_0_5971;
   wire n_8_0_5423;
   wire n_8_0_5392;
   wire n_8_0_5405;
   wire n_8_0_5362;
   wire n_8_0_5374;
   wire n_8_0_5186;
   wire n_8_0_4375;
   wire n_8_0_4211;
   wire n_8_0_4100;
   wire n_8_0_4079;
   wire n_8_0_3904;
   wire n_8_0_3587;
   wire n_8_0_3591;
   wire n_8_0_3548;
   wire n_8_0_3558;
   wire n_8_0_3302;
   wire n_8_0_3298;
   wire n_8_0_3200;
   wire n_8_0_3142;
   wire n_8_0_3139;
   wire n_8_0_3102;
   wire n_8_0_3114;
   wire n_8_0_3085;
   wire n_8_0_3095;
   wire n_8_0_2753;
   wire n_8_0_3886;
   wire n_8_0_3892;
   wire n_8_0_2979;
   wire n_8_0_3903;
   wire n_8_0_3905;
   wire n_8_0_3906;
   wire n_8_0_3907;
   wire n_8_0_3917;
   wire n_8_0_3918;
   wire n_8_0_3285;
   wire n_8_0_3919;
   wire n_8_0_3940;
   wire n_8_0_3941;
   wire n_8_0_3995;
   wire n_8_0_3996;
   wire n_8_0_4002;
   wire n_8_0_4003;
   wire n_8_0_4020;
   wire n_8_0_4021;
   wire n_8_0_4023;
   wire n_8_0_4024;
   wire n_8_0_4037;
   wire n_8_0_4046;
   wire n_8_0_4047;
   wire n_8_0_4048;
   wire n_8_0_4051;
   wire n_8_0_4052;
   wire n_8_0_4075;
   wire n_8_0_4076;
   wire n_8_0_4077;
   wire n_8_0_4080;
   wire n_8_0_4081;
   wire n_8_0_4116;
   wire n_8_0_4136;
   wire n_8_0_4137;
   wire n_8_0_4156;
   wire n_8_0_4160;
   wire n_8_0_4161;
   wire n_8_0_4162;
   wire n_8_0_4163;
   wire n_8_0_4164;
   wire n_8_0_4185;
   wire n_8_0_4190;
   wire n_8_0_4206;
   wire n_8_0_4207;
   wire n_8_0_4246;
   wire n_8_0_4256;
   wire n_8_0_4258;
   wire n_8_0_4115;
   wire n_8_0_4266;
   wire n_8_0_4275;
   wire n_8_0_4276;
   wire n_8_0_4277;
   wire n_8_0_4291;
   wire n_8_0_4294;
   wire n_8_0_4301;
   wire n_8_0_4302;
   wire n_8_0_4318;
   wire n_8_0_4332;
   wire n_8_0_4333;
   wire n_8_0_4334;
   wire n_8_0_4355;
   wire n_8_0_4356;
   wire n_8_0_4371;
   wire n_8_0_4372;
   wire n_8_0_4379;
   wire n_8_0_4388;
   wire n_8_0_4404;
   wire n_8_0_4408;
   wire n_8_0_4410;
   wire n_8_0_4444;
   wire n_8_0_4459;
   wire n_8_0_4460;
   wire n_8_0_4469;
   wire n_8_0_4470;
   wire n_8_0_6988;
   wire n_8_0_4474;
   wire n_8_0_4475;
   wire n_8_0_4476;
   wire n_8_0_4500;
   wire n_8_0_4502;
   wire n_8_0_2761;
   wire n_8_0_2758;
   wire n_8_0_4566;
   wire n_8_0_2765;
   wire n_8_0_4567;
   wire n_8_0_4568;
   wire n_8_0_4569;
   wire n_8_0_4613;
   wire n_8_0_4614;
   wire n_8_0_2982;
   wire n_8_0_4615;
   wire n_8_0_4616;
   wire n_8_0_4814;
   wire n_8_0_4815;
   wire n_8_0_4821;
   wire n_8_0_4822;
   wire n_8_0_4830;
   wire n_8_0_4844;
   wire n_8_0_4845;
   wire n_8_0_2935;
   wire n_8_0_2939;
   wire n_8_0_2928;
   wire n_8_0_4846;
   wire n_8_0_2943;
   wire n_8_0_4847;
   wire n_8_0_2981;
   wire n_8_0_4849;
   wire n_8_0_4850;
   wire n_8_0_5059;
   wire n_8_0_5060;
   wire n_8_0_5061;
   wire n_8_0_5062;
   wire n_8_0_5063;
   wire n_8_0_5064;
   wire n_8_0_5068;
   wire n_8_0_5171;
   wire n_8_0_5172;
   wire n_8_0_5173;
   wire n_8_0_5174;
   wire n_8_0_5175;
   wire n_8_0_5356;
   wire n_8_0_5357;
   wire n_8_0_5358;
   wire n_8_0_5359;
   wire n_8_0_5361;
   wire n_8_0_5380;
   wire n_8_0_5381;
   wire n_8_0_5391;
   wire n_8_0_5401;
   wire n_8_0_5402;
   wire n_8_0_5410;
   wire n_8_0_5411;
   wire n_8_0_5412;
   wire n_8_0_5413;
   wire n_8_0_5437;
   wire n_8_0_5962;
   wire n_8_0_5963;
   wire n_8_0_6859;
   wire n_8_0_5964;
   wire n_8_0_5967;
   wire n_8_0_5968;
   wire n_8_0_5972;
   wire n_8_0_3145;
   wire n_8_0_5974;
   wire n_8_0_6102;
   wire n_8_0_6103;
   wire n_8_0_6104;
   wire n_8_0_6116;
   wire n_8_0_6119;
   wire n_8_0_6137;
   wire n_8_0_6176;
   wire n_8_0_6177;
   wire n_8_0_3187;
   wire n_8_0_6178;
   wire n_8_0_3177;
   wire n_8_0_3196;
   wire n_8_0_6200;
   wire n_8_0_3209;
   wire n_8_0_6202;
   wire n_8_0_6238;
   wire n_8_0_3211;
   wire n_8_0_6257;
   wire n_8_0_6258;
   wire n_8_0_6259;
   wire n_8_0_6260;
   wire n_8_0_6277;
   wire n_8_0_6377;
   wire n_8_0_3231;
   wire n_8_0_3228;
   wire n_8_0_3219;
   wire n_8_0_3235;
   wire n_8_0_3241;
   wire n_8_0_6388;
   wire n_8_0_3244;
   wire n_8_0_3243;
   wire n_8_0_6402;
   wire n_8_0_6415;
   wire n_8_0_6470;
   wire n_8_0_6567;
   wire n_8_0_6568;
   wire n_8_0_6615;
   wire n_8_0_3280;
   wire n_8_0_3296;
   wire n_8_0_6616;
   wire n_8_0_6720;
   wire n_8_0_6732;
   wire n_8_0_6733;
   wire n_8_0_6734;
   wire n_8_0_6080;
   wire n_8_0_6735;
   wire n_8_0_3352;
   wire n_8_0_6736;
   wire n_8_0_6737;
   wire n_8_0_6738;
   wire n_8_0_6866;
   wire n_8_0_6868;
   wire n_8_0_6870;
   wire n_8_0_6871;
   wire n_8_0_3372;
   wire n_8_0_3365;
   wire n_8_0_6872;
   wire n_8_0_6987;
   wire n_8_0_7001;
   wire n_8_0_7005;
   wire n_8_0_7090;
   wire n_8_0_6201;
   wire n_8_0_7091;
   wire n_8_0_7092;
   wire n_8_0_7093;
   wire n_8_0_7094;
   wire n_8_0_3468;
   wire n_8_0_7095;
   wire n_8_0_7096;
   wire n_8_0_7097;
   wire n_8_0_3478;
   wire n_8_0_7098;
   wire n_8_0_3692;
   wire n_8_0_7099;
   wire n_8_0_7100;
   wire n_8_0_7101;
   wire n_8_0_3477;
   wire n_8_0_7102;
   wire n_8_0_4422;
   wire n_8_0_7103;
   wire n_8_0_7104;
   wire n_8_0_7105;
   wire n_8_0_7106;
   wire n_8_0_7107;
   wire n_8_0_7108;
   wire n_8_0_7109;
   wire n_8_0_3561;
   wire n_8_0_3566;
   wire n_8_0_7110;
   wire n_8_0_7111;
   wire n_8_0_7112;
   wire n_8_0_7113;
   wire n_8_0_3557;
   wire n_8_0_3554;
   wire n_8_0_7114;
   wire n_8_0_7115;
   wire n_8_0_7116;
   wire n_8_0_7117;
   wire n_8_0_7118;
   wire n_8_0_7119;
   wire n_8_0_7120;
   wire n_8_0_7121;
   wire n_8_0_7122;
   wire n_8_0_7123;
   wire n_8_0_7124;
   wire n_8_0_7125;
   wire n_8_0_7126;
   wire n_8_0_7127;
   wire n_8_0_7128;
   wire n_8_0_3577;
   wire n_8_0_7129;
   wire n_8_0_3594;
   wire n_8_0_3574;
   wire n_8_0_3580;
   wire n_8_0_7130;
   wire n_8_0_7131;
   wire n_8_0_7132;
   wire n_8_0_7133;
   wire n_8_0_7134;
   wire n_8_0_7135;
   wire n_8_0_7136;
   wire n_8_0_7137;
   wire n_8_0_7138;
   wire n_8_0_3615;
   wire n_8_0_7139;
   wire n_8_0_7140;
   wire n_8_0_3601;
   wire n_8_0_7141;
   wire n_8_0_7142;
   wire n_8_0_7143;
   wire n_8_0_3658;
   wire n_8_0_3659;
   wire n_8_0_7144;
   wire n_8_0_7145;
   wire n_8_0_7146;
   wire n_8_0_7147;
   wire n_8_0_3694;
   wire n_8_0_3682;
   wire n_8_0_3681;
   wire n_8_0_3687;
   wire n_8_0_3689;
   wire n_8_0_7148;
   wire n_8_0_3691;
   wire n_8_0_7149;
   wire n_8_0_4424;
   wire n_8_0_7150;
   wire n_8_0_7151;
   wire n_8_0_7152;
   wire n_8_0_3705;
   wire n_8_0_3702;
   wire n_8_0_3699;
   wire n_8_0_7153;
   wire n_8_0_7154;
   wire n_8_0_4503;
   wire n_8_0_6041;
   wire n_8_0_7155;
   wire n_8_0_4409;
   wire n_8_0_7156;
   wire n_8_0_7157;
   wire n_8_0_7158;
   wire n_8_0_7159;
   wire n_8_0_7160;
   wire n_8_0_7161;
   wire n_8_0_7162;
   wire n_8_0_3835;
   wire n_8_0_7163;
   wire n_8_0_7164;
   wire n_8_0_7165;
   wire n_8_0_7166;
   wire n_8_0_7167;
   wire n_8_0_7168;
   wire n_8_0_7169;
   wire n_8_0_7170;
   wire n_8_0_7171;
   wire n_8_0_3855;
   wire n_8_0_7172;
   wire n_8_0_7173;
   wire n_8_0_5674;
   wire n_8_0_7174;
   wire n_8_0_7175;
   wire n_8_0_7176;
   wire n_8_0_7177;
   wire n_8_0_7178;
   wire n_8_0_7179;
   wire n_8_0_5975;
   wire n_8_0_7180;
   wire n_8_0_7181;
   wire n_8_0_7182;
   wire n_8_0_4001;
   wire n_8_0_7183;
   wire n_8_0_7184;
   wire n_8_0_5954;
   wire n_8_0_7185;
   wire n_8_0_7186;
   wire n_8_0_7187;
   wire n_8_0_7188;
   wire n_8_0_7189;
   wire n_8_0_7190;
   wire n_8_0_4090;
   wire n_8_0_4096;
   wire n_8_0_4083;
   wire n_8_0_7191;
   wire n_8_0_7192;
   wire n_8_0_4598;
   wire n_8_0_4599;
   wire n_8_0_7193;
   wire n_8_0_7194;
   wire n_8_0_7195;
   wire n_8_0_7196;
   wire n_8_0_7197;
   wire n_8_0_7198;
   wire n_8_0_7199;
   wire n_8_0_7200;
   wire n_8_0_7201;
   wire n_8_0_7202;
   wire n_8_0_7203;
   wire n_8_0_7204;
   wire n_8_0_7205;
   wire n_8_0_7206;
   wire n_8_0_7207;
   wire n_8_0_7208;
   wire n_8_0_6118;
   wire n_8_0_7209;
   wire n_8_0_7210;
   wire n_8_0_7211;
   wire n_8_0_4363;
   wire n_8_0_7212;
   wire n_8_0_7213;
   wire n_8_0_4370;
   wire n_8_0_7214;
   wire n_8_0_7215;
   wire n_8_0_7216;
   wire n_8_0_7217;
   wire n_8_0_7218;
   wire n_8_0_7219;
   wire n_8_0_7220;
   wire n_8_0_7221;
   wire n_8_0_4532;
   wire n_8_0_7222;
   wire n_8_0_7223;
   wire n_8_0_7224;
   wire n_8_0_7225;
   wire n_8_0_7226;
   wire n_8_0_7227;
   wire n_8_0_7228;
   wire n_8_0_4465;
   wire n_8_0_7229;
   wire n_8_0_4471;
   wire n_8_0_4468;
   wire n_8_0_4595;
   wire n_8_0_7230;
   wire n_8_0_7231;
   wire n_8_0_7232;
   wire n_8_0_6465;
   wire n_8_0_6466;
   wire n_8_0_7233;
   wire n_8_0_6468;
   wire n_8_0_6467;
   wire n_8_0_7234;
   wire n_8_0_7235;
   wire n_8_0_7236;
   wire n_8_0_7237;
   wire n_8_0_7238;
   wire n_8_0_7239;
   wire n_8_0_7240;
   wire n_8_0_7241;
   wire n_8_0_7242;
   wire n_8_0_4618;
   wire n_8_0_4617;
   wire n_8_0_4619;
   wire n_8_0_4624;
   wire n_8_0_4623;
   wire n_8_0_4625;
   wire n_8_0_7243;
   wire n_8_0_7244;
   wire n_8_0_7245;
   wire n_8_0_7246;
   wire n_8_0_7247;
   wire n_8_0_7248;
   wire n_8_0_4827;
   wire n_8_0_4816;
   wire n_8_0_7249;
   wire n_8_0_4824;
   wire n_8_0_4820;
   wire n_8_0_7250;
   wire n_8_0_7251;
   wire n_8_0_7252;
   wire n_8_0_7253;
   wire n_8_0_7254;
   wire n_8_0_4823;
   wire n_8_0_7255;
   wire n_8_0_7256;
   wire n_8_0_7257;
   wire n_8_0_7258;
   wire n_8_0_4851;
   wire n_8_0_7259;
   wire n_8_0_7260;
   wire n_8_0_7261;
   wire n_8_0_4861;
   wire n_8_0_4864;
   wire n_8_0_4867;
   wire n_8_0_7262;
   wire n_8_0_4848;
   wire n_8_0_7263;
   wire n_8_0_7264;
   wire n_8_0_7265;
   wire n_8_0_5056;
   wire n_8_0_6362;
   wire n_8_0_7266;
   wire n_8_0_7267;
   wire n_8_0_7268;
   wire n_8_0_7269;
   wire n_8_0_7270;
   wire n_8_0_7271;
   wire n_8_0_7272;
   wire n_8_0_6054;
   wire n_8_0_7273;
   wire n_8_0_7274;
   wire n_8_0_7275;
   wire n_8_0_7276;
   wire n_8_0_5074;
   wire n_8_0_5077;
   wire n_8_0_5082;
   wire n_8_0_5065;
   wire n_8_0_7277;
   wire n_8_0_7278;
   wire n_8_0_5071;
   wire n_8_0_7279;
   wire n_8_0_7280;
   wire n_8_0_7281;
   wire n_8_0_5081;
   wire n_8_0_6042;
   wire n_8_0_6157;
   wire n_8_0_7282;
   wire n_8_0_7283;
   wire n_8_0_7284;
   wire n_8_0_7285;
   wire n_8_0_7286;
   wire n_8_0_7287;
   wire n_8_0_7288;
   wire n_8_0_5188;
   wire n_8_0_7289;
   wire n_8_0_7290;
   wire n_8_0_7291;
   wire n_8_0_7292;
   wire n_8_0_5178;
   wire n_8_0_5195;
   wire n_8_0_7293;
   wire n_8_0_7294;
   wire n_8_0_5176;
   wire n_8_0_7295;
   wire n_8_0_5182;
   wire n_8_0_5192;
   wire n_8_0_7296;
   wire n_8_0_5193;
   wire n_8_0_7297;
   wire n_8_0_7298;
   wire n_8_0_7299;
   wire n_8_0_7300;
   wire n_8_0_7301;
   wire n_8_0_7302;
   wire n_8_0_5365;
   wire n_8_0_7303;
   wire n_8_0_7304;
   wire n_8_0_7305;
   wire n_8_0_7306;
   wire n_8_0_5371;
   wire n_8_0_5377;
   wire n_8_0_7307;
   wire n_8_0_5480;
   wire n_8_0_7308;
   wire n_8_0_7309;
   wire n_8_0_7310;
   wire n_8_0_7311;
   wire n_8_0_7312;
   wire n_8_0_7313;
   wire n_8_0_7314;
   wire n_8_0_7315;
   wire n_8_0_7316;
   wire n_8_0_7317;
   wire n_8_0_7318;
   wire n_8_0_7319;
   wire n_8_0_5398;
   wire n_8_0_7320;
   wire n_8_0_7321;
   wire n_8_0_7322;
   wire n_8_0_5388;
   wire n_8_0_5407;
   wire n_8_0_7323;
   wire n_8_0_7324;
   wire n_8_0_7325;
   wire n_8_0_5403;
   wire n_8_0_5404;
   wire n_8_0_6540;
   wire n_8_0_7326;
   wire n_8_0_7327;
   wire n_8_0_7328;
   wire n_8_0_7329;
   wire n_8_0_7330;
   wire n_8_0_7331;
   wire n_8_0_7332;
   wire n_8_0_7333;
   wire n_8_0_6249;
   wire n_8_0_6593;
   wire n_8_0_6247;
   wire n_8_0_7334;
   wire n_8_0_7335;
   wire n_8_0_7336;
   wire n_8_0_5430;
   wire n_8_0_7337;
   wire n_8_0_7338;
   wire n_8_0_7339;
   wire n_8_0_7340;
   wire n_8_0_7341;
   wire n_8_0_7342;
   wire n_8_0_5414;
   wire n_8_0_5438;
   wire n_8_0_5416;
   wire n_8_0_5420;
   wire n_8_0_7343;
   wire n_8_0_5436;
   wire n_8_0_6724;
   wire n_8_0_6727;
   wire n_8_0_6233;
   wire n_8_0_6232;
   wire n_8_0_7344;
   wire n_8_0_7345;
   wire n_8_0_7346;
   wire n_8_0_7347;
   wire n_8_0_5985;
   wire n_8_0_7348;
   wire n_8_0_5993;
   wire n_8_0_7349;
   wire n_8_0_7350;
   wire n_8_0_7351;
   wire n_8_0_7352;
   wire n_8_0_7353;
   wire n_8_0_6752;
   wire n_8_0_7354;
   wire n_8_0_7355;
   wire n_8_0_7356;
   wire n_8_0_7357;
   wire n_8_0_7358;
   wire n_8_0_5973;
   wire n_8_0_7359;
   wire n_8_0_7360;
   wire n_8_0_7361;
   wire n_8_0_7362;
   wire n_8_0_7363;
   wire n_8_0_7364;
   wire n_8_0_7365;
   wire n_8_0_6595;
   wire n_8_0_7366;
   wire n_8_0_7367;
   wire n_8_0_6124;
   wire n_8_0_6129;
   wire n_8_0_7368;
   wire n_8_0_7369;
   wire n_8_0_7370;
   wire n_8_0_7371;
   wire n_8_0_6105;
   wire n_8_0_6110;
   wire n_8_0_6115;
   wire n_8_0_7372;
   wire n_8_0_6117;
   wire n_8_0_7373;
   wire n_8_0_7374;
   wire n_8_0_7375;
   wire n_8_0_7376;
   wire n_8_0_7377;
   wire n_8_0_6203;
   wire n_8_0_6179;
   wire n_8_0_6212;
   wire n_8_0_6186;
   wire n_8_0_7378;
   wire n_8_0_6207;
   wire n_8_0_6193;
   wire n_8_0_6199;
   wire n_8_0_7379;
   wire n_8_0_7380;
   wire n_8_0_7381;
   wire n_8_0_6729;
   wire n_8_0_7382;
   wire n_8_0_7383;
   wire n_8_0_7384;
   wire n_8_0_7385;
   wire n_8_0_7386;
   wire n_8_0_7387;
   wire n_8_0_7388;
   wire n_8_0_7389;
   wire n_8_0_7390;
   wire n_8_0_7391;
   wire n_8_0_7392;
   wire n_8_0_6811;
   wire n_8_0_7393;
   wire n_8_0_7394;
   wire n_8_0_7395;
   wire n_8_0_6280;
   wire n_8_0_6302;
   wire n_8_0_6272;
   wire n_8_0_6296;
   wire n_8_0_6289;
   wire n_8_0_7396;
   wire n_8_0_7397;
   wire n_8_0_7398;
   wire n_8_0_7399;
   wire n_8_0_7400;
   wire n_8_0_6279;
   wire n_8_0_7401;
   wire n_8_0_7402;
   wire n_8_0_6389;
   wire n_8_0_7403;
   wire n_8_0_7404;
   wire n_8_0_7405;
   wire n_8_0_7406;
   wire n_8_0_6396;
   wire n_8_0_7407;
   wire n_8_0_7408;
   wire n_8_0_7409;
   wire n_8_0_6378;
   wire n_8_0_7410;
   wire n_8_0_7411;
   wire n_8_0_7412;
   wire n_8_0_7413;
   wire n_8_0_6406;
   wire n_8_0_6383;
   wire n_8_0_6401;
   wire n_8_0_7414;
   wire n_8_0_7415;
   wire n_8_0_7416;
   wire n_8_0_6403;
   wire n_8_0_6715;
   wire n_8_0_7417;
   wire n_8_0_7418;
   wire n_8_0_7419;
   wire n_8_0_6602;
   wire n_8_0_6582;
   wire n_8_0_6755;
   wire n_8_0_6614;
   wire n_8_0_7420;
   wire n_8_0_6730;
   wire n_8_0_6731;
   wire n_8_0_7421;
   wire n_8_0_7422;
   wire n_8_0_7423;
   wire n_8_0_7424;
   wire n_8_0_7425;
   wire n_8_0_7426;
   wire n_8_0_7427;
   wire n_8_0_7428;
   wire n_8_0_6996;
   wire n_8_0_7429;
   wire n_8_0_6997;
   wire n_8_0_7003;
   wire n_8_0_7004;
   wire n_8_0_6998;
   wire n_8_0_6999;
   wire n_8_0_7000;
   wire n_8_0_7430;
   wire n_8_0_7431;
   wire n_8_0_7432;
   wire n_8_0_7433;
   wire n_8_0_7434;
   wire n_8_0_7435;
   wire n_8_0_6854;
   wire n_8_0_6853;
   wire n_8_0_7436;
   wire n_0_39;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_6;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire [6:0]buf_flush_i;
   wire n_0_170;
   wire n_0_296;
   wire [6:0]buf_fill_i;
   wire buf_is_empty;
   wire n_0_171;
   wire n_0_40;
   wire n_0_7;
   wire n_0_1_0;
   wire n_0_1_1;
   wire n_0_8;
   wire n_0_1_2;
   wire n_0_1_3;
   wire n_0_9;
   wire n_0_1_4;
   wire n_0_1_5;
   wire n_0_10;
   wire n_0_1_6;
   wire n_0_1_7;
   wire n_0_11;
   wire n_0_1_8;
   wire n_0_1_9;
   wire n_0_12;
   wire n_0_1_10;
   wire n_0_1_11;
   wire n_0_13;
   wire n_0_1_12;
   wire n_0_1_13;
   wire n_0_14;
   wire n_0_1_14;
   wire n_0_1_15;
   wire n_0_15;
   wire n_0_1_16;
   wire n_0_1_17;
   wire n_0_16;
   wire n_0_1_18;
   wire n_0_1_19;
   wire n_0_17;
   wire n_0_1_20;
   wire n_0_1_21;
   wire n_0_18;
   wire n_0_1_22;
   wire n_0_1_23;
   wire n_0_19;
   wire n_0_1_24;
   wire n_0_1_25;
   wire n_0_20;
   wire n_0_1_26;
   wire n_0_1_27;
   wire n_0_21;
   wire n_0_1_28;
   wire n_0_1_29;
   wire n_0_22;
   wire n_0_1_30;
   wire n_0_1_31;
   wire n_0_23;
   wire n_0_1_32;
   wire n_0_1_33;
   wire n_0_24;
   wire n_0_1_34;
   wire n_0_1_35;
   wire n_0_25;
   wire n_0_1_36;
   wire n_0_1_37;
   wire n_0_26;
   wire n_0_1_38;
   wire n_0_1_39;
   wire n_0_27;
   wire n_0_1_40;
   wire n_0_1_41;
   wire n_0_28;
   wire n_0_1_42;
   wire n_0_1_43;
   wire n_0_29;
   wire n_0_1_44;
   wire n_0_1_45;
   wire n_0_30;
   wire n_0_1_46;
   wire n_0_1_47;
   wire n_0_31;
   wire n_0_1_48;
   wire n_0_1_49;
   wire n_0_32;
   wire n_0_1_50;
   wire n_0_1_51;
   wire n_0_33;
   wire n_0_1_52;
   wire n_0_1_53;
   wire n_0_34;
   wire n_0_1_54;
   wire n_0_1_55;
   wire n_0_35;
   wire n_0_1_56;
   wire n_0_1_57;
   wire n_0_36;
   wire n_0_1_58;
   wire n_0_1_59;
   wire n_0_37;
   wire n_0_1_60;
   wire n_0_1_61;
   wire n_0_38;
   wire n_0_1_62;
   wire n_0_1_63;
   wire n_0_1_64;
   wire n_0_1_65;
   wire n_0_1_66;
   wire n_0_163;
   wire n_0_1_67;
   wire n_0_5;
   wire n_0_1_68;
   wire n_0_1_69;
   wire n_0_1_70;
   wire n_0_1_71;
   wire n_0_1_72;
   wire n_0_1_73;
   wire n_0_1_74;
   wire n_0_1_75;
   wire n_0_1_76;
   wire n_0_1_77;
   wire n_0_169;
   wire n_0_1_78;
   wire n_0_1_79;
   wire error_success_reg_enable_mux_n_0;
   wire n_0_164;
   wire n_0_295;
   wire n_0_294;
   wire n_0_293;
   wire n_0_292;
   wire n_0_291;
   wire n_0_290;
   wire n_0_289;
   wire n_0_288;
   wire n_0_287;
   wire n_0_286;
   wire n_0_285;
   wire n_0_284;
   wire n_0_283;
   wire n_0_282;
   wire n_0_281;
   wire n_0_280;
   wire n_0_279;
   wire n_0_278;
   wire n_0_277;
   wire n_0_276;
   wire n_0_275;
   wire n_0_274;
   wire n_0_273;
   wire n_0_272;
   wire n_0_271;
   wire n_0_270;
   wire n_0_269;
   wire n_0_268;
   wire n_0_267;
   wire n_0_266;
   wire n_0_265;
   wire n_0_264;
   wire n_0_263;
   wire n_0_262;
   wire n_0_261;
   wire n_0_260;
   wire n_0_259;
   wire n_0_258;
   wire n_0_257;
   wire n_0_256;
   wire n_0_255;
   wire n_0_254;
   wire n_0_253;
   wire n_0_252;
   wire n_0_251;
   wire n_0_250;
   wire n_0_249;
   wire n_0_248;
   wire n_0_247;
   wire n_0_246;
   wire n_0_245;
   wire n_0_244;
   wire n_0_243;
   wire n_0_242;
   wire n_0_241;
   wire n_0_240;
   wire n_0_239;
   wire n_0_238;
   wire n_0_237;
   wire n_0_236;
   wire n_0_235;
   wire n_0_234;
   wire n_0_233;
   wire n_0_232;
   wire n_0_231;
   wire n_0_230;
   wire n_0_229;
   wire n_0_228;
   wire n_0_227;
   wire n_0_226;
   wire n_0_225;
   wire n_0_224;
   wire n_0_222;
   wire n_0_221;
   wire n_0_220;
   wire n_0_219;
   wire n_0_218;
   wire n_0_217;
   wire n_0_216;
   wire n_0_215;
   wire n_0_214;
   wire n_0_213;
   wire n_0_212;
   wire n_0_211;
   wire n_0_210;
   wire n_0_209;
   wire n_0_208;
   wire n_0_207;
   wire n_0_206;
   wire n_0_205;
   wire n_0_204;
   wire n_0_203;
   wire n_0_202;
   wire n_0_201;
   wire n_0_200;
   wire n_0_199;
   wire n_0_198;
   wire n_0_197;
   wire n_0_196;
   wire n_0_195;
   wire n_0_194;
   wire n_0_193;
   wire n_0_192;
   wire n_0_191;
   wire n_0_190;
   wire n_0_189;
   wire n_0_188;
   wire n_0_187;
   wire n_0_186;
   wire n_0_185;
   wire n_0_184;
   wire n_0_183;
   wire n_0_182;
   wire n_0_181;
   wire n_0_180;
   wire n_0_179;
   wire n_0_178;
   wire n_0_177;
   wire n_0_176;
   wire n_0_175;
   wire n_0_174;
   wire n_0_173;
   wire n_0_172;
   wire n_0_168;
   wire n_0_167;
   wire n_0_166;
   wire n_0_165;
   wire n_0_223;
   wire n_0_0_0;
   wire n_0_0_1;
   wire [6:0]\out_bs[0] ;
   wire [6:0]\out_as[0] ;
   wire [6:0]buf_flush_i_inc;
   wire [6:0]buf_fill_flush_diff;
   wire [6:0]\out_bs[1] ;
   wire [6:0]\out_as[1] ;
   wire [6:0]\out_bs[2] ;
   wire [6:0]\out_as[2] ;
   wire [6:0]\out_bs[3] ;
   wire [6:0]\out_as[3] ;
   wire [6:0]\out_bs[4] ;
   wire [6:0]\out_as[4] ;
   wire [6:0]\out_bs[5] ;
   wire [6:0]\out_as[5] ;
   wire [6:0]\out_bs[6] ;
   wire [6:0]\out_as[6] ;
   wire [6:0]\out_bs[7] ;
   wire [6:0]\out_as[7] ;
   wire [6:0]buf_flush_i_inv;

   HA_X1 i_8_0_0 (.A(\out_as[0] [6]), .B(n_8_0_1165), .CO(n_8_0_5), .S());
   HA_X1 i_8_0_1 (.A(\out_as[0] [6]), .B(n_8_0_1164), .CO(n_8_0_4), .S());
   HA_X1 i_8_0_2 (.A(\out_as[0] [6]), .B(n_8_0_1162), .CO(n_8_0_0), .S());
   HA_X1 i_8_0_3 (.A(\out_as[0] [6]), .B(n_8_0_1166), .CO(n_8_0_3), .S());
   HA_X1 i_8_0_4 (.A(\out_as[0] [6]), .B(n_8_0_1243), .CO(n_8_0_1), .S());
   HA_X1 i_8_0_5 (.A(\out_as[0] [6]), .B(n_8_0_1161), .CO(n_8_0_2), .S());
   HA_X1 i_8_0_6 (.A(\out_as[0] [6]), .B(n_8_0_1160), .CO(n_8_0_6), .S());
   HA_X1 i_8_0_7 (.A(\out_as[0] [6]), .B(n_8_0_1294), .CO(n_8_0_7), .S());
   HA_X1 i_8_0_8 (.A(\out_as[0] [6]), .B(n_8_0_1302), .CO(n_8_0_8), .S());
   HA_X1 i_8_0_9 (.A(\out_as[0] [6]), .B(n_8_0_1159), .CO(n_8_0_9), .S());
   HA_X1 i_8_0_10 (.A(\out_as[0] [6]), .B(n_8_0_1158), .CO(n_8_0_10), .S());
   HA_X1 i_8_0_11 (.A(\out_as[0] [6]), .B(n_8_0_1157), .CO(n_8_0_11), .S());
   HA_X1 i_8_0_12 (.A(\out_as[0] [6]), .B(n_8_0_1156), .CO(n_8_0_12), .S());
   HA_X1 i_8_0_13 (.A(\out_as[0] [6]), .B(n_8_0_1155), .CO(n_8_0_13), .S());
   HA_X1 i_8_0_14 (.A(\out_as[0] [6]), .B(n_8_0_1154), .CO(n_8_0_14), .S());
   HA_X1 i_8_0_15 (.A(\out_as[0] [6]), .B(n_8_0_1359), .CO(n_8_0_15), .S());
   HA_X1 i_8_0_16 (.A(\out_as[0] [6]), .B(n_8_0_1153), .CO(n_8_0_16), .S());
   HA_X1 i_8_0_17 (.A(\out_as[0] [6]), .B(n_8_0_1368), .CO(n_8_0_17), .S());
   HA_X1 i_8_0_18 (.A(\out_as[0] [6]), .B(n_8_0_1152), .CO(n_8_0_18), .S());
   HA_X1 i_8_0_19 (.A(\out_as[0] [6]), .B(n_8_0_1377), .CO(n_8_0_19), .S());
   HA_X1 i_8_0_20 (.A(\out_as[0] [6]), .B(n_8_0_1378), .CO(n_8_0_20), .S());
   HA_X1 i_8_0_21 (.A(\out_as[0] [6]), .B(n_8_0_1151), .CO(n_8_0_21), .S());
   HA_X1 i_8_0_22 (.A(\out_as[0] [6]), .B(n_8_0_1150), .CO(n_8_0_22), .S());
   HA_X1 i_8_0_23 (.A(\out_as[0] [6]), .B(n_8_0_1149), .CO(n_8_0_23), .S());
   HA_X1 i_8_0_24 (.A(\out_as[0] [6]), .B(n_8_0_1148), .CO(n_8_0_24), .S());
   HA_X1 i_8_0_25 (.A(\out_as[0] [6]), .B(n_8_0_1147), .CO(n_8_0_25), .S());
   HA_X1 i_8_0_26 (.A(\out_as[0] [6]), .B(n_8_0_1396), .CO(n_8_0_26), .S());
   HA_X1 i_8_0_27 (.A(\out_as[0] [6]), .B(n_8_0_1146), .CO(n_8_0_27), .S());
   HA_X1 i_8_0_28 (.A(\out_as[0] [6]), .B(n_8_0_1406), .CO(n_8_0_28), .S());
   HA_X1 i_8_0_29 (.A(\out_as[0] [6]), .B(n_8_0_1145), .CO(n_8_0_29), .S());
   HA_X1 i_8_0_30 (.A(\out_as[0] [6]), .B(n_8_0_1144), .CO(n_8_0_30), .S());
   HA_X1 i_8_0_31 (.A(\out_as[0] [6]), .B(\out_as[0] [5]), .CO(n_8_0_31), .S());
   HA_X1 i_8_0_32 (.A(\out_as[0] [6]), .B(n_8_0_959), .CO(n_8_0_32), .S());
   HA_X1 i_8_0_33 (.A(\out_as[0] [6]), .B(n_8_0_951), .CO(n_8_0_33), .S());
   HA_X1 i_8_0_34 (.A(\out_as[0] [6]), .B(n_8_0_943), .CO(n_8_0_34), .S());
   HA_X1 i_8_0_35 (.A(\out_as[0] [6]), .B(n_8_0_935), .CO(n_8_0_35), .S());
   HA_X1 i_8_0_36 (.A(\out_as[0] [6]), .B(n_8_0_927), .CO(n_8_0_36), .S());
   HA_X1 i_8_0_37 (.A(\out_as[0] [6]), .B(n_8_0_919), .CO(n_8_0_37), .S());
   HA_X1 i_8_0_38 (.A(\out_as[0] [6]), .B(n_8_0_911), .CO(n_8_0_38), .S());
   HA_X1 i_8_0_39 (.A(\out_as[0] [6]), .B(n_8_0_903), .CO(n_8_0_39), .S());
   HA_X1 i_8_0_40 (.A(\out_as[0] [6]), .B(n_8_0_895), .CO(n_8_0_40), .S());
   HA_X1 i_8_0_41 (.A(\out_as[0] [6]), .B(n_8_0_887), .CO(n_8_0_41), .S());
   HA_X1 i_8_0_42 (.A(\out_as[0] [6]), .B(n_8_0_879), .CO(n_8_0_42), .S());
   HA_X1 i_8_0_43 (.A(\out_as[0] [6]), .B(n_8_0_871), .CO(n_8_0_43), .S());
   HA_X1 i_8_0_44 (.A(\out_as[0] [6]), .B(n_8_0_863), .CO(n_8_0_44), .S());
   HA_X1 i_8_0_45 (.A(\out_as[0] [6]), .B(n_8_0_855), .CO(n_8_0_45), .S());
   HA_X1 i_8_0_46 (.A(\out_as[0] [6]), .B(n_8_0_847), .CO(n_8_0_46), .S());
   HA_X1 i_8_0_47 (.A(\out_as[0] [6]), .B(n_8_0_839), .CO(n_8_0_47), .S());
   HA_X1 i_8_0_48 (.A(\out_as[0] [6]), .B(n_8_0_831), .CO(n_8_0_48), .S());
   HA_X1 i_8_0_49 (.A(\out_as[0] [6]), .B(n_8_0_815), .CO(n_8_0_49), .S());
   HA_X1 i_8_0_50 (.A(\out_as[0] [6]), .B(n_8_0_799), .CO(n_8_0_50), .S());
   HA_X1 i_8_0_51 (.A(\out_as[0] [6]), .B(n_8_0_783), .CO(n_8_0_51), .S());
   HA_X1 i_8_0_52 (.A(\out_as[0] [6]), .B(n_8_0_767), .CO(n_8_0_52), .S());
   HA_X1 i_8_0_53 (.A(\out_as[0] [6]), .B(n_8_0_751), .CO(n_8_0_53), .S());
   HA_X1 i_8_0_54 (.A(\out_as[0] [6]), .B(n_8_0_735), .CO(n_8_0_54), .S());
   HA_X1 i_8_0_55 (.A(\out_as[0] [6]), .B(n_8_0_719), .CO(n_8_0_55), .S());
   HA_X1 i_8_0_56 (.A(\out_as[0] [6]), .B(n_8_0_703), .CO(n_8_0_56), .S());
   HA_X1 i_8_0_57 (.A(\out_as[0] [6]), .B(n_8_0_679), .CO(n_8_0_57), .S());
   HA_X1 i_8_0_58 (.A(\out_as[0] [6]), .B(n_8_0_655), .CO(n_8_0_58), .S());
   HA_X1 i_8_0_59 (.A(\out_as[0] [6]), .B(n_8_0_631), .CO(n_8_0_59), .S());
   HA_X1 i_8_0_60 (.A(\out_as[0] [6]), .B(n_8_0_607), .CO(n_8_0_60), .S());
   HA_X1 i_8_0_61 (.A(\out_as[0] [6]), .B(n_8_0_575), .CO(n_8_0_61), .S());
   HA_X1 i_8_0_62 (.A(\out_as[0] [6]), .B(n_8_0_543), .CO(n_8_0_62), .S());
   HA_X1 i_8_0_63 (.A(\out_as[1] [6]), .B(n_8_0_1141), .CO(n_8_0_63), .S());
   HA_X1 i_8_0_64 (.A(\out_as[1] [6]), .B(n_8_0_1142), .CO(n_8_0_64), .S());
   HA_X1 i_8_0_65 (.A(\out_as[1] [6]), .B(n_8_0_1138), .CO(n_8_0_65), .S());
   HA_X1 i_8_0_66 (.A(\out_as[1] [6]), .B(n_8_0_1229), .CO(n_8_0_66), .S());
   HA_X1 i_8_0_67 (.A(\out_as[1] [6]), .B(n_8_0_1136), .CO(n_8_0_67), .S());
   HA_X1 i_8_0_68 (.A(\out_as[1] [6]), .B(n_8_0_1265), .CO(n_8_0_68), .S());
   HA_X1 i_8_0_69 (.A(\out_as[1] [6]), .B(n_8_0_1279), .CO(n_8_0_69), .S());
   HA_X1 i_8_0_70 (.A(\out_as[1] [6]), .B(n_8_0_1230), .CO(n_8_0_70), .S());
   HA_X1 i_8_0_71 (.A(\out_as[1] [6]), .B(n_8_0_1135), .CO(n_8_0_71), .S());
   HA_X1 i_8_0_72 (.A(\out_as[1] [6]), .B(n_8_0_1134), .CO(n_8_0_72), .S());
   HA_X1 i_8_0_73 (.A(\out_as[1] [6]), .B(n_8_0_1133), .CO(n_8_0_73), .S());
   HA_X1 i_8_0_74 (.A(\out_as[1] [6]), .B(n_8_0_1132), .CO(n_8_0_74), .S());
   HA_X1 i_8_0_75 (.A(\out_as[1] [6]), .B(n_8_0_1131), .CO(n_8_0_75), .S());
   HA_X1 i_8_0_76 (.A(\out_as[1] [6]), .B(n_8_0_1130), .CO(n_8_0_76), .S());
   HA_X1 i_8_0_77 (.A(\out_as[1] [6]), .B(n_8_0_1129), .CO(n_8_0_77), .S());
   HA_X1 i_8_0_78 (.A(\out_as[1] [6]), .B(n_8_0_1356), .CO(n_8_0_78), .S());
   HA_X1 i_8_0_79 (.A(\out_as[1] [6]), .B(n_8_0_1361), .CO(n_8_0_79), .S());
   HA_X1 i_8_0_80 (.A(\out_as[1] [6]), .B(n_8_0_1369), .CO(n_8_0_80), .S());
   HA_X1 i_8_0_81 (.A(\out_as[1] [6]), .B(n_8_0_1373), .CO(n_8_0_81), .S());
   HA_X1 i_8_0_82 (.A(\out_as[1] [6]), .B(n_8_0_1376), .CO(n_8_0_82), .S());
   HA_X1 i_8_0_83 (.A(\out_as[1] [6]), .B(n_8_0_1128), .CO(n_8_0_83), .S());
   HA_X1 i_8_0_84 (.A(\out_as[1] [6]), .B(n_8_0_1380), .CO(n_8_0_84), .S());
   HA_X1 i_8_0_85 (.A(\out_as[1] [6]), .B(n_8_0_1383), .CO(n_8_0_85), .S());
   HA_X1 i_8_0_86 (.A(\out_as[1] [6]), .B(n_8_0_1127), .CO(n_8_0_86), .S());
   HA_X1 i_8_0_87 (.A(\out_as[1] [6]), .B(n_8_0_1388), .CO(n_8_0_87), .S());
   HA_X1 i_8_0_88 (.A(\out_as[1] [6]), .B(n_8_0_1126), .CO(n_8_0_88), .S());
   HA_X1 i_8_0_89 (.A(\out_as[1] [6]), .B(n_8_0_1125), .CO(n_8_0_89), .S());
   HA_X1 i_8_0_90 (.A(\out_as[1] [6]), .B(n_8_0_1398), .CO(n_8_0_90), .S());
   HA_X1 i_8_0_91 (.A(\out_as[1] [6]), .B(n_8_0_1402), .CO(n_8_0_91), .S());
   HA_X1 i_8_0_92 (.A(\out_as[1] [6]), .B(n_8_0_1124), .CO(n_8_0_92), .S());
   HA_X1 i_8_0_93 (.A(\out_as[1] [6]), .B(n_8_0_1412), .CO(n_8_0_93), .S());
   HA_X1 i_8_0_94 (.A(\out_as[1] [6]), .B(\out_as[1] [5]), .CO(n_8_0_94), .S());
   HA_X1 i_8_0_95 (.A(\out_as[1] [6]), .B(n_8_0_958), .CO(n_8_0_95), .S());
   HA_X1 i_8_0_96 (.A(\out_as[1] [6]), .B(n_8_0_950), .CO(n_8_0_96), .S());
   HA_X1 i_8_0_97 (.A(\out_as[1] [6]), .B(n_8_0_942), .CO(n_8_0_97), .S());
   HA_X1 i_8_0_98 (.A(\out_as[1] [6]), .B(n_8_0_934), .CO(n_8_0_98), .S());
   HA_X1 i_8_0_99 (.A(\out_as[1] [6]), .B(n_8_0_926), .CO(n_8_0_99), .S());
   HA_X1 i_8_0_100 (.A(\out_as[1] [6]), .B(n_8_0_918), .CO(n_8_0_100), .S());
   HA_X1 i_8_0_101 (.A(\out_as[1] [6]), .B(n_8_0_910), .CO(n_8_0_101), .S());
   HA_X1 i_8_0_102 (.A(\out_as[1] [6]), .B(n_8_0_902), .CO(n_8_0_102), .S());
   HA_X1 i_8_0_103 (.A(\out_as[1] [6]), .B(n_8_0_894), .CO(n_8_0_103), .S());
   HA_X1 i_8_0_104 (.A(\out_as[1] [6]), .B(n_8_0_886), .CO(n_8_0_104), .S());
   HA_X1 i_8_0_105 (.A(\out_as[1] [6]), .B(n_8_0_878), .CO(n_8_0_105), .S());
   HA_X1 i_8_0_106 (.A(\out_as[1] [6]), .B(n_8_0_870), .CO(n_8_0_106), .S());
   HA_X1 i_8_0_107 (.A(\out_as[1] [6]), .B(n_8_0_862), .CO(n_8_0_107), .S());
   HA_X1 i_8_0_108 (.A(\out_as[1] [6]), .B(n_8_0_854), .CO(n_8_0_108), .S());
   HA_X1 i_8_0_109 (.A(\out_as[1] [6]), .B(n_8_0_846), .CO(n_8_0_109), .S());
   HA_X1 i_8_0_110 (.A(\out_as[1] [6]), .B(n_8_0_838), .CO(n_8_0_110), .S());
   HA_X1 i_8_0_111 (.A(\out_as[1] [6]), .B(n_8_0_829), .CO(n_8_0_111), .S());
   HA_X1 i_8_0_112 (.A(\out_as[1] [6]), .B(n_8_0_813), .CO(n_8_0_112), .S());
   HA_X1 i_8_0_113 (.A(\out_as[1] [6]), .B(n_8_0_797), .CO(n_8_0_113), .S());
   HA_X1 i_8_0_114 (.A(\out_as[1] [6]), .B(n_8_0_781), .CO(n_8_0_114), .S());
   HA_X1 i_8_0_115 (.A(\out_as[1] [6]), .B(n_8_0_765), .CO(n_8_0_115), .S());
   HA_X1 i_8_0_116 (.A(\out_as[1] [6]), .B(n_8_0_749), .CO(n_8_0_116), .S());
   HA_X1 i_8_0_117 (.A(\out_as[1] [6]), .B(n_8_0_733), .CO(n_8_0_117), .S());
   HA_X1 i_8_0_118 (.A(\out_as[1] [6]), .B(n_8_0_717), .CO(n_8_0_118), .S());
   HA_X1 i_8_0_119 (.A(\out_as[1] [6]), .B(n_8_0_700), .CO(n_8_0_119), .S());
   HA_X1 i_8_0_120 (.A(\out_as[1] [6]), .B(n_8_0_676), .CO(n_8_0_120), .S());
   HA_X1 i_8_0_121 (.A(\out_as[1] [6]), .B(n_8_0_652), .CO(n_8_0_121), .S());
   HA_X1 i_8_0_122 (.A(\out_as[1] [6]), .B(n_8_0_628), .CO(n_8_0_122), .S());
   HA_X1 i_8_0_123 (.A(\out_as[1] [6]), .B(n_8_0_603), .CO(n_8_0_123), .S());
   HA_X1 i_8_0_124 (.A(\out_as[1] [6]), .B(n_8_0_571), .CO(n_8_0_124), .S());
   HA_X1 i_8_0_125 (.A(\out_as[1] [6]), .B(n_8_0_538), .CO(n_8_0_125), .S());
   HA_X1 i_8_0_126 (.A(\out_as[2] [6]), .B(n_8_0_1123), .CO(n_8_0_126), .S());
   HA_X1 i_8_0_127 (.A(\out_as[2] [6]), .B(n_8_0_1120), .CO(n_8_0_127), .S());
   HA_X1 i_8_0_128 (.A(\out_as[2] [6]), .B(n_8_0_1117), .CO(n_8_0_128), .S());
   HA_X1 i_8_0_129 (.A(\out_as[2] [6]), .B(n_8_0_1222), .CO(n_8_0_129), .S());
   HA_X1 i_8_0_130 (.A(\out_as[2] [6]), .B(n_8_0_1115), .CO(n_8_0_130), .S());
   HA_X1 i_8_0_131 (.A(\out_as[2] [6]), .B(n_8_0_1114), .CO(n_8_0_131), .S());
   HA_X1 i_8_0_132 (.A(\out_as[2] [6]), .B(n_8_0_1282), .CO(n_8_0_132), .S());
   HA_X1 i_8_0_133 (.A(\out_as[2] [6]), .B(n_8_0_1121), .CO(n_8_0_133), .S());
   HA_X1 i_8_0_134 (.A(\out_as[2] [6]), .B(n_8_0_1113), .CO(n_8_0_134), .S());
   HA_X1 i_8_0_135 (.A(\out_as[2] [6]), .B(n_8_0_1112), .CO(n_8_0_135), .S());
   HA_X1 i_8_0_136 (.A(\out_as[2] [6]), .B(n_8_0_1111), .CO(n_8_0_136), .S());
   HA_X1 i_8_0_137 (.A(\out_as[2] [6]), .B(n_8_0_1325), .CO(n_8_0_137), .S());
   HA_X1 i_8_0_138 (.A(\out_as[2] [6]), .B(n_8_0_1110), .CO(n_8_0_138), .S());
   HA_X1 i_8_0_139 (.A(\out_as[2] [6]), .B(n_8_0_1109), .CO(n_8_0_139), .S());
   HA_X1 i_8_0_140 (.A(\out_as[2] [6]), .B(n_8_0_1108), .CO(n_8_0_140), .S());
   HA_X1 i_8_0_141 (.A(\out_as[2] [6]), .B(n_8_0_1355), .CO(n_8_0_141), .S());
   HA_X1 i_8_0_142 (.A(\out_as[2] [6]), .B(n_8_0_1364), .CO(n_8_0_142), .S());
   HA_X1 i_8_0_143 (.A(\out_as[2] [6]), .B(n_8_0_1370), .CO(n_8_0_143), .S());
   HA_X1 i_8_0_144 (.A(\out_as[2] [6]), .B(n_8_0_1374), .CO(n_8_0_144), .S());
   HA_X1 i_8_0_145 (.A(\out_as[2] [6]), .B(n_8_0_1107), .CO(n_8_0_145), .S());
   HA_X1 i_8_0_146 (.A(\out_as[2] [6]), .B(n_8_0_1106), .CO(n_8_0_146), .S());
   HA_X1 i_8_0_147 (.A(\out_as[2] [6]), .B(n_8_0_1105), .CO(n_8_0_147), .S());
   HA_X1 i_8_0_148 (.A(\out_as[2] [6]), .B(n_8_0_1382), .CO(n_8_0_148), .S());
   HA_X1 i_8_0_149 (.A(\out_as[2] [6]), .B(n_8_0_1385), .CO(n_8_0_149), .S());
   HA_X1 i_8_0_150 (.A(\out_as[2] [6]), .B(n_8_0_1390), .CO(n_8_0_150), .S());
   HA_X1 i_8_0_151 (.A(\out_as[2] [6]), .B(n_8_0_1104), .CO(n_8_0_151), .S());
   HA_X1 i_8_0_152 (.A(\out_as[2] [6]), .B(n_8_0_1103), .CO(n_8_0_152), .S());
   HA_X1 i_8_0_153 (.A(\out_as[2] [6]), .B(n_8_0_1102), .CO(n_8_0_153), .S());
   HA_X1 i_8_0_154 (.A(\out_as[2] [6]), .B(n_8_0_1101), .CO(n_8_0_154), .S());
   HA_X1 i_8_0_155 (.A(\out_as[2] [6]), .B(n_8_0_1100), .CO(n_8_0_155), .S());
   HA_X1 i_8_0_156 (.A(\out_as[2] [6]), .B(n_8_0_1413), .CO(n_8_0_156), .S());
   HA_X1 i_8_0_157 (.A(\out_as[2] [6]), .B(\out_as[2] [5]), .CO(n_8_0_157), 
      .S());
   HA_X1 i_8_0_158 (.A(\out_as[2] [6]), .B(n_8_0_957), .CO(n_8_0_158), .S());
   HA_X1 i_8_0_159 (.A(\out_as[2] [6]), .B(n_8_0_949), .CO(n_8_0_159), .S());
   HA_X1 i_8_0_160 (.A(\out_as[2] [6]), .B(n_8_0_941), .CO(n_8_0_160), .S());
   HA_X1 i_8_0_161 (.A(\out_as[2] [6]), .B(n_8_0_933), .CO(n_8_0_161), .S());
   HA_X1 i_8_0_162 (.A(\out_as[2] [6]), .B(n_8_0_925), .CO(n_8_0_162), .S());
   HA_X1 i_8_0_163 (.A(\out_as[2] [6]), .B(n_8_0_917), .CO(n_8_0_163), .S());
   HA_X1 i_8_0_164 (.A(\out_as[2] [6]), .B(n_8_0_909), .CO(n_8_0_164), .S());
   HA_X1 i_8_0_165 (.A(\out_as[2] [6]), .B(n_8_0_901), .CO(n_8_0_165), .S());
   HA_X1 i_8_0_166 (.A(\out_as[2] [6]), .B(n_8_0_893), .CO(n_8_0_166), .S());
   HA_X1 i_8_0_167 (.A(\out_as[2] [6]), .B(n_8_0_885), .CO(n_8_0_167), .S());
   HA_X1 i_8_0_168 (.A(\out_as[2] [6]), .B(n_8_0_877), .CO(n_8_0_168), .S());
   HA_X1 i_8_0_169 (.A(\out_as[2] [6]), .B(n_8_0_869), .CO(n_8_0_169), .S());
   HA_X1 i_8_0_170 (.A(\out_as[2] [6]), .B(n_8_0_861), .CO(n_8_0_170), .S());
   HA_X1 i_8_0_171 (.A(\out_as[2] [6]), .B(n_8_0_853), .CO(n_8_0_171), .S());
   HA_X1 i_8_0_172 (.A(\out_as[2] [6]), .B(n_8_0_845), .CO(n_8_0_172), .S());
   HA_X1 i_8_0_173 (.A(\out_as[2] [6]), .B(n_8_0_837), .CO(n_8_0_173), .S());
   HA_X1 i_8_0_174 (.A(\out_as[2] [6]), .B(n_8_0_827), .CO(n_8_0_174), .S());
   HA_X1 i_8_0_175 (.A(\out_as[2] [6]), .B(n_8_0_811), .CO(n_8_0_175), .S());
   HA_X1 i_8_0_176 (.A(\out_as[2] [6]), .B(n_8_0_795), .CO(n_8_0_176), .S());
   HA_X1 i_8_0_177 (.A(\out_as[2] [6]), .B(n_8_0_779), .CO(n_8_0_177), .S());
   HA_X1 i_8_0_178 (.A(\out_as[2] [6]), .B(n_8_0_763), .CO(n_8_0_178), .S());
   HA_X1 i_8_0_179 (.A(\out_as[2] [6]), .B(n_8_0_747), .CO(n_8_0_179), .S());
   HA_X1 i_8_0_180 (.A(\out_as[2] [6]), .B(n_8_0_731), .CO(n_8_0_180), .S());
   HA_X1 i_8_0_181 (.A(\out_as[2] [6]), .B(n_8_0_715), .CO(n_8_0_181), .S());
   HA_X1 i_8_0_182 (.A(\out_as[2] [6]), .B(n_8_0_697), .CO(n_8_0_182), .S());
   HA_X1 i_8_0_183 (.A(\out_as[2] [6]), .B(n_8_0_673), .CO(n_8_0_183), .S());
   HA_X1 i_8_0_184 (.A(\out_as[2] [6]), .B(n_8_0_649), .CO(n_8_0_184), .S());
   HA_X1 i_8_0_185 (.A(\out_as[2] [6]), .B(n_8_0_625), .CO(n_8_0_185), .S());
   HA_X1 i_8_0_186 (.A(\out_as[2] [6]), .B(n_8_0_599), .CO(n_8_0_186), .S());
   HA_X1 i_8_0_187 (.A(\out_as[2] [6]), .B(n_8_0_567), .CO(n_8_0_187), .S());
   HA_X1 i_8_0_188 (.A(\out_as[2] [6]), .B(n_8_0_533), .CO(n_8_0_188), .S());
   HA_X1 i_8_0_189 (.A(\out_as[3] [6]), .B(n_8_0_1097), .CO(n_8_0_189), .S());
   HA_X1 i_8_0_190 (.A(\out_as[3] [6]), .B(n_8_0_1095), .CO(n_8_0_190), .S());
   HA_X1 i_8_0_191 (.A(\out_as[3] [6]), .B(n_8_0_1093), .CO(n_8_0_191), .S());
   HA_X1 i_8_0_192 (.A(\out_as[3] [6]), .B(n_8_0_1092), .CO(n_8_0_192), .S());
   HA_X1 i_8_0_193 (.A(\out_as[3] [6]), .B(n_8_0_1248), .CO(n_8_0_193), .S());
   HA_X1 i_8_0_194 (.A(\out_as[3] [6]), .B(n_8_0_1253), .CO(n_8_0_194), .S());
   HA_X1 i_8_0_195 (.A(\out_as[3] [6]), .B(n_8_0_1091), .CO(n_8_0_195), .S());
   HA_X1 i_8_0_196 (.A(\out_as[3] [6]), .B(n_8_0_1254), .CO(n_8_0_196), .S());
   HA_X1 i_8_0_197 (.A(\out_as[3] [6]), .B(n_8_0_1300), .CO(n_8_0_197), .S());
   HA_X1 i_8_0_198 (.A(\out_as[3] [6]), .B(n_8_0_1090), .CO(n_8_0_198), .S());
   HA_X1 i_8_0_199 (.A(\out_as[3] [6]), .B(n_8_0_1089), .CO(n_8_0_199), .S());
   HA_X1 i_8_0_200 (.A(\out_as[3] [6]), .B(n_8_0_1088), .CO(n_8_0_200), .S());
   HA_X1 i_8_0_201 (.A(\out_as[3] [6]), .B(n_8_0_1087), .CO(n_8_0_201), .S());
   HA_X1 i_8_0_202 (.A(\out_as[3] [6]), .B(n_8_0_1086), .CO(n_8_0_202), .S());
   HA_X1 i_8_0_203 (.A(\out_as[3] [6]), .B(n_8_0_1085), .CO(n_8_0_203), .S());
   HA_X1 i_8_0_204 (.A(\out_as[3] [6]), .B(n_8_0_1353), .CO(n_8_0_204), .S());
   HA_X1 i_8_0_205 (.A(\out_as[3] [6]), .B(n_8_0_1363), .CO(n_8_0_205), .S());
   HA_X1 i_8_0_206 (.A(\out_as[3] [6]), .B(n_8_0_1084), .CO(n_8_0_206), .S());
   HA_X1 i_8_0_207 (.A(\out_as[3] [6]), .B(n_8_0_1083), .CO(n_8_0_207), .S());
   HA_X1 i_8_0_208 (.A(\out_as[3] [6]), .B(n_8_0_1082), .CO(n_8_0_208), .S());
   HA_X1 i_8_0_209 (.A(\out_as[3] [6]), .B(n_8_0_1081), .CO(n_8_0_209), .S());
   HA_X1 i_8_0_210 (.A(\out_as[3] [6]), .B(n_8_0_1080), .CO(n_8_0_210), .S());
   HA_X1 i_8_0_211 (.A(\out_as[3] [6]), .B(n_8_0_1079), .CO(n_8_0_211), .S());
   HA_X1 i_8_0_212 (.A(\out_as[3] [6]), .B(n_8_0_1387), .CO(n_8_0_212), .S());
   HA_X1 i_8_0_213 (.A(\out_as[3] [6]), .B(n_8_0_1078), .CO(n_8_0_213), .S());
   HA_X1 i_8_0_214 (.A(\out_as[3] [6]), .B(n_8_0_1077), .CO(n_8_0_214), .S());
   HA_X1 i_8_0_215 (.A(\out_as[3] [6]), .B(n_8_0_1076), .CO(n_8_0_215), .S());
   HA_X1 i_8_0_216 (.A(\out_as[3] [6]), .B(n_8_0_1400), .CO(n_8_0_216), .S());
   HA_X1 i_8_0_217 (.A(\out_as[3] [6]), .B(n_8_0_1407), .CO(n_8_0_217), .S());
   HA_X1 i_8_0_218 (.A(\out_as[3] [6]), .B(n_8_0_1410), .CO(n_8_0_218), .S());
   HA_X1 i_8_0_219 (.A(\out_as[3] [6]), .B(n_8_0_1075), .CO(n_8_0_219), .S());
   HA_X1 i_8_0_220 (.A(\out_as[3] [6]), .B(\out_as[3] [5]), .CO(n_8_0_220), 
      .S());
   HA_X1 i_8_0_221 (.A(\out_as[3] [6]), .B(n_8_0_956), .CO(n_8_0_221), .S());
   HA_X1 i_8_0_222 (.A(\out_as[3] [6]), .B(n_8_0_948), .CO(n_8_0_222), .S());
   HA_X1 i_8_0_223 (.A(\out_as[3] [6]), .B(n_8_0_940), .CO(n_8_0_223), .S());
   HA_X1 i_8_0_224 (.A(\out_as[3] [6]), .B(n_8_0_932), .CO(n_8_0_224), .S());
   HA_X1 i_8_0_225 (.A(\out_as[3] [6]), .B(n_8_0_924), .CO(n_8_0_225), .S());
   HA_X1 i_8_0_226 (.A(\out_as[3] [6]), .B(n_8_0_916), .CO(n_8_0_226), .S());
   HA_X1 i_8_0_227 (.A(\out_as[3] [6]), .B(n_8_0_908), .CO(n_8_0_227), .S());
   HA_X1 i_8_0_228 (.A(\out_as[3] [6]), .B(n_8_0_900), .CO(n_8_0_228), .S());
   HA_X1 i_8_0_229 (.A(\out_as[3] [6]), .B(n_8_0_892), .CO(n_8_0_229), .S());
   HA_X1 i_8_0_230 (.A(\out_as[3] [6]), .B(n_8_0_884), .CO(n_8_0_230), .S());
   HA_X1 i_8_0_231 (.A(\out_as[3] [6]), .B(n_8_0_876), .CO(n_8_0_231), .S());
   HA_X1 i_8_0_232 (.A(\out_as[3] [6]), .B(n_8_0_868), .CO(n_8_0_232), .S());
   HA_X1 i_8_0_233 (.A(\out_as[3] [6]), .B(n_8_0_860), .CO(n_8_0_233), .S());
   HA_X1 i_8_0_234 (.A(\out_as[3] [6]), .B(n_8_0_852), .CO(n_8_0_234), .S());
   HA_X1 i_8_0_235 (.A(\out_as[3] [6]), .B(n_8_0_844), .CO(n_8_0_235), .S());
   HA_X1 i_8_0_236 (.A(\out_as[3] [6]), .B(n_8_0_836), .CO(n_8_0_236), .S());
   HA_X1 i_8_0_237 (.A(\out_as[3] [6]), .B(n_8_0_825), .CO(n_8_0_237), .S());
   HA_X1 i_8_0_238 (.A(\out_as[3] [6]), .B(n_8_0_809), .CO(n_8_0_238), .S());
   HA_X1 i_8_0_239 (.A(\out_as[3] [6]), .B(n_8_0_793), .CO(n_8_0_239), .S());
   HA_X1 i_8_0_240 (.A(\out_as[3] [6]), .B(n_8_0_777), .CO(n_8_0_240), .S());
   HA_X1 i_8_0_241 (.A(\out_as[3] [6]), .B(n_8_0_761), .CO(n_8_0_241), .S());
   HA_X1 i_8_0_242 (.A(\out_as[3] [6]), .B(n_8_0_745), .CO(n_8_0_242), .S());
   HA_X1 i_8_0_243 (.A(\out_as[3] [6]), .B(n_8_0_729), .CO(n_8_0_243), .S());
   HA_X1 i_8_0_244 (.A(\out_as[3] [6]), .B(n_8_0_713), .CO(n_8_0_244), .S());
   HA_X1 i_8_0_245 (.A(\out_as[3] [6]), .B(n_8_0_694), .CO(n_8_0_245), .S());
   HA_X1 i_8_0_246 (.A(\out_as[3] [6]), .B(n_8_0_670), .CO(n_8_0_246), .S());
   HA_X1 i_8_0_247 (.A(\out_as[3] [6]), .B(n_8_0_646), .CO(n_8_0_247), .S());
   HA_X1 i_8_0_248 (.A(\out_as[3] [6]), .B(n_8_0_622), .CO(n_8_0_248), .S());
   HA_X1 i_8_0_249 (.A(\out_as[3] [6]), .B(n_8_0_595), .CO(n_8_0_249), .S());
   HA_X1 i_8_0_250 (.A(\out_as[3] [6]), .B(n_8_0_563), .CO(n_8_0_250), .S());
   HA_X1 i_8_0_251 (.A(\out_as[3] [6]), .B(n_8_0_528), .CO(n_8_0_251), .S());
   HA_X1 i_8_0_252 (.A(\out_as[4] [6]), .B(n_8_0_1072), .CO(n_8_0_252), .S());
   HA_X1 i_8_0_253 (.A(\out_as[4] [6]), .B(n_8_0_1070), .CO(n_8_0_253), .S());
   HA_X1 i_8_0_254 (.A(\out_as[4] [6]), .B(n_8_0_1068), .CO(n_8_0_254), .S());
   HA_X1 i_8_0_255 (.A(\out_as[4] [6]), .B(n_8_0_1067), .CO(n_8_0_255), .S());
   HA_X1 i_8_0_256 (.A(\out_as[4] [6]), .B(n_8_0_1234), .CO(n_8_0_256), .S());
   HA_X1 i_8_0_257 (.A(\out_as[4] [6]), .B(n_8_0_1066), .CO(n_8_0_257), .S());
   HA_X1 i_8_0_258 (.A(\out_as[4] [6]), .B(n_8_0_1065), .CO(n_8_0_258), .S());
   HA_X1 i_8_0_259 (.A(\out_as[4] [6]), .B(n_8_0_1074), .CO(n_8_0_259), .S());
   HA_X1 i_8_0_260 (.A(\out_as[4] [6]), .B(n_8_0_1064), .CO(n_8_0_260), .S());
   HA_X1 i_8_0_261 (.A(\out_as[4] [6]), .B(n_8_0_1063), .CO(n_8_0_261), .S());
   HA_X1 i_8_0_262 (.A(\out_as[4] [6]), .B(n_8_0_1062), .CO(n_8_0_262), .S());
   HA_X1 i_8_0_263 (.A(\out_as[4] [6]), .B(n_8_0_1061), .CO(n_8_0_263), .S());
   HA_X1 i_8_0_264 (.A(\out_as[4] [6]), .B(n_8_0_1060), .CO(n_8_0_264), .S());
   HA_X1 i_8_0_265 (.A(\out_as[4] [6]), .B(n_8_0_1059), .CO(n_8_0_265), .S());
   HA_X1 i_8_0_266 (.A(\out_as[4] [6]), .B(n_8_0_1058), .CO(n_8_0_266), .S());
   HA_X1 i_8_0_267 (.A(\out_as[4] [6]), .B(n_8_0_1357), .CO(n_8_0_267), .S());
   HA_X1 i_8_0_268 (.A(\out_as[4] [6]), .B(n_8_0_1362), .CO(n_8_0_268), .S());
   HA_X1 i_8_0_269 (.A(\out_as[4] [6]), .B(n_8_0_1057), .CO(n_8_0_269), .S());
   HA_X1 i_8_0_270 (.A(\out_as[4] [6]), .B(n_8_0_1056), .CO(n_8_0_270), .S());
   HA_X1 i_8_0_271 (.A(\out_as[4] [6]), .B(n_8_0_1055), .CO(n_8_0_271), .S());
   HA_X1 i_8_0_272 (.A(\out_as[4] [6]), .B(n_8_0_1054), .CO(n_8_0_272), .S());
   HA_X1 i_8_0_273 (.A(\out_as[4] [6]), .B(n_8_0_1053), .CO(n_8_0_273), .S());
   HA_X1 i_8_0_274 (.A(\out_as[4] [6]), .B(n_8_0_1052), .CO(n_8_0_274), .S());
   HA_X1 i_8_0_275 (.A(\out_as[4] [6]), .B(n_8_0_1386), .CO(n_8_0_275), .S());
   HA_X1 i_8_0_276 (.A(\out_as[4] [6]), .B(n_8_0_1051), .CO(n_8_0_276), .S());
   HA_X1 i_8_0_277 (.A(\out_as[4] [6]), .B(n_8_0_1050), .CO(n_8_0_277), .S());
   HA_X1 i_8_0_278 (.A(\out_as[4] [6]), .B(n_8_0_1395), .CO(n_8_0_278), .S());
   HA_X1 i_8_0_279 (.A(\out_as[4] [6]), .B(n_8_0_1401), .CO(n_8_0_279), .S());
   HA_X1 i_8_0_280 (.A(\out_as[4] [6]), .B(n_8_0_1405), .CO(n_8_0_280), .S());
   HA_X1 i_8_0_281 (.A(\out_as[4] [6]), .B(n_8_0_1049), .CO(n_8_0_281), .S());
   HA_X1 i_8_0_282 (.A(\out_as[4] [6]), .B(n_8_0_1414), .CO(n_8_0_282), .S());
   HA_X1 i_8_0_283 (.A(\out_as[4] [6]), .B(\out_as[4] [5]), .CO(n_8_0_283), 
      .S());
   HA_X1 i_8_0_284 (.A(\out_as[4] [6]), .B(n_8_0_955), .CO(n_8_0_284), .S());
   HA_X1 i_8_0_285 (.A(\out_as[4] [6]), .B(n_8_0_947), .CO(n_8_0_285), .S());
   HA_X1 i_8_0_286 (.A(\out_as[4] [6]), .B(n_8_0_939), .CO(n_8_0_286), .S());
   HA_X1 i_8_0_287 (.A(\out_as[4] [6]), .B(n_8_0_931), .CO(n_8_0_287), .S());
   HA_X1 i_8_0_288 (.A(\out_as[4] [6]), .B(n_8_0_923), .CO(n_8_0_288), .S());
   HA_X1 i_8_0_289 (.A(\out_as[4] [6]), .B(n_8_0_915), .CO(n_8_0_289), .S());
   HA_X1 i_8_0_290 (.A(\out_as[4] [6]), .B(n_8_0_907), .CO(n_8_0_290), .S());
   HA_X1 i_8_0_291 (.A(\out_as[4] [6]), .B(n_8_0_899), .CO(n_8_0_291), .S());
   HA_X1 i_8_0_292 (.A(\out_as[4] [6]), .B(n_8_0_891), .CO(n_8_0_292), .S());
   HA_X1 i_8_0_293 (.A(\out_as[4] [6]), .B(n_8_0_883), .CO(n_8_0_293), .S());
   HA_X1 i_8_0_294 (.A(\out_as[4] [6]), .B(n_8_0_875), .CO(n_8_0_294), .S());
   HA_X1 i_8_0_295 (.A(\out_as[4] [6]), .B(n_8_0_867), .CO(n_8_0_295), .S());
   HA_X1 i_8_0_296 (.A(\out_as[4] [6]), .B(n_8_0_859), .CO(n_8_0_296), .S());
   HA_X1 i_8_0_297 (.A(\out_as[4] [6]), .B(n_8_0_851), .CO(n_8_0_297), .S());
   HA_X1 i_8_0_298 (.A(\out_as[4] [6]), .B(n_8_0_843), .CO(n_8_0_298), .S());
   HA_X1 i_8_0_299 (.A(\out_as[4] [6]), .B(n_8_0_835), .CO(n_8_0_299), .S());
   HA_X1 i_8_0_300 (.A(\out_as[4] [6]), .B(n_8_0_823), .CO(n_8_0_300), .S());
   HA_X1 i_8_0_301 (.A(\out_as[4] [6]), .B(n_8_0_807), .CO(n_8_0_301), .S());
   HA_X1 i_8_0_302 (.A(\out_as[4] [6]), .B(n_8_0_791), .CO(n_8_0_302), .S());
   HA_X1 i_8_0_303 (.A(\out_as[4] [6]), .B(n_8_0_775), .CO(n_8_0_303), .S());
   HA_X1 i_8_0_304 (.A(\out_as[4] [6]), .B(n_8_0_759), .CO(n_8_0_304), .S());
   HA_X1 i_8_0_305 (.A(\out_as[4] [6]), .B(n_8_0_743), .CO(n_8_0_305), .S());
   HA_X1 i_8_0_306 (.A(\out_as[4] [6]), .B(n_8_0_727), .CO(n_8_0_306), .S());
   HA_X1 i_8_0_307 (.A(\out_as[4] [6]), .B(n_8_0_711), .CO(n_8_0_307), .S());
   HA_X1 i_8_0_308 (.A(\out_as[4] [6]), .B(n_8_0_691), .CO(n_8_0_308), .S());
   HA_X1 i_8_0_309 (.A(\out_as[4] [6]), .B(n_8_0_667), .CO(n_8_0_309), .S());
   HA_X1 i_8_0_310 (.A(\out_as[4] [6]), .B(n_8_0_643), .CO(n_8_0_310), .S());
   HA_X1 i_8_0_311 (.A(\out_as[4] [6]), .B(n_8_0_619), .CO(n_8_0_311), .S());
   HA_X1 i_8_0_312 (.A(\out_as[4] [6]), .B(n_8_0_591), .CO(n_8_0_312), .S());
   HA_X1 i_8_0_313 (.A(\out_as[4] [6]), .B(n_8_0_559), .CO(n_8_0_313), .S());
   HA_X1 i_8_0_314 (.A(\out_as[4] [6]), .B(n_8_0_523), .CO(n_8_0_314), .S());
   HA_X1 i_8_0_315 (.A(\out_as[5] [6]), .B(n_8_0_1045), .CO(n_8_0_315), .S());
   HA_X1 i_8_0_316 (.A(\out_as[5] [6]), .B(n_8_0_1198), .CO(n_8_0_316), .S());
   HA_X1 i_8_0_317 (.A(\out_as[5] [6]), .B(n_8_0_1043), .CO(n_8_0_317), .S());
   HA_X1 i_8_0_318 (.A(\out_as[5] [6]), .B(n_8_0_1215), .CO(n_8_0_318), .S());
   HA_X1 i_8_0_319 (.A(\out_as[5] [6]), .B(n_8_0_1042), .CO(n_8_0_319), .S());
   HA_X1 i_8_0_320 (.A(\out_as[5] [6]), .B(n_8_0_1041), .CO(n_8_0_320), .S());
   HA_X1 i_8_0_321 (.A(\out_as[5] [6]), .B(n_8_0_1274), .CO(n_8_0_321), .S());
   HA_X1 i_8_0_322 (.A(\out_as[5] [6]), .B(n_8_0_1216), .CO(n_8_0_322), .S());
   HA_X1 i_8_0_323 (.A(\out_as[5] [6]), .B(n_8_0_1040), .CO(n_8_0_323), .S());
   HA_X1 i_8_0_324 (.A(\out_as[5] [6]), .B(n_8_0_1039), .CO(n_8_0_324), .S());
   HA_X1 i_8_0_325 (.A(\out_as[5] [6]), .B(n_8_0_1037), .CO(n_8_0_325), .S());
   HA_X1 i_8_0_326 (.A(\out_as[5] [6]), .B(n_8_0_1035), .CO(n_8_0_326), .S());
   HA_X1 i_8_0_327 (.A(\out_as[5] [6]), .B(n_8_0_1033), .CO(n_8_0_327), .S());
   HA_X1 i_8_0_328 (.A(\out_as[5] [6]), .B(n_8_0_1031), .CO(n_8_0_328), .S());
   HA_X1 i_8_0_329 (.A(\out_as[5] [6]), .B(n_8_0_1030), .CO(n_8_0_329), .S());
   HA_X1 i_8_0_330 (.A(\out_as[5] [6]), .B(n_8_0_1354), .CO(n_8_0_330), .S());
   HA_X1 i_8_0_331 (.A(\out_as[5] [6]), .B(n_8_0_1029), .CO(n_8_0_331), .S());
   HA_X1 i_8_0_332 (.A(\out_as[5] [6]), .B(n_8_0_1028), .CO(n_8_0_332), .S());
   HA_X1 i_8_0_333 (.A(\out_as[5] [6]), .B(n_8_0_1027), .CO(n_8_0_333), .S());
   HA_X1 i_8_0_334 (.A(\out_as[5] [6]), .B(n_8_0_1026), .CO(n_8_0_334), .S());
   HA_X1 i_8_0_335 (.A(\out_as[5] [6]), .B(n_8_0_1025), .CO(n_8_0_335), .S());
   HA_X1 i_8_0_336 (.A(\out_as[5] [6]), .B(n_8_0_1024), .CO(n_8_0_336), .S());
   HA_X1 i_8_0_337 (.A(\out_as[5] [6]), .B(n_8_0_1023), .CO(n_8_0_337), .S());
   HA_X1 i_8_0_338 (.A(\out_as[5] [6]), .B(n_8_0_1022), .CO(n_8_0_338), .S());
   HA_X1 i_8_0_339 (.A(\out_as[5] [6]), .B(n_8_0_1021), .CO(n_8_0_339), .S());
   HA_X1 i_8_0_340 (.A(\out_as[5] [6]), .B(n_8_0_1392), .CO(n_8_0_340), .S());
   HA_X1 i_8_0_341 (.A(\out_as[5] [6]), .B(n_8_0_1020), .CO(n_8_0_341), .S());
   HA_X1 i_8_0_342 (.A(\out_as[5] [6]), .B(n_8_0_1019), .CO(n_8_0_342), .S());
   HA_X1 i_8_0_343 (.A(\out_as[5] [6]), .B(n_8_0_1018), .CO(n_8_0_343), .S());
   HA_X1 i_8_0_344 (.A(\out_as[5] [6]), .B(n_8_0_1017), .CO(n_8_0_344), .S());
   HA_X1 i_8_0_345 (.A(\out_as[5] [6]), .B(n_8_0_1016), .CO(n_8_0_345), .S());
   HA_X1 i_8_0_346 (.A(\out_as[5] [6]), .B(\out_as[5] [5]), .CO(n_8_0_346), 
      .S());
   HA_X1 i_8_0_347 (.A(\out_as[5] [6]), .B(n_8_0_954), .CO(n_8_0_347), .S());
   HA_X1 i_8_0_348 (.A(\out_as[5] [6]), .B(n_8_0_946), .CO(n_8_0_348), .S());
   HA_X1 i_8_0_349 (.A(\out_as[5] [6]), .B(n_8_0_938), .CO(n_8_0_349), .S());
   HA_X1 i_8_0_350 (.A(\out_as[5] [6]), .B(n_8_0_930), .CO(n_8_0_350), .S());
   HA_X1 i_8_0_351 (.A(\out_as[5] [6]), .B(n_8_0_922), .CO(n_8_0_351), .S());
   HA_X1 i_8_0_352 (.A(\out_as[5] [6]), .B(n_8_0_914), .CO(n_8_0_352), .S());
   HA_X1 i_8_0_353 (.A(\out_as[5] [6]), .B(n_8_0_906), .CO(n_8_0_353), .S());
   HA_X1 i_8_0_354 (.A(\out_as[5] [6]), .B(n_8_0_898), .CO(n_8_0_354), .S());
   HA_X1 i_8_0_355 (.A(\out_as[5] [6]), .B(n_8_0_890), .CO(n_8_0_355), .S());
   HA_X1 i_8_0_356 (.A(\out_as[5] [6]), .B(n_8_0_882), .CO(n_8_0_356), .S());
   HA_X1 i_8_0_357 (.A(\out_as[5] [6]), .B(n_8_0_874), .CO(n_8_0_357), .S());
   HA_X1 i_8_0_358 (.A(\out_as[5] [6]), .B(n_8_0_866), .CO(n_8_0_358), .S());
   HA_X1 i_8_0_359 (.A(\out_as[5] [6]), .B(n_8_0_858), .CO(n_8_0_359), .S());
   HA_X1 i_8_0_360 (.A(\out_as[5] [6]), .B(n_8_0_850), .CO(n_8_0_360), .S());
   HA_X1 i_8_0_361 (.A(\out_as[5] [6]), .B(n_8_0_842), .CO(n_8_0_361), .S());
   HA_X1 i_8_0_362 (.A(\out_as[5] [6]), .B(n_8_0_834), .CO(n_8_0_362), .S());
   HA_X1 i_8_0_363 (.A(\out_as[5] [6]), .B(n_8_0_821), .CO(n_8_0_363), .S());
   HA_X1 i_8_0_364 (.A(\out_as[5] [6]), .B(n_8_0_805), .CO(n_8_0_364), .S());
   HA_X1 i_8_0_365 (.A(\out_as[5] [6]), .B(n_8_0_789), .CO(n_8_0_365), .S());
   HA_X1 i_8_0_366 (.A(\out_as[5] [6]), .B(n_8_0_773), .CO(n_8_0_366), .S());
   HA_X1 i_8_0_367 (.A(\out_as[5] [6]), .B(n_8_0_757), .CO(n_8_0_367), .S());
   HA_X1 i_8_0_368 (.A(\out_as[5] [6]), .B(n_8_0_741), .CO(n_8_0_368), .S());
   HA_X1 i_8_0_369 (.A(\out_as[5] [6]), .B(n_8_0_725), .CO(n_8_0_369), .S());
   HA_X1 i_8_0_370 (.A(\out_as[5] [6]), .B(n_8_0_709), .CO(n_8_0_370), .S());
   HA_X1 i_8_0_371 (.A(\out_as[5] [6]), .B(n_8_0_688), .CO(n_8_0_371), .S());
   HA_X1 i_8_0_372 (.A(\out_as[5] [6]), .B(n_8_0_664), .CO(n_8_0_372), .S());
   HA_X1 i_8_0_373 (.A(\out_as[5] [6]), .B(n_8_0_640), .CO(n_8_0_373), .S());
   HA_X1 i_8_0_374 (.A(\out_as[5] [6]), .B(n_8_0_616), .CO(n_8_0_374), .S());
   HA_X1 i_8_0_375 (.A(\out_as[5] [6]), .B(n_8_0_587), .CO(n_8_0_375), .S());
   HA_X1 i_8_0_376 (.A(\out_as[5] [6]), .B(n_8_0_555), .CO(n_8_0_376), .S());
   HA_X1 i_8_0_377 (.A(\out_as[5] [6]), .B(n_8_0_518), .CO(n_8_0_377), .S());
   HA_X1 i_8_0_378 (.A(\out_as[6] [6]), .B(n_8_0_1015), .CO(n_8_0_378), .S());
   HA_X1 i_8_0_379 (.A(\out_as[6] [6]), .B(n_8_0_1014), .CO(n_8_0_379), .S());
   HA_X1 i_8_0_380 (.A(\out_as[6] [6]), .B(n_8_0_1012), .CO(n_8_0_380), .S());
   HA_X1 i_8_0_381 (.A(\out_as[6] [6]), .B(n_8_0_1219), .CO(n_8_0_381), .S());
   HA_X1 i_8_0_382 (.A(\out_as[6] [6]), .B(n_8_0_1245), .CO(n_8_0_382), .S());
   HA_X1 i_8_0_383 (.A(\out_as[6] [6]), .B(n_8_0_1259), .CO(n_8_0_383), .S());
   HA_X1 i_8_0_384 (.A(\out_as[6] [6]), .B(n_8_0_1270), .CO(n_8_0_384), .S());
   HA_X1 i_8_0_385 (.A(\out_as[6] [6]), .B(n_8_0_1271), .CO(n_8_0_385), .S());
   HA_X1 i_8_0_386 (.A(\out_as[6] [6]), .B(n_8_0_1011), .CO(n_8_0_386), .S());
   HA_X1 i_8_0_387 (.A(\out_as[6] [6]), .B(n_8_0_1009), .CO(n_8_0_387), .S());
   HA_X1 i_8_0_388 (.A(\out_as[6] [6]), .B(n_8_0_1008), .CO(n_8_0_388), .S());
   HA_X1 i_8_0_389 (.A(\out_as[6] [6]), .B(n_8_0_1327), .CO(n_8_0_389), .S());
   HA_X1 i_8_0_390 (.A(\out_as[6] [6]), .B(n_8_0_1007), .CO(n_8_0_390), .S());
   HA_X1 i_8_0_391 (.A(\out_as[6] [6]), .B(n_8_0_1006), .CO(n_8_0_391), .S());
   HA_X1 i_8_0_392 (.A(\out_as[6] [6]), .B(n_8_0_1005), .CO(n_8_0_392), .S());
   HA_X1 i_8_0_393 (.A(\out_as[6] [6]), .B(n_8_0_1358), .CO(n_8_0_393), .S());
   HA_X1 i_8_0_394 (.A(\out_as[6] [6]), .B(n_8_0_1365), .CO(n_8_0_394), .S());
   HA_X1 i_8_0_395 (.A(\out_as[6] [6]), .B(n_8_0_1371), .CO(n_8_0_395), .S());
   HA_X1 i_8_0_396 (.A(\out_as[6] [6]), .B(n_8_0_1372), .CO(n_8_0_396), .S());
   HA_X1 i_8_0_397 (.A(\out_as[6] [6]), .B(n_8_0_1375), .CO(n_8_0_397), .S());
   HA_X1 i_8_0_398 (.A(\out_as[6] [6]), .B(n_8_0_1379), .CO(n_8_0_398), .S());
   HA_X1 i_8_0_399 (.A(\out_as[6] [6]), .B(n_8_0_1004), .CO(n_8_0_399), .S());
   HA_X1 i_8_0_400 (.A(\out_as[6] [6]), .B(n_8_0_1381), .CO(n_8_0_400), .S());
   HA_X1 i_8_0_401 (.A(\out_as[6] [6]), .B(n_8_0_1003), .CO(n_8_0_401), .S());
   HA_X1 i_8_0_402 (.A(\out_as[6] [6]), .B(n_8_0_1391), .CO(n_8_0_402), .S());
   HA_X1 i_8_0_403 (.A(\out_as[6] [6]), .B(n_8_0_1393), .CO(n_8_0_403), .S());
   HA_X1 i_8_0_404 (.A(\out_as[6] [6]), .B(n_8_0_1397), .CO(n_8_0_404), .S());
   HA_X1 i_8_0_405 (.A(\out_as[6] [6]), .B(n_8_0_1002), .CO(n_8_0_405), .S());
   HA_X1 i_8_0_406 (.A(\out_as[6] [6]), .B(n_8_0_1403), .CO(n_8_0_406), .S());
   HA_X1 i_8_0_407 (.A(\out_as[6] [6]), .B(n_8_0_1408), .CO(n_8_0_407), .S());
   HA_X1 i_8_0_408 (.A(\out_as[6] [6]), .B(n_8_0_1415), .CO(n_8_0_408), .S());
   HA_X1 i_8_0_409 (.A(\out_as[6] [6]), .B(\out_as[6] [5]), .CO(n_8_0_409), 
      .S());
   HA_X1 i_8_0_410 (.A(\out_as[6] [6]), .B(n_8_0_953), .CO(n_8_0_410), .S());
   HA_X1 i_8_0_411 (.A(\out_as[6] [6]), .B(n_8_0_945), .CO(n_8_0_411), .S());
   HA_X1 i_8_0_412 (.A(\out_as[6] [6]), .B(n_8_0_937), .CO(n_8_0_412), .S());
   HA_X1 i_8_0_413 (.A(\out_as[6] [6]), .B(n_8_0_929), .CO(n_8_0_413), .S());
   HA_X1 i_8_0_414 (.A(\out_as[6] [6]), .B(n_8_0_921), .CO(n_8_0_414), .S());
   HA_X1 i_8_0_415 (.A(\out_as[6] [6]), .B(n_8_0_913), .CO(n_8_0_415), .S());
   HA_X1 i_8_0_416 (.A(\out_as[6] [6]), .B(n_8_0_905), .CO(n_8_0_416), .S());
   HA_X1 i_8_0_417 (.A(\out_as[6] [6]), .B(n_8_0_897), .CO(n_8_0_417), .S());
   HA_X1 i_8_0_418 (.A(\out_as[6] [6]), .B(n_8_0_889), .CO(n_8_0_418), .S());
   HA_X1 i_8_0_419 (.A(\out_as[6] [6]), .B(n_8_0_881), .CO(n_8_0_419), .S());
   HA_X1 i_8_0_420 (.A(\out_as[6] [6]), .B(n_8_0_873), .CO(n_8_0_420), .S());
   HA_X1 i_8_0_421 (.A(\out_as[6] [6]), .B(n_8_0_865), .CO(n_8_0_421), .S());
   HA_X1 i_8_0_422 (.A(\out_as[6] [6]), .B(n_8_0_857), .CO(n_8_0_422), .S());
   HA_X1 i_8_0_423 (.A(\out_as[6] [6]), .B(n_8_0_849), .CO(n_8_0_423), .S());
   HA_X1 i_8_0_424 (.A(\out_as[6] [6]), .B(n_8_0_841), .CO(n_8_0_424), .S());
   HA_X1 i_8_0_425 (.A(\out_as[6] [6]), .B(n_8_0_833), .CO(n_8_0_425), .S());
   HA_X1 i_8_0_426 (.A(\out_as[6] [6]), .B(n_8_0_819), .CO(n_8_0_426), .S());
   HA_X1 i_8_0_427 (.A(\out_as[6] [6]), .B(n_8_0_803), .CO(n_8_0_427), .S());
   HA_X1 i_8_0_428 (.A(\out_as[6] [6]), .B(n_8_0_787), .CO(n_8_0_428), .S());
   HA_X1 i_8_0_429 (.A(\out_as[6] [6]), .B(n_8_0_771), .CO(n_8_0_429), .S());
   HA_X1 i_8_0_430 (.A(\out_as[6] [6]), .B(n_8_0_755), .CO(n_8_0_430), .S());
   HA_X1 i_8_0_431 (.A(\out_as[6] [6]), .B(n_8_0_739), .CO(n_8_0_431), .S());
   HA_X1 i_8_0_432 (.A(\out_as[6] [6]), .B(n_8_0_723), .CO(n_8_0_432), .S());
   HA_X1 i_8_0_433 (.A(\out_as[6] [6]), .B(n_8_0_707), .CO(n_8_0_433), .S());
   HA_X1 i_8_0_434 (.A(\out_as[6] [6]), .B(n_8_0_685), .CO(n_8_0_434), .S());
   HA_X1 i_8_0_435 (.A(\out_as[6] [6]), .B(n_8_0_661), .CO(n_8_0_435), .S());
   HA_X1 i_8_0_436 (.A(\out_as[6] [6]), .B(n_8_0_637), .CO(n_8_0_436), .S());
   HA_X1 i_8_0_437 (.A(\out_as[6] [6]), .B(n_8_0_613), .CO(n_8_0_437), .S());
   HA_X1 i_8_0_438 (.A(\out_as[6] [6]), .B(n_8_0_583), .CO(n_8_0_438), .S());
   HA_X1 i_8_0_439 (.A(\out_as[6] [6]), .B(n_8_0_551), .CO(n_8_0_439), .S());
   HA_X1 i_8_0_440 (.A(\out_as[6] [6]), .B(n_8_0_513), .CO(n_8_0_440), .S());
   HA_X1 i_8_0_441 (.A(\out_as[7] [6]), .B(n_8_0_998), .CO(n_8_0_441), .S());
   HA_X1 i_8_0_442 (.A(\out_as[7] [6]), .B(n_8_0_996), .CO(n_8_0_442), .S());
   HA_X1 i_8_0_443 (.A(\out_as[7] [6]), .B(n_8_0_994), .CO(n_8_0_443), .S());
   HA_X1 i_8_0_444 (.A(\out_as[7] [6]), .B(n_8_0_993), .CO(n_8_0_444), .S());
   HA_X1 i_8_0_445 (.A(\out_as[7] [6]), .B(n_8_0_992), .CO(n_8_0_445), .S());
   HA_X1 i_8_0_446 (.A(\out_as[7] [6]), .B(n_8_0_990), .CO(n_8_0_446), .S());
   HA_X1 i_8_0_447 (.A(\out_as[7] [6]), .B(n_8_0_989), .CO(n_8_0_447), .S());
   HA_X1 i_8_0_448 (.A(\out_as[7] [6]), .B(n_8_0_999), .CO(n_8_0_448), .S());
   HA_X1 i_8_0_449 (.A(\out_as[7] [6]), .B(n_8_0_988), .CO(n_8_0_449), .S());
   HA_X1 i_8_0_450 (.A(\out_as[7] [6]), .B(n_8_0_987), .CO(n_8_0_450), .S());
   HA_X1 i_8_0_451 (.A(\out_as[7] [6]), .B(n_8_0_986), .CO(n_8_0_451), .S());
   HA_X1 i_8_0_452 (.A(\out_as[7] [6]), .B(n_8_0_985), .CO(n_8_0_452), .S());
   HA_X1 i_8_0_453 (.A(\out_as[7] [6]), .B(n_8_0_984), .CO(n_8_0_453), .S());
   HA_X1 i_8_0_454 (.A(\out_as[7] [6]), .B(n_8_0_983), .CO(n_8_0_454), .S());
   HA_X1 i_8_0_455 (.A(\out_as[7] [6]), .B(n_8_0_982), .CO(n_8_0_455), .S());
   HA_X1 i_8_0_456 (.A(\out_as[7] [6]), .B(n_8_0_1360), .CO(n_8_0_456), .S());
   HA_X1 i_8_0_457 (.A(\out_as[7] [6]), .B(n_8_0_1366), .CO(n_8_0_457), .S());
   HA_X1 i_8_0_458 (.A(\out_as[7] [6]), .B(n_8_0_1367), .CO(n_8_0_458), .S());
   HA_X1 i_8_0_459 (.A(\out_as[7] [6]), .B(n_8_0_981), .CO(n_8_0_459), .S());
   HA_X1 i_8_0_460 (.A(\out_as[7] [6]), .B(n_8_0_980), .CO(n_8_0_460), .S());
   HA_X1 i_8_0_461 (.A(\out_as[7] [6]), .B(n_8_0_979), .CO(n_8_0_461), .S());
   HA_X1 i_8_0_462 (.A(\out_as[7] [6]), .B(n_8_0_978), .CO(n_8_0_462), .S());
   HA_X1 i_8_0_463 (.A(\out_as[7] [6]), .B(n_8_0_1384), .CO(n_8_0_463), .S());
   HA_X1 i_8_0_464 (.A(\out_as[7] [6]), .B(n_8_0_977), .CO(n_8_0_464), .S());
   HA_X1 i_8_0_465 (.A(\out_as[7] [6]), .B(n_8_0_1389), .CO(n_8_0_465), .S());
   HA_X1 i_8_0_466 (.A(\out_as[7] [6]), .B(n_8_0_976), .CO(n_8_0_466), .S());
   HA_X1 i_8_0_467 (.A(\out_as[7] [6]), .B(n_8_0_1394), .CO(n_8_0_467), .S());
   HA_X1 i_8_0_468 (.A(\out_as[7] [6]), .B(n_8_0_1399), .CO(n_8_0_468), .S());
   HA_X1 i_8_0_469 (.A(\out_as[7] [6]), .B(n_8_0_1404), .CO(n_8_0_469), .S());
   HA_X1 i_8_0_470 (.A(\out_as[7] [6]), .B(n_8_0_1409), .CO(n_8_0_470), .S());
   HA_X1 i_8_0_471 (.A(\out_as[7] [6]), .B(n_8_0_1411), .CO(n_8_0_471), .S());
   HA_X1 i_8_0_472 (.A(\out_as[7] [6]), .B(\out_as[7] [5]), .CO(n_8_0_472), 
      .S());
   HA_X1 i_8_0_473 (.A(\out_as[7] [6]), .B(n_8_0_952), .CO(n_8_0_473), .S());
   HA_X1 i_8_0_474 (.A(\out_as[7] [6]), .B(n_8_0_944), .CO(n_8_0_474), .S());
   HA_X1 i_8_0_475 (.A(\out_as[7] [6]), .B(n_8_0_936), .CO(n_8_0_475), .S());
   HA_X1 i_8_0_476 (.A(\out_as[7] [6]), .B(n_8_0_928), .CO(n_8_0_476), .S());
   HA_X1 i_8_0_477 (.A(\out_as[7] [6]), .B(n_8_0_920), .CO(n_8_0_477), .S());
   HA_X1 i_8_0_478 (.A(\out_as[7] [6]), .B(n_8_0_912), .CO(n_8_0_478), .S());
   HA_X1 i_8_0_479 (.A(\out_as[7] [6]), .B(n_8_0_904), .CO(n_8_0_479), .S());
   HA_X1 i_8_0_480 (.A(\out_as[7] [6]), .B(n_8_0_896), .CO(n_8_0_480), .S());
   HA_X1 i_8_0_481 (.A(\out_as[7] [6]), .B(n_8_0_888), .CO(n_8_0_481), .S());
   HA_X1 i_8_0_482 (.A(\out_as[7] [6]), .B(n_8_0_880), .CO(n_8_0_482), .S());
   HA_X1 i_8_0_483 (.A(\out_as[7] [6]), .B(n_8_0_872), .CO(n_8_0_483), .S());
   HA_X1 i_8_0_484 (.A(\out_as[7] [6]), .B(n_8_0_864), .CO(n_8_0_484), .S());
   HA_X1 i_8_0_485 (.A(\out_as[7] [6]), .B(n_8_0_856), .CO(n_8_0_485), .S());
   HA_X1 i_8_0_486 (.A(\out_as[7] [6]), .B(n_8_0_848), .CO(n_8_0_486), .S());
   HA_X1 i_8_0_487 (.A(\out_as[7] [6]), .B(n_8_0_840), .CO(n_8_0_487), .S());
   HA_X1 i_8_0_488 (.A(\out_as[7] [6]), .B(n_8_0_832), .CO(n_8_0_488), .S());
   HA_X1 i_8_0_489 (.A(\out_as[7] [6]), .B(n_8_0_817), .CO(n_8_0_489), .S());
   HA_X1 i_8_0_490 (.A(\out_as[7] [6]), .B(n_8_0_801), .CO(n_8_0_490), .S());
   HA_X1 i_8_0_491 (.A(\out_as[7] [6]), .B(n_8_0_785), .CO(n_8_0_491), .S());
   HA_X1 i_8_0_492 (.A(\out_as[7] [6]), .B(n_8_0_769), .CO(n_8_0_492), .S());
   HA_X1 i_8_0_493 (.A(\out_as[7] [6]), .B(n_8_0_753), .CO(n_8_0_493), .S());
   HA_X1 i_8_0_494 (.A(\out_as[7] [6]), .B(n_8_0_737), .CO(n_8_0_494), .S());
   HA_X1 i_8_0_495 (.A(\out_as[7] [6]), .B(n_8_0_721), .CO(n_8_0_495), .S());
   HA_X1 i_8_0_496 (.A(\out_as[7] [6]), .B(n_8_0_705), .CO(n_8_0_496), .S());
   HA_X1 i_8_0_497 (.A(\out_as[7] [6]), .B(n_8_0_682), .CO(n_8_0_497), .S());
   HA_X1 i_8_0_498 (.A(\out_as[7] [6]), .B(n_8_0_658), .CO(n_8_0_498), .S());
   HA_X1 i_8_0_499 (.A(\out_as[7] [6]), .B(n_8_0_634), .CO(n_8_0_499), .S());
   HA_X1 i_8_0_500 (.A(\out_as[7] [6]), .B(n_8_0_610), .CO(n_8_0_500), .S());
   HA_X1 i_8_0_501 (.A(\out_as[7] [6]), .B(n_8_0_579), .CO(n_8_0_501), .S());
   HA_X1 i_8_0_502 (.A(\out_as[7] [6]), .B(n_8_0_547), .CO(n_8_0_502), .S());
   HA_X1 i_8_0_503 (.A(\out_as[7] [6]), .B(n_8_0_508), .CO(n_8_0_503), .S());
   HA_X1 i_8_0_504 (.A(\out_as[7] [1]), .B(\out_as[7] [0]), .CO(n_8_0_504), 
      .S());
   HA_X1 i_8_0_505 (.A(\out_as[7] [2]), .B(n_8_0_504), .CO(n_8_0_505), .S());
   HA_X1 i_8_0_506 (.A(\out_as[7] [3]), .B(n_8_0_505), .CO(n_8_0_506), .S());
   HA_X1 i_8_0_507 (.A(\out_as[7] [4]), .B(n_8_0_506), .CO(n_8_0_507), .S());
   HA_X1 i_8_0_508 (.A(\out_as[7] [5]), .B(n_8_0_507), .CO(n_8_0_508), .S());
   HA_X1 i_8_0_509 (.A(\out_as[6] [1]), .B(\out_as[6] [0]), .CO(n_8_0_509), 
      .S());
   HA_X1 i_8_0_510 (.A(\out_as[6] [2]), .B(n_8_0_509), .CO(n_8_0_510), .S());
   HA_X1 i_8_0_511 (.A(\out_as[6] [3]), .B(n_8_0_510), .CO(n_8_0_511), .S());
   HA_X1 i_8_0_512 (.A(\out_as[6] [4]), .B(n_8_0_511), .CO(n_8_0_512), .S());
   HA_X1 i_8_0_513 (.A(\out_as[6] [5]), .B(n_8_0_512), .CO(n_8_0_513), .S());
   HA_X1 i_8_0_514 (.A(\out_as[5] [1]), .B(\out_as[5] [0]), .CO(n_8_0_514), 
      .S());
   HA_X1 i_8_0_515 (.A(\out_as[5] [2]), .B(n_8_0_514), .CO(n_8_0_515), .S());
   HA_X1 i_8_0_516 (.A(\out_as[5] [3]), .B(n_8_0_515), .CO(n_8_0_516), .S());
   HA_X1 i_8_0_517 (.A(\out_as[5] [4]), .B(n_8_0_516), .CO(n_8_0_517), .S());
   HA_X1 i_8_0_518 (.A(\out_as[5] [5]), .B(n_8_0_517), .CO(n_8_0_518), .S());
   HA_X1 i_8_0_519 (.A(\out_as[4] [1]), .B(\out_as[4] [0]), .CO(n_8_0_519), 
      .S());
   HA_X1 i_8_0_520 (.A(\out_as[4] [2]), .B(n_8_0_519), .CO(n_8_0_520), .S());
   HA_X1 i_8_0_521 (.A(\out_as[4] [3]), .B(n_8_0_520), .CO(n_8_0_521), .S());
   HA_X1 i_8_0_522 (.A(\out_as[4] [4]), .B(n_8_0_521), .CO(n_8_0_522), .S());
   HA_X1 i_8_0_523 (.A(\out_as[4] [5]), .B(n_8_0_522), .CO(n_8_0_523), .S());
   HA_X1 i_8_0_524 (.A(\out_as[3] [1]), .B(\out_as[3] [0]), .CO(n_8_0_524), 
      .S());
   HA_X1 i_8_0_525 (.A(\out_as[3] [2]), .B(n_8_0_524), .CO(n_8_0_525), .S());
   HA_X1 i_8_0_526 (.A(\out_as[3] [3]), .B(n_8_0_525), .CO(n_8_0_526), .S());
   HA_X1 i_8_0_527 (.A(\out_as[3] [4]), .B(n_8_0_526), .CO(n_8_0_527), .S());
   HA_X1 i_8_0_528 (.A(\out_as[3] [5]), .B(n_8_0_527), .CO(n_8_0_528), .S());
   HA_X1 i_8_0_529 (.A(\out_as[2] [1]), .B(\out_as[2] [0]), .CO(n_8_0_529), 
      .S());
   HA_X1 i_8_0_530 (.A(\out_as[2] [2]), .B(n_8_0_529), .CO(n_8_0_530), .S());
   HA_X1 i_8_0_531 (.A(\out_as[2] [3]), .B(n_8_0_530), .CO(n_8_0_531), .S());
   HA_X1 i_8_0_532 (.A(\out_as[2] [4]), .B(n_8_0_531), .CO(n_8_0_532), .S());
   HA_X1 i_8_0_533 (.A(\out_as[2] [5]), .B(n_8_0_532), .CO(n_8_0_533), .S());
   HA_X1 i_8_0_534 (.A(\out_as[1] [1]), .B(\out_as[1] [0]), .CO(n_8_0_534), 
      .S());
   HA_X1 i_8_0_535 (.A(\out_as[1] [2]), .B(n_8_0_534), .CO(n_8_0_535), .S());
   HA_X1 i_8_0_536 (.A(\out_as[1] [3]), .B(n_8_0_535), .CO(n_8_0_536), .S());
   HA_X1 i_8_0_537 (.A(\out_as[1] [4]), .B(n_8_0_536), .CO(n_8_0_537), .S());
   HA_X1 i_8_0_538 (.A(\out_as[1] [5]), .B(n_8_0_537), .CO(n_8_0_538), .S());
   HA_X1 i_8_0_539 (.A(\out_as[0] [1]), .B(\out_as[0] [0]), .CO(n_8_0_539), 
      .S());
   HA_X1 i_8_0_540 (.A(\out_as[0] [2]), .B(n_8_0_539), .CO(n_8_0_540), .S());
   HA_X1 i_8_0_541 (.A(\out_as[0] [3]), .B(n_8_0_540), .CO(n_8_0_541), .S());
   HA_X1 i_8_0_542 (.A(\out_as[0] [4]), .B(n_8_0_541), .CO(n_8_0_542), .S());
   HA_X1 i_8_0_543 (.A(\out_as[0] [5]), .B(n_8_0_542), .CO(n_8_0_543), .S());
   HA_X1 i_8_0_544 (.A(\out_as[7] [2]), .B(\out_as[7] [1]), .CO(n_8_0_544), 
      .S());
   HA_X1 i_8_0_545 (.A(\out_as[7] [3]), .B(n_8_0_544), .CO(n_8_0_545), .S());
   HA_X1 i_8_0_546 (.A(\out_as[7] [4]), .B(n_8_0_545), .CO(n_8_0_546), .S());
   HA_X1 i_8_0_547 (.A(\out_as[7] [5]), .B(n_8_0_546), .CO(n_8_0_547), .S());
   HA_X1 i_8_0_548 (.A(\out_as[6] [2]), .B(\out_as[6] [1]), .CO(n_8_0_548), 
      .S());
   HA_X1 i_8_0_549 (.A(\out_as[6] [3]), .B(n_8_0_548), .CO(n_8_0_549), .S());
   HA_X1 i_8_0_550 (.A(\out_as[6] [4]), .B(n_8_0_549), .CO(n_8_0_550), .S());
   HA_X1 i_8_0_551 (.A(\out_as[6] [5]), .B(n_8_0_550), .CO(n_8_0_551), .S());
   HA_X1 i_8_0_552 (.A(\out_as[5] [2]), .B(\out_as[5] [1]), .CO(n_8_0_552), 
      .S());
   HA_X1 i_8_0_553 (.A(\out_as[5] [3]), .B(n_8_0_552), .CO(n_8_0_553), .S());
   HA_X1 i_8_0_554 (.A(\out_as[5] [4]), .B(n_8_0_553), .CO(n_8_0_554), .S());
   HA_X1 i_8_0_555 (.A(\out_as[5] [5]), .B(n_8_0_554), .CO(n_8_0_555), .S());
   HA_X1 i_8_0_556 (.A(\out_as[4] [2]), .B(\out_as[4] [1]), .CO(n_8_0_556), 
      .S());
   HA_X1 i_8_0_557 (.A(\out_as[4] [3]), .B(n_8_0_556), .CO(n_8_0_557), .S());
   HA_X1 i_8_0_558 (.A(\out_as[4] [4]), .B(n_8_0_557), .CO(n_8_0_558), .S());
   HA_X1 i_8_0_559 (.A(\out_as[4] [5]), .B(n_8_0_558), .CO(n_8_0_559), .S());
   HA_X1 i_8_0_560 (.A(\out_as[3] [2]), .B(\out_as[3] [1]), .CO(n_8_0_560), 
      .S());
   HA_X1 i_8_0_561 (.A(\out_as[3] [3]), .B(n_8_0_560), .CO(n_8_0_561), .S());
   HA_X1 i_8_0_562 (.A(\out_as[3] [4]), .B(n_8_0_561), .CO(n_8_0_562), .S());
   HA_X1 i_8_0_563 (.A(\out_as[3] [5]), .B(n_8_0_562), .CO(n_8_0_563), .S());
   HA_X1 i_8_0_564 (.A(\out_as[2] [2]), .B(\out_as[2] [1]), .CO(n_8_0_564), 
      .S());
   HA_X1 i_8_0_565 (.A(\out_as[2] [3]), .B(n_8_0_564), .CO(n_8_0_565), .S());
   HA_X1 i_8_0_566 (.A(\out_as[2] [4]), .B(n_8_0_565), .CO(n_8_0_566), .S());
   HA_X1 i_8_0_567 (.A(\out_as[2] [5]), .B(n_8_0_566), .CO(n_8_0_567), .S());
   HA_X1 i_8_0_568 (.A(\out_as[1] [2]), .B(\out_as[1] [1]), .CO(n_8_0_568), 
      .S());
   HA_X1 i_8_0_569 (.A(\out_as[1] [3]), .B(n_8_0_568), .CO(n_8_0_569), .S());
   HA_X1 i_8_0_570 (.A(\out_as[1] [4]), .B(n_8_0_569), .CO(n_8_0_570), .S());
   HA_X1 i_8_0_571 (.A(\out_as[1] [5]), .B(n_8_0_570), .CO(n_8_0_571), .S());
   HA_X1 i_8_0_572 (.A(\out_as[0] [2]), .B(\out_as[0] [1]), .CO(n_8_0_572), 
      .S());
   HA_X1 i_8_0_573 (.A(\out_as[0] [3]), .B(n_8_0_572), .CO(n_8_0_573), .S());
   HA_X1 i_8_0_574 (.A(\out_as[0] [4]), .B(n_8_0_573), .CO(n_8_0_574), .S());
   HA_X1 i_8_0_575 (.A(\out_as[0] [5]), .B(n_8_0_574), .CO(n_8_0_575), .S());
   HA_X1 i_8_0_576 (.A(\out_as[7] [2]), .B(n_8_0_1183), .CO(n_8_0_576), .S());
   HA_X1 i_8_0_577 (.A(\out_as[7] [3]), .B(n_8_0_576), .CO(n_8_0_577), .S());
   HA_X1 i_8_0_578 (.A(\out_as[7] [4]), .B(n_8_0_577), .CO(n_8_0_578), .S());
   HA_X1 i_8_0_579 (.A(\out_as[7] [5]), .B(n_8_0_578), .CO(n_8_0_579), .S());
   HA_X1 i_8_0_580 (.A(\out_as[6] [2]), .B(n_8_0_1181), .CO(n_8_0_580), .S());
   HA_X1 i_8_0_581 (.A(\out_as[6] [3]), .B(n_8_0_580), .CO(n_8_0_581), .S());
   HA_X1 i_8_0_582 (.A(\out_as[6] [4]), .B(n_8_0_581), .CO(n_8_0_582), .S());
   HA_X1 i_8_0_583 (.A(\out_as[6] [5]), .B(n_8_0_582), .CO(n_8_0_583), .S());
   HA_X1 i_8_0_584 (.A(\out_as[5] [2]), .B(n_8_0_1048), .CO(n_8_0_584), .S());
   HA_X1 i_8_0_585 (.A(\out_as[5] [3]), .B(n_8_0_584), .CO(n_8_0_585), .S());
   HA_X1 i_8_0_586 (.A(\out_as[5] [4]), .B(n_8_0_585), .CO(n_8_0_586), .S());
   HA_X1 i_8_0_587 (.A(\out_as[5] [5]), .B(n_8_0_586), .CO(n_8_0_587), .S());
   HA_X1 i_8_0_588 (.A(\out_as[4] [2]), .B(n_8_0_1174), .CO(n_8_0_588), .S());
   HA_X1 i_8_0_589 (.A(\out_as[4] [3]), .B(n_8_0_588), .CO(n_8_0_589), .S());
   HA_X1 i_8_0_590 (.A(\out_as[4] [4]), .B(n_8_0_589), .CO(n_8_0_590), .S());
   HA_X1 i_8_0_591 (.A(\out_as[4] [5]), .B(n_8_0_590), .CO(n_8_0_591), .S());
   HA_X1 i_8_0_592 (.A(\out_as[3] [2]), .B(n_8_0_1179), .CO(n_8_0_592), .S());
   HA_X1 i_8_0_593 (.A(\out_as[3] [3]), .B(n_8_0_592), .CO(n_8_0_593), .S());
   HA_X1 i_8_0_594 (.A(\out_as[3] [4]), .B(n_8_0_593), .CO(n_8_0_594), .S());
   HA_X1 i_8_0_595 (.A(\out_as[3] [5]), .B(n_8_0_594), .CO(n_8_0_595), .S());
   HA_X1 i_8_0_596 (.A(\out_as[2] [2]), .B(n_8_0_1168), .CO(n_8_0_596), .S());
   HA_X1 i_8_0_597 (.A(\out_as[2] [3]), .B(n_8_0_596), .CO(n_8_0_597), .S());
   HA_X1 i_8_0_598 (.A(\out_as[2] [4]), .B(n_8_0_597), .CO(n_8_0_598), .S());
   HA_X1 i_8_0_599 (.A(\out_as[2] [5]), .B(n_8_0_598), .CO(n_8_0_599), .S());
   HA_X1 i_8_0_600 (.A(\out_as[1] [2]), .B(n_8_0_1171), .CO(n_8_0_600), .S());
   HA_X1 i_8_0_601 (.A(\out_as[1] [3]), .B(n_8_0_600), .CO(n_8_0_601), .S());
   HA_X1 i_8_0_602 (.A(\out_as[1] [4]), .B(n_8_0_601), .CO(n_8_0_602), .S());
   HA_X1 i_8_0_603 (.A(\out_as[1] [5]), .B(n_8_0_602), .CO(n_8_0_603), .S());
   HA_X1 i_8_0_604 (.A(\out_as[0] [2]), .B(n_8_0_1176), .CO(n_8_0_604), .S());
   HA_X1 i_8_0_605 (.A(\out_as[0] [3]), .B(n_8_0_604), .CO(n_8_0_605), .S());
   HA_X1 i_8_0_606 (.A(\out_as[0] [4]), .B(n_8_0_605), .CO(n_8_0_606), .S());
   HA_X1 i_8_0_607 (.A(\out_as[0] [5]), .B(n_8_0_606), .CO(n_8_0_607), .S());
   HA_X1 i_8_0_608 (.A(\out_as[7] [3]), .B(\out_as[7] [2]), .CO(n_8_0_608), 
      .S());
   HA_X1 i_8_0_609 (.A(\out_as[7] [4]), .B(n_8_0_608), .CO(n_8_0_609), .S());
   HA_X1 i_8_0_610 (.A(\out_as[7] [5]), .B(n_8_0_609), .CO(n_8_0_610), .S());
   HA_X1 i_8_0_611 (.A(\out_as[6] [3]), .B(\out_as[6] [2]), .CO(n_8_0_611), 
      .S());
   HA_X1 i_8_0_612 (.A(\out_as[6] [4]), .B(n_8_0_611), .CO(n_8_0_612), .S());
   HA_X1 i_8_0_613 (.A(\out_as[6] [5]), .B(n_8_0_612), .CO(n_8_0_613), .S());
   HA_X1 i_8_0_614 (.A(\out_as[5] [3]), .B(\out_as[5] [2]), .CO(n_8_0_614), 
      .S());
   HA_X1 i_8_0_615 (.A(\out_as[5] [4]), .B(n_8_0_614), .CO(n_8_0_615), .S());
   HA_X1 i_8_0_616 (.A(\out_as[5] [5]), .B(n_8_0_615), .CO(n_8_0_616), .S());
   HA_X1 i_8_0_617 (.A(\out_as[4] [3]), .B(\out_as[4] [2]), .CO(n_8_0_617), 
      .S());
   HA_X1 i_8_0_618 (.A(\out_as[4] [4]), .B(n_8_0_617), .CO(n_8_0_618), .S());
   HA_X1 i_8_0_619 (.A(\out_as[4] [5]), .B(n_8_0_618), .CO(n_8_0_619), .S());
   HA_X1 i_8_0_620 (.A(\out_as[3] [3]), .B(\out_as[3] [2]), .CO(n_8_0_620), 
      .S());
   HA_X1 i_8_0_621 (.A(\out_as[3] [4]), .B(n_8_0_620), .CO(n_8_0_621), .S());
   HA_X1 i_8_0_622 (.A(\out_as[3] [5]), .B(n_8_0_621), .CO(n_8_0_622), .S());
   HA_X1 i_8_0_623 (.A(\out_as[2] [3]), .B(\out_as[2] [2]), .CO(n_8_0_623), 
      .S());
   HA_X1 i_8_0_624 (.A(\out_as[2] [4]), .B(n_8_0_623), .CO(n_8_0_624), .S());
   HA_X1 i_8_0_625 (.A(\out_as[2] [5]), .B(n_8_0_624), .CO(n_8_0_625), .S());
   HA_X1 i_8_0_626 (.A(\out_as[1] [3]), .B(\out_as[1] [2]), .CO(n_8_0_626), 
      .S());
   HA_X1 i_8_0_627 (.A(\out_as[1] [4]), .B(n_8_0_626), .CO(n_8_0_627), .S());
   HA_X1 i_8_0_628 (.A(\out_as[1] [5]), .B(n_8_0_627), .CO(n_8_0_628), .S());
   HA_X1 i_8_0_629 (.A(\out_as[0] [3]), .B(\out_as[0] [2]), .CO(n_8_0_629), 
      .S());
   HA_X1 i_8_0_630 (.A(\out_as[0] [4]), .B(n_8_0_629), .CO(n_8_0_630), .S());
   HA_X1 i_8_0_631 (.A(\out_as[0] [5]), .B(n_8_0_630), .CO(n_8_0_631), .S());
   HA_X1 i_8_0_632 (.A(\out_as[7] [3]), .B(n_8_0_1212), .CO(n_8_0_632), .S());
   HA_X1 i_8_0_633 (.A(\out_as[7] [4]), .B(n_8_0_632), .CO(n_8_0_633), .S());
   HA_X1 i_8_0_634 (.A(\out_as[7] [5]), .B(n_8_0_633), .CO(n_8_0_634), .S());
   HA_X1 i_8_0_635 (.A(\out_as[6] [3]), .B(n_8_0_1206), .CO(n_8_0_635), .S());
   HA_X1 i_8_0_636 (.A(\out_as[6] [4]), .B(n_8_0_635), .CO(n_8_0_636), .S());
   HA_X1 i_8_0_637 (.A(\out_as[6] [5]), .B(n_8_0_636), .CO(n_8_0_637), .S());
   HA_X1 i_8_0_638 (.A(\out_as[5] [3]), .B(n_8_0_1210), .CO(n_8_0_638), .S());
   HA_X1 i_8_0_639 (.A(\out_as[5] [4]), .B(n_8_0_638), .CO(n_8_0_639), .S());
   HA_X1 i_8_0_640 (.A(\out_as[5] [5]), .B(n_8_0_639), .CO(n_8_0_640), .S());
   HA_X1 i_8_0_641 (.A(\out_as[4] [3]), .B(n_8_0_1204), .CO(n_8_0_641), .S());
   HA_X1 i_8_0_642 (.A(\out_as[4] [4]), .B(n_8_0_641), .CO(n_8_0_642), .S());
   HA_X1 i_8_0_643 (.A(\out_as[4] [5]), .B(n_8_0_642), .CO(n_8_0_643), .S());
   HA_X1 i_8_0_644 (.A(\out_as[3] [3]), .B(n_8_0_1213), .CO(n_8_0_644), .S());
   HA_X1 i_8_0_645 (.A(\out_as[3] [4]), .B(n_8_0_644), .CO(n_8_0_645), .S());
   HA_X1 i_8_0_646 (.A(\out_as[3] [5]), .B(n_8_0_645), .CO(n_8_0_646), .S());
   HA_X1 i_8_0_647 (.A(\out_as[2] [3]), .B(n_8_0_1119), .CO(n_8_0_647), .S());
   HA_X1 i_8_0_648 (.A(\out_as[2] [4]), .B(n_8_0_647), .CO(n_8_0_648), .S());
   HA_X1 i_8_0_649 (.A(\out_as[2] [5]), .B(n_8_0_648), .CO(n_8_0_649), .S());
   HA_X1 i_8_0_650 (.A(\out_as[1] [3]), .B(n_8_0_1208), .CO(n_8_0_650), .S());
   HA_X1 i_8_0_651 (.A(\out_as[1] [4]), .B(n_8_0_650), .CO(n_8_0_651), .S());
   HA_X1 i_8_0_652 (.A(\out_as[1] [5]), .B(n_8_0_651), .CO(n_8_0_652), .S());
   HA_X1 i_8_0_653 (.A(\out_as[0] [3]), .B(n_8_0_1203), .CO(n_8_0_653), .S());
   HA_X1 i_8_0_654 (.A(\out_as[0] [4]), .B(n_8_0_653), .CO(n_8_0_654), .S());
   HA_X1 i_8_0_655 (.A(\out_as[0] [5]), .B(n_8_0_654), .CO(n_8_0_655), .S());
   HA_X1 i_8_0_656 (.A(\out_as[7] [3]), .B(n_8_0_1193), .CO(n_8_0_656), .S());
   HA_X1 i_8_0_657 (.A(\out_as[7] [4]), .B(n_8_0_656), .CO(n_8_0_657), .S());
   HA_X1 i_8_0_658 (.A(\out_as[7] [5]), .B(n_8_0_657), .CO(n_8_0_658), .S());
   HA_X1 i_8_0_659 (.A(\out_as[6] [3]), .B(n_8_0_1185), .CO(n_8_0_659), .S());
   HA_X1 i_8_0_660 (.A(\out_as[6] [4]), .B(n_8_0_659), .CO(n_8_0_660), .S());
   HA_X1 i_8_0_661 (.A(\out_as[6] [5]), .B(n_8_0_660), .CO(n_8_0_661), .S());
   HA_X1 i_8_0_662 (.A(\out_as[5] [3]), .B(n_8_0_1201), .CO(n_8_0_662), .S());
   HA_X1 i_8_0_663 (.A(\out_as[5] [4]), .B(n_8_0_662), .CO(n_8_0_663), .S());
   HA_X1 i_8_0_664 (.A(\out_as[5] [5]), .B(n_8_0_663), .CO(n_8_0_664), .S());
   HA_X1 i_8_0_665 (.A(\out_as[4] [3]), .B(n_8_0_1188), .CO(n_8_0_665), .S());
   HA_X1 i_8_0_666 (.A(\out_as[4] [4]), .B(n_8_0_665), .CO(n_8_0_666), .S());
   HA_X1 i_8_0_667 (.A(\out_as[4] [5]), .B(n_8_0_666), .CO(n_8_0_667), .S());
   HA_X1 i_8_0_668 (.A(\out_as[3] [3]), .B(n_8_0_1187), .CO(n_8_0_668), .S());
   HA_X1 i_8_0_669 (.A(\out_as[3] [4]), .B(n_8_0_668), .CO(n_8_0_669), .S());
   HA_X1 i_8_0_670 (.A(\out_as[3] [5]), .B(n_8_0_669), .CO(n_8_0_670), .S());
   HA_X1 i_8_0_671 (.A(\out_as[2] [3]), .B(n_8_0_1195), .CO(n_8_0_671), .S());
   HA_X1 i_8_0_672 (.A(\out_as[2] [4]), .B(n_8_0_671), .CO(n_8_0_672), .S());
   HA_X1 i_8_0_673 (.A(\out_as[2] [5]), .B(n_8_0_672), .CO(n_8_0_673), .S());
   HA_X1 i_8_0_674 (.A(\out_as[1] [3]), .B(n_8_0_1197), .CO(n_8_0_674), .S());
   HA_X1 i_8_0_675 (.A(\out_as[1] [4]), .B(n_8_0_674), .CO(n_8_0_675), .S());
   HA_X1 i_8_0_676 (.A(\out_as[1] [5]), .B(n_8_0_675), .CO(n_8_0_676), .S());
   HA_X1 i_8_0_677 (.A(\out_as[0] [3]), .B(n_8_0_1191), .CO(n_8_0_677), .S());
   HA_X1 i_8_0_678 (.A(\out_as[0] [4]), .B(n_8_0_677), .CO(n_8_0_678), .S());
   HA_X1 i_8_0_679 (.A(\out_as[0] [5]), .B(n_8_0_678), .CO(n_8_0_679), .S());
   HA_X1 i_8_0_680 (.A(\out_as[7] [3]), .B(n_8_0_1182), .CO(n_8_0_680), .S());
   HA_X1 i_8_0_681 (.A(\out_as[7] [4]), .B(n_8_0_680), .CO(n_8_0_681), .S());
   HA_X1 i_8_0_682 (.A(\out_as[7] [5]), .B(n_8_0_681), .CO(n_8_0_682), .S());
   HA_X1 i_8_0_683 (.A(\out_as[6] [3]), .B(n_8_0_975), .CO(n_8_0_683), .S());
   HA_X1 i_8_0_684 (.A(\out_as[6] [4]), .B(n_8_0_683), .CO(n_8_0_684), .S());
   HA_X1 i_8_0_685 (.A(\out_as[6] [5]), .B(n_8_0_684), .CO(n_8_0_685), .S());
   HA_X1 i_8_0_686 (.A(\out_as[5] [3]), .B(n_8_0_1047), .CO(n_8_0_686), .S());
   HA_X1 i_8_0_687 (.A(\out_as[5] [4]), .B(n_8_0_686), .CO(n_8_0_687), .S());
   HA_X1 i_8_0_688 (.A(\out_as[5] [5]), .B(n_8_0_687), .CO(n_8_0_688), .S());
   HA_X1 i_8_0_689 (.A(\out_as[4] [3]), .B(n_8_0_1173), .CO(n_8_0_689), .S());
   HA_X1 i_8_0_690 (.A(\out_as[4] [4]), .B(n_8_0_689), .CO(n_8_0_690), .S());
   HA_X1 i_8_0_691 (.A(\out_as[4] [5]), .B(n_8_0_690), .CO(n_8_0_691), .S());
   HA_X1 i_8_0_692 (.A(\out_as[3] [3]), .B(n_8_0_1178), .CO(n_8_0_692), .S());
   HA_X1 i_8_0_693 (.A(\out_as[3] [4]), .B(n_8_0_692), .CO(n_8_0_693), .S());
   HA_X1 i_8_0_694 (.A(\out_as[3] [5]), .B(n_8_0_693), .CO(n_8_0_694), .S());
   HA_X1 i_8_0_695 (.A(\out_as[2] [3]), .B(n_8_0_974), .CO(n_8_0_695), .S());
   HA_X1 i_8_0_696 (.A(\out_as[2] [4]), .B(n_8_0_695), .CO(n_8_0_696), .S());
   HA_X1 i_8_0_697 (.A(\out_as[2] [5]), .B(n_8_0_696), .CO(n_8_0_697), .S());
   HA_X1 i_8_0_698 (.A(\out_as[1] [3]), .B(n_8_0_1170), .CO(n_8_0_698), .S());
   HA_X1 i_8_0_699 (.A(\out_as[1] [4]), .B(n_8_0_698), .CO(n_8_0_699), .S());
   HA_X1 i_8_0_700 (.A(\out_as[1] [5]), .B(n_8_0_699), .CO(n_8_0_700), .S());
   HA_X1 i_8_0_701 (.A(\out_as[0] [3]), .B(n_8_0_973), .CO(n_8_0_701), .S());
   HA_X1 i_8_0_702 (.A(\out_as[0] [4]), .B(n_8_0_701), .CO(n_8_0_702), .S());
   HA_X1 i_8_0_703 (.A(\out_as[0] [5]), .B(n_8_0_702), .CO(n_8_0_703), .S());
   HA_X1 i_8_0_704 (.A(\out_as[7] [4]), .B(\out_as[7] [3]), .CO(n_8_0_704), 
      .S());
   HA_X1 i_8_0_705 (.A(\out_as[7] [5]), .B(n_8_0_704), .CO(n_8_0_705), .S());
   HA_X1 i_8_0_706 (.A(\out_as[6] [4]), .B(\out_as[6] [3]), .CO(n_8_0_706), 
      .S());
   HA_X1 i_8_0_707 (.A(\out_as[6] [5]), .B(n_8_0_706), .CO(n_8_0_707), .S());
   HA_X1 i_8_0_708 (.A(\out_as[5] [4]), .B(\out_as[5] [3]), .CO(n_8_0_708), 
      .S());
   HA_X1 i_8_0_709 (.A(\out_as[5] [5]), .B(n_8_0_708), .CO(n_8_0_709), .S());
   HA_X1 i_8_0_710 (.A(\out_as[4] [4]), .B(\out_as[4] [3]), .CO(n_8_0_710), 
      .S());
   HA_X1 i_8_0_711 (.A(\out_as[4] [5]), .B(n_8_0_710), .CO(n_8_0_711), .S());
   HA_X1 i_8_0_712 (.A(\out_as[3] [4]), .B(\out_as[3] [3]), .CO(n_8_0_712), 
      .S());
   HA_X1 i_8_0_713 (.A(\out_as[3] [5]), .B(n_8_0_712), .CO(n_8_0_713), .S());
   HA_X1 i_8_0_714 (.A(\out_as[2] [4]), .B(\out_as[2] [3]), .CO(n_8_0_714), 
      .S());
   HA_X1 i_8_0_715 (.A(\out_as[2] [5]), .B(n_8_0_714), .CO(n_8_0_715), .S());
   HA_X1 i_8_0_716 (.A(\out_as[1] [4]), .B(\out_as[1] [3]), .CO(n_8_0_716), 
      .S());
   HA_X1 i_8_0_717 (.A(\out_as[1] [5]), .B(n_8_0_716), .CO(n_8_0_717), .S());
   HA_X1 i_8_0_718 (.A(\out_as[0] [4]), .B(\out_as[0] [3]), .CO(n_8_0_718), 
      .S());
   HA_X1 i_8_0_719 (.A(\out_as[0] [5]), .B(n_8_0_718), .CO(n_8_0_719), .S());
   HA_X1 i_8_0_720 (.A(\out_as[7] [4]), .B(n_8_0_1286), .CO(n_8_0_720), .S());
   HA_X1 i_8_0_721 (.A(\out_as[7] [5]), .B(n_8_0_720), .CO(n_8_0_721), .S());
   HA_X1 i_8_0_722 (.A(\out_as[6] [4]), .B(n_8_0_1273), .CO(n_8_0_722), .S());
   HA_X1 i_8_0_723 (.A(\out_as[6] [5]), .B(n_8_0_722), .CO(n_8_0_723), .S());
   HA_X1 i_8_0_724 (.A(\out_as[5] [4]), .B(n_8_0_1276), .CO(n_8_0_724), .S());
   HA_X1 i_8_0_725 (.A(\out_as[5] [5]), .B(n_8_0_724), .CO(n_8_0_725), .S());
   HA_X1 i_8_0_726 (.A(\out_as[4] [4]), .B(n_8_0_1269), .CO(n_8_0_726), .S());
   HA_X1 i_8_0_727 (.A(\out_as[4] [5]), .B(n_8_0_726), .CO(n_8_0_727), .S());
   HA_X1 i_8_0_728 (.A(\out_as[3] [4]), .B(n_8_0_1288), .CO(n_8_0_728), .S());
   HA_X1 i_8_0_729 (.A(\out_as[3] [5]), .B(n_8_0_728), .CO(n_8_0_729), .S());
   HA_X1 i_8_0_730 (.A(\out_as[2] [4]), .B(n_8_0_1284), .CO(n_8_0_730), .S());
   HA_X1 i_8_0_731 (.A(\out_as[2] [5]), .B(n_8_0_730), .CO(n_8_0_731), .S());
   HA_X1 i_8_0_732 (.A(\out_as[1] [4]), .B(n_8_0_1281), .CO(n_8_0_732), .S());
   HA_X1 i_8_0_733 (.A(\out_as[1] [5]), .B(n_8_0_732), .CO(n_8_0_733), .S());
   HA_X1 i_8_0_734 (.A(\out_as[0] [4]), .B(n_8_0_1278), .CO(n_8_0_734), .S());
   HA_X1 i_8_0_735 (.A(\out_as[0] [5]), .B(n_8_0_734), .CO(n_8_0_735), .S());
   HA_X1 i_8_0_736 (.A(\out_as[7] [4]), .B(n_8_0_1262), .CO(n_8_0_736), .S());
   HA_X1 i_8_0_737 (.A(\out_as[7] [5]), .B(n_8_0_736), .CO(n_8_0_737), .S());
   HA_X1 i_8_0_738 (.A(\out_as[6] [4]), .B(n_8_0_1261), .CO(n_8_0_738), .S());
   HA_X1 i_8_0_739 (.A(\out_as[6] [5]), .B(n_8_0_738), .CO(n_8_0_739), .S());
   HA_X1 i_8_0_740 (.A(\out_as[5] [4]), .B(n_8_0_1258), .CO(n_8_0_740), .S());
   HA_X1 i_8_0_741 (.A(\out_as[5] [5]), .B(n_8_0_740), .CO(n_8_0_741), .S());
   HA_X1 i_8_0_742 (.A(\out_as[4] [4]), .B(n_8_0_1252), .CO(n_8_0_742), .S());
   HA_X1 i_8_0_743 (.A(\out_as[4] [5]), .B(n_8_0_742), .CO(n_8_0_743), .S());
   HA_X1 i_8_0_744 (.A(\out_as[3] [4]), .B(n_8_0_1256), .CO(n_8_0_744), .S());
   HA_X1 i_8_0_745 (.A(\out_as[3] [5]), .B(n_8_0_744), .CO(n_8_0_745), .S());
   HA_X1 i_8_0_746 (.A(\out_as[2] [4]), .B(n_8_0_1264), .CO(n_8_0_746), .S());
   HA_X1 i_8_0_747 (.A(\out_as[2] [5]), .B(n_8_0_746), .CO(n_8_0_747), .S());
   HA_X1 i_8_0_748 (.A(\out_as[1] [4]), .B(n_8_0_1267), .CO(n_8_0_748), .S());
   HA_X1 i_8_0_749 (.A(\out_as[1] [5]), .B(n_8_0_748), .CO(n_8_0_749), .S());
   HA_X1 i_8_0_750 (.A(\out_as[0] [4]), .B(n_8_0_1251), .CO(n_8_0_750), .S());
   HA_X1 i_8_0_751 (.A(\out_as[0] [5]), .B(n_8_0_750), .CO(n_8_0_751), .S());
   HA_X1 i_8_0_752 (.A(\out_as[7] [4]), .B(n_8_0_1240), .CO(n_8_0_752), .S());
   HA_X1 i_8_0_753 (.A(\out_as[7] [5]), .B(n_8_0_752), .CO(n_8_0_753), .S());
   HA_X1 i_8_0_754 (.A(\out_as[6] [4]), .B(n_8_0_1247), .CO(n_8_0_754), .S());
   HA_X1 i_8_0_755 (.A(\out_as[6] [5]), .B(n_8_0_754), .CO(n_8_0_755), .S());
   HA_X1 i_8_0_756 (.A(\out_as[5] [4]), .B(n_8_0_1238), .CO(n_8_0_756), .S());
   HA_X1 i_8_0_757 (.A(\out_as[5] [5]), .B(n_8_0_756), .CO(n_8_0_757), .S());
   HA_X1 i_8_0_758 (.A(\out_as[4] [4]), .B(n_8_0_1236), .CO(n_8_0_758), .S());
   HA_X1 i_8_0_759 (.A(\out_as[4] [5]), .B(n_8_0_758), .CO(n_8_0_759), .S());
   HA_X1 i_8_0_760 (.A(\out_as[3] [4]), .B(n_8_0_1250), .CO(n_8_0_760), .S());
   HA_X1 i_8_0_761 (.A(\out_as[3] [5]), .B(n_8_0_760), .CO(n_8_0_761), .S());
   HA_X1 i_8_0_762 (.A(\out_as[2] [4]), .B(n_8_0_1241), .CO(n_8_0_762), .S());
   HA_X1 i_8_0_763 (.A(\out_as[2] [5]), .B(n_8_0_762), .CO(n_8_0_763), .S());
   HA_X1 i_8_0_764 (.A(\out_as[1] [4]), .B(n_8_0_1242), .CO(n_8_0_764), .S());
   HA_X1 i_8_0_765 (.A(\out_as[1] [5]), .B(n_8_0_764), .CO(n_8_0_765), .S());
   HA_X1 i_8_0_766 (.A(\out_as[0] [4]), .B(n_8_0_1244), .CO(n_8_0_766), .S());
   HA_X1 i_8_0_767 (.A(\out_as[0] [5]), .B(n_8_0_766), .CO(n_8_0_767), .S());
   HA_X1 i_8_0_768 (.A(\out_as[7] [4]), .B(n_8_0_1226), .CO(n_8_0_768), .S());
   HA_X1 i_8_0_769 (.A(\out_as[7] [5]), .B(n_8_0_768), .CO(n_8_0_769), .S());
   HA_X1 i_8_0_770 (.A(\out_as[6] [4]), .B(n_8_0_1221), .CO(n_8_0_770), .S());
   HA_X1 i_8_0_771 (.A(\out_as[6] [5]), .B(n_8_0_770), .CO(n_8_0_771), .S());
   HA_X1 i_8_0_772 (.A(\out_as[5] [4]), .B(n_8_0_1218), .CO(n_8_0_772), .S());
   HA_X1 i_8_0_773 (.A(\out_as[5] [5]), .B(n_8_0_772), .CO(n_8_0_773), .S());
   HA_X1 i_8_0_774 (.A(\out_as[4] [4]), .B(n_8_0_1233), .CO(n_8_0_774), .S());
   HA_X1 i_8_0_775 (.A(\out_as[4] [5]), .B(n_8_0_774), .CO(n_8_0_775), .S());
   HA_X1 i_8_0_776 (.A(\out_as[3] [4]), .B(n_8_0_1214), .CO(n_8_0_776), .S());
   HA_X1 i_8_0_777 (.A(\out_as[3] [5]), .B(n_8_0_776), .CO(n_8_0_777), .S());
   HA_X1 i_8_0_778 (.A(\out_as[2] [4]), .B(n_8_0_1224), .CO(n_8_0_778), .S());
   HA_X1 i_8_0_779 (.A(\out_as[2] [5]), .B(n_8_0_778), .CO(n_8_0_779), .S());
   HA_X1 i_8_0_780 (.A(\out_as[1] [4]), .B(n_8_0_1231), .CO(n_8_0_780), .S());
   HA_X1 i_8_0_781 (.A(\out_as[1] [5]), .B(n_8_0_780), .CO(n_8_0_781), .S());
   HA_X1 i_8_0_782 (.A(\out_as[0] [4]), .B(n_8_0_1228), .CO(n_8_0_782), .S());
   HA_X1 i_8_0_783 (.A(\out_as[0] [5]), .B(n_8_0_782), .CO(n_8_0_783), .S());
   HA_X1 i_8_0_784 (.A(\out_as[7] [4]), .B(n_8_0_1211), .CO(n_8_0_784), .S());
   HA_X1 i_8_0_785 (.A(\out_as[7] [5]), .B(n_8_0_784), .CO(n_8_0_785), .S());
   HA_X1 i_8_0_786 (.A(\out_as[6] [4]), .B(n_8_0_1205), .CO(n_8_0_786), .S());
   HA_X1 i_8_0_787 (.A(\out_as[6] [5]), .B(n_8_0_786), .CO(n_8_0_787), .S());
   HA_X1 i_8_0_788 (.A(\out_as[5] [4]), .B(n_8_0_1209), .CO(n_8_0_788), .S());
   HA_X1 i_8_0_789 (.A(\out_as[5] [5]), .B(n_8_0_788), .CO(n_8_0_789), .S());
   HA_X1 i_8_0_790 (.A(\out_as[4] [4]), .B(n_8_0_972), .CO(n_8_0_790), .S());
   HA_X1 i_8_0_791 (.A(\out_as[4] [5]), .B(n_8_0_790), .CO(n_8_0_791), .S());
   HA_X1 i_8_0_792 (.A(\out_as[3] [4]), .B(n_8_0_971), .CO(n_8_0_792), .S());
   HA_X1 i_8_0_793 (.A(\out_as[3] [5]), .B(n_8_0_792), .CO(n_8_0_793), .S());
   HA_X1 i_8_0_794 (.A(\out_as[2] [4]), .B(n_8_0_1118), .CO(n_8_0_794), .S());
   HA_X1 i_8_0_795 (.A(\out_as[2] [5]), .B(n_8_0_794), .CO(n_8_0_795), .S());
   HA_X1 i_8_0_796 (.A(\out_as[1] [4]), .B(n_8_0_1207), .CO(n_8_0_796), .S());
   HA_X1 i_8_0_797 (.A(\out_as[1] [5]), .B(n_8_0_796), .CO(n_8_0_797), .S());
   HA_X1 i_8_0_798 (.A(\out_as[0] [4]), .B(n_8_0_1163), .CO(n_8_0_798), .S());
   HA_X1 i_8_0_799 (.A(\out_as[0] [5]), .B(n_8_0_798), .CO(n_8_0_799), .S());
   HA_X1 i_8_0_800 (.A(\out_as[7] [4]), .B(n_8_0_1192), .CO(n_8_0_800), .S());
   HA_X1 i_8_0_801 (.A(\out_as[7] [5]), .B(n_8_0_800), .CO(n_8_0_801), .S());
   HA_X1 i_8_0_802 (.A(\out_as[6] [4]), .B(n_8_0_1184), .CO(n_8_0_802), .S());
   HA_X1 i_8_0_803 (.A(\out_as[6] [5]), .B(n_8_0_802), .CO(n_8_0_803), .S());
   HA_X1 i_8_0_804 (.A(\out_as[5] [4]), .B(n_8_0_1200), .CO(n_8_0_804), .S());
   HA_X1 i_8_0_805 (.A(\out_as[5] [5]), .B(n_8_0_804), .CO(n_8_0_805), .S());
   HA_X1 i_8_0_806 (.A(\out_as[4] [4]), .B(n_8_0_970), .CO(n_8_0_806), .S());
   HA_X1 i_8_0_807 (.A(\out_as[4] [5]), .B(n_8_0_806), .CO(n_8_0_807), .S());
   HA_X1 i_8_0_808 (.A(\out_as[3] [4]), .B(n_8_0_1186), .CO(n_8_0_808), .S());
   HA_X1 i_8_0_809 (.A(\out_as[3] [5]), .B(n_8_0_808), .CO(n_8_0_809), .S());
   HA_X1 i_8_0_810 (.A(\out_as[2] [4]), .B(n_8_0_1194), .CO(n_8_0_810), .S());
   HA_X1 i_8_0_811 (.A(\out_as[2] [5]), .B(n_8_0_810), .CO(n_8_0_811), .S());
   HA_X1 i_8_0_812 (.A(\out_as[1] [4]), .B(n_8_0_1196), .CO(n_8_0_812), .S());
   HA_X1 i_8_0_813 (.A(\out_as[1] [5]), .B(n_8_0_812), .CO(n_8_0_813), .S());
   HA_X1 i_8_0_814 (.A(\out_as[0] [4]), .B(n_8_0_1190), .CO(n_8_0_814), .S());
   HA_X1 i_8_0_815 (.A(\out_as[0] [5]), .B(n_8_0_814), .CO(n_8_0_815), .S());
   HA_X1 i_8_0_816 (.A(\out_as[7] [4]), .B(n_8_0_1001), .CO(n_8_0_816), .S());
   HA_X1 i_8_0_817 (.A(\out_as[7] [5]), .B(n_8_0_816), .CO(n_8_0_817), .S());
   HA_X1 i_8_0_818 (.A(\out_as[6] [4]), .B(n_8_0_1180), .CO(n_8_0_818), .S());
   HA_X1 i_8_0_819 (.A(\out_as[6] [5]), .B(n_8_0_818), .CO(n_8_0_819), .S());
   HA_X1 i_8_0_820 (.A(\out_as[5] [4]), .B(n_8_0_969), .CO(n_8_0_820), .S());
   HA_X1 i_8_0_821 (.A(\out_as[5] [5]), .B(n_8_0_820), .CO(n_8_0_821), .S());
   HA_X1 i_8_0_822 (.A(\out_as[4] [4]), .B(n_8_0_1172), .CO(n_8_0_822), .S());
   HA_X1 i_8_0_823 (.A(\out_as[4] [5]), .B(n_8_0_822), .CO(n_8_0_823), .S());
   HA_X1 i_8_0_824 (.A(\out_as[3] [4]), .B(n_8_0_1177), .CO(n_8_0_824), .S());
   HA_X1 i_8_0_825 (.A(\out_as[3] [5]), .B(n_8_0_824), .CO(n_8_0_825), .S());
   HA_X1 i_8_0_826 (.A(\out_as[2] [4]), .B(n_8_0_1167), .CO(n_8_0_826), .S());
   HA_X1 i_8_0_827 (.A(\out_as[2] [5]), .B(n_8_0_826), .CO(n_8_0_827), .S());
   HA_X1 i_8_0_828 (.A(\out_as[1] [4]), .B(n_8_0_1169), .CO(n_8_0_828), .S());
   HA_X1 i_8_0_829 (.A(\out_as[1] [5]), .B(n_8_0_828), .CO(n_8_0_829), .S());
   HA_X1 i_8_0_830 (.A(\out_as[0] [4]), .B(n_8_0_1175), .CO(n_8_0_830), .S());
   HA_X1 i_8_0_831 (.A(\out_as[0] [5]), .B(n_8_0_830), .CO(n_8_0_831), .S());
   HA_X1 i_8_0_832 (.A(\out_as[7] [5]), .B(\out_as[7] [4]), .CO(n_8_0_832), 
      .S());
   HA_X1 i_8_0_833 (.A(\out_as[6] [5]), .B(\out_as[6] [4]), .CO(n_8_0_833), 
      .S());
   HA_X1 i_8_0_834 (.A(\out_as[5] [5]), .B(\out_as[5] [4]), .CO(n_8_0_834), 
      .S());
   HA_X1 i_8_0_835 (.A(\out_as[4] [5]), .B(\out_as[4] [4]), .CO(n_8_0_835), 
      .S());
   HA_X1 i_8_0_836 (.A(\out_as[3] [5]), .B(\out_as[3] [4]), .CO(n_8_0_836), 
      .S());
   HA_X1 i_8_0_837 (.A(\out_as[2] [5]), .B(\out_as[2] [4]), .CO(n_8_0_837), 
      .S());
   HA_X1 i_8_0_838 (.A(\out_as[1] [5]), .B(\out_as[1] [4]), .CO(n_8_0_838), 
      .S());
   HA_X1 i_8_0_839 (.A(\out_as[0] [5]), .B(\out_as[0] [4]), .CO(n_8_0_839), 
      .S());
   HA_X1 i_8_0_840 (.A(\out_as[7] [5]), .B(n_8_0_1352), .CO(n_8_0_840), .S());
   HA_X1 i_8_0_841 (.A(\out_as[6] [5]), .B(n_8_0_1348), .CO(n_8_0_841), .S());
   HA_X1 i_8_0_842 (.A(\out_as[5] [5]), .B(n_8_0_1345), .CO(n_8_0_842), .S());
   HA_X1 i_8_0_843 (.A(\out_as[4] [5]), .B(n_8_0_1346), .CO(n_8_0_843), .S());
   HA_X1 i_8_0_844 (.A(\out_as[3] [5]), .B(n_8_0_1347), .CO(n_8_0_844), .S());
   HA_X1 i_8_0_845 (.A(\out_as[2] [5]), .B(n_8_0_1349), .CO(n_8_0_845), .S());
   HA_X1 i_8_0_846 (.A(\out_as[1] [5]), .B(n_8_0_1351), .CO(n_8_0_846), .S());
   HA_X1 i_8_0_847 (.A(\out_as[0] [5]), .B(n_8_0_1350), .CO(n_8_0_847), .S());
   HA_X1 i_8_0_848 (.A(\out_as[7] [5]), .B(n_8_0_1343), .CO(n_8_0_848), .S());
   HA_X1 i_8_0_849 (.A(\out_as[6] [5]), .B(n_8_0_1339), .CO(n_8_0_849), .S());
   HA_X1 i_8_0_850 (.A(\out_as[5] [5]), .B(n_8_0_1032), .CO(n_8_0_850), .S());
   HA_X1 i_8_0_851 (.A(\out_as[4] [5]), .B(n_8_0_1338), .CO(n_8_0_851), .S());
   HA_X1 i_8_0_852 (.A(\out_as[3] [5]), .B(n_8_0_1344), .CO(n_8_0_852), .S());
   HA_X1 i_8_0_853 (.A(\out_as[2] [5]), .B(n_8_0_1341), .CO(n_8_0_853), .S());
   HA_X1 i_8_0_854 (.A(\out_as[1] [5]), .B(n_8_0_1340), .CO(n_8_0_854), .S());
   HA_X1 i_8_0_855 (.A(\out_as[0] [5]), .B(n_8_0_1342), .CO(n_8_0_855), .S());
   HA_X1 i_8_0_856 (.A(\out_as[7] [5]), .B(n_8_0_1336), .CO(n_8_0_856), .S());
   HA_X1 i_8_0_857 (.A(\out_as[6] [5]), .B(n_8_0_1332), .CO(n_8_0_857), .S());
   HA_X1 i_8_0_858 (.A(\out_as[5] [5]), .B(n_8_0_1034), .CO(n_8_0_858), .S());
   HA_X1 i_8_0_859 (.A(\out_as[4] [5]), .B(n_8_0_1333), .CO(n_8_0_859), .S());
   HA_X1 i_8_0_860 (.A(\out_as[3] [5]), .B(n_8_0_1337), .CO(n_8_0_860), .S());
   HA_X1 i_8_0_861 (.A(\out_as[2] [5]), .B(n_8_0_1335), .CO(n_8_0_861), .S());
   HA_X1 i_8_0_862 (.A(\out_as[1] [5]), .B(n_8_0_1334), .CO(n_8_0_862), .S());
   HA_X1 i_8_0_863 (.A(\out_as[0] [5]), .B(n_8_0_1331), .CO(n_8_0_863), .S());
   HA_X1 i_8_0_864 (.A(\out_as[7] [5]), .B(n_8_0_1322), .CO(n_8_0_864), .S());
   HA_X1 i_8_0_865 (.A(\out_as[6] [5]), .B(n_8_0_1328), .CO(n_8_0_865), .S());
   HA_X1 i_8_0_866 (.A(\out_as[5] [5]), .B(n_8_0_1036), .CO(n_8_0_866), .S());
   HA_X1 i_8_0_867 (.A(\out_as[4] [5]), .B(n_8_0_1329), .CO(n_8_0_867), .S());
   HA_X1 i_8_0_868 (.A(\out_as[3] [5]), .B(n_8_0_1330), .CO(n_8_0_868), .S());
   HA_X1 i_8_0_869 (.A(\out_as[2] [5]), .B(n_8_0_1326), .CO(n_8_0_869), .S());
   HA_X1 i_8_0_870 (.A(\out_as[1] [5]), .B(n_8_0_1324), .CO(n_8_0_870), .S());
   HA_X1 i_8_0_871 (.A(\out_as[0] [5]), .B(n_8_0_1323), .CO(n_8_0_871), .S());
   HA_X1 i_8_0_872 (.A(\out_as[7] [5]), .B(n_8_0_1315), .CO(n_8_0_872), .S());
   HA_X1 i_8_0_873 (.A(\out_as[6] [5]), .B(n_8_0_1318), .CO(n_8_0_873), .S());
   HA_X1 i_8_0_874 (.A(\out_as[5] [5]), .B(n_8_0_1038), .CO(n_8_0_874), .S());
   HA_X1 i_8_0_875 (.A(\out_as[4] [5]), .B(n_8_0_1319), .CO(n_8_0_875), .S());
   HA_X1 i_8_0_876 (.A(\out_as[3] [5]), .B(n_8_0_1321), .CO(n_8_0_876), .S());
   HA_X1 i_8_0_877 (.A(\out_as[2] [5]), .B(n_8_0_1320), .CO(n_8_0_877), .S());
   HA_X1 i_8_0_878 (.A(\out_as[1] [5]), .B(n_8_0_1317), .CO(n_8_0_878), .S());
   HA_X1 i_8_0_879 (.A(\out_as[0] [5]), .B(n_8_0_1316), .CO(n_8_0_879), .S());
   HA_X1 i_8_0_880 (.A(\out_as[7] [5]), .B(n_8_0_1311), .CO(n_8_0_880), .S());
   HA_X1 i_8_0_881 (.A(\out_as[6] [5]), .B(n_8_0_1010), .CO(n_8_0_881), .S());
   HA_X1 i_8_0_882 (.A(\out_as[5] [5]), .B(n_8_0_1310), .CO(n_8_0_882), .S());
   HA_X1 i_8_0_883 (.A(\out_as[4] [5]), .B(n_8_0_1309), .CO(n_8_0_883), .S());
   HA_X1 i_8_0_884 (.A(\out_as[3] [5]), .B(n_8_0_1308), .CO(n_8_0_884), .S());
   HA_X1 i_8_0_885 (.A(\out_as[2] [5]), .B(n_8_0_1312), .CO(n_8_0_885), .S());
   HA_X1 i_8_0_886 (.A(\out_as[1] [5]), .B(n_8_0_1314), .CO(n_8_0_886), .S());
   HA_X1 i_8_0_887 (.A(\out_as[0] [5]), .B(n_8_0_1313), .CO(n_8_0_887), .S());
   HA_X1 i_8_0_888 (.A(\out_as[7] [5]), .B(n_8_0_1305), .CO(n_8_0_888), .S());
   HA_X1 i_8_0_889 (.A(\out_as[6] [5]), .B(n_8_0_1304), .CO(n_8_0_889), .S());
   HA_X1 i_8_0_890 (.A(\out_as[5] [5]), .B(n_8_0_1298), .CO(n_8_0_890), .S());
   HA_X1 i_8_0_891 (.A(\out_as[4] [5]), .B(n_8_0_1299), .CO(n_8_0_891), .S());
   HA_X1 i_8_0_892 (.A(\out_as[3] [5]), .B(n_8_0_1301), .CO(n_8_0_892), .S());
   HA_X1 i_8_0_893 (.A(\out_as[2] [5]), .B(n_8_0_1307), .CO(n_8_0_893), .S());
   HA_X1 i_8_0_894 (.A(\out_as[1] [5]), .B(n_8_0_1306), .CO(n_8_0_894), .S());
   HA_X1 i_8_0_895 (.A(\out_as[0] [5]), .B(n_8_0_1303), .CO(n_8_0_895), .S());
   HA_X1 i_8_0_896 (.A(\out_as[7] [5]), .B(n_8_0_1296), .CO(n_8_0_896), .S());
   HA_X1 i_8_0_897 (.A(\out_as[6] [5]), .B(n_8_0_1291), .CO(n_8_0_897), .S());
   HA_X1 i_8_0_898 (.A(\out_as[5] [5]), .B(n_8_0_1289), .CO(n_8_0_898), .S());
   HA_X1 i_8_0_899 (.A(\out_as[4] [5]), .B(n_8_0_1297), .CO(n_8_0_899), .S());
   HA_X1 i_8_0_900 (.A(\out_as[3] [5]), .B(n_8_0_1290), .CO(n_8_0_900), .S());
   HA_X1 i_8_0_901 (.A(\out_as[2] [5]), .B(n_8_0_1293), .CO(n_8_0_901), .S());
   HA_X1 i_8_0_902 (.A(\out_as[1] [5]), .B(n_8_0_1292), .CO(n_8_0_902), .S());
   HA_X1 i_8_0_903 (.A(\out_as[0] [5]), .B(n_8_0_1295), .CO(n_8_0_903), .S());
   HA_X1 i_8_0_904 (.A(\out_as[7] [5]), .B(n_8_0_1285), .CO(n_8_0_904), .S());
   HA_X1 i_8_0_905 (.A(\out_as[6] [5]), .B(n_8_0_1272), .CO(n_8_0_905), .S());
   HA_X1 i_8_0_906 (.A(\out_as[5] [5]), .B(n_8_0_1275), .CO(n_8_0_906), .S());
   HA_X1 i_8_0_907 (.A(\out_as[4] [5]), .B(n_8_0_1268), .CO(n_8_0_907), .S());
   HA_X1 i_8_0_908 (.A(\out_as[3] [5]), .B(n_8_0_1287), .CO(n_8_0_908), .S());
   HA_X1 i_8_0_909 (.A(\out_as[2] [5]), .B(n_8_0_1283), .CO(n_8_0_909), .S());
   HA_X1 i_8_0_910 (.A(\out_as[1] [5]), .B(n_8_0_1280), .CO(n_8_0_910), .S());
   HA_X1 i_8_0_911 (.A(\out_as[0] [5]), .B(n_8_0_1277), .CO(n_8_0_911), .S());
   HA_X1 i_8_0_912 (.A(\out_as[7] [5]), .B(n_8_0_991), .CO(n_8_0_912), .S());
   HA_X1 i_8_0_913 (.A(\out_as[6] [5]), .B(n_8_0_1260), .CO(n_8_0_913), .S());
   HA_X1 i_8_0_914 (.A(\out_as[5] [5]), .B(n_8_0_1257), .CO(n_8_0_914), .S());
   HA_X1 i_8_0_915 (.A(\out_as[4] [5]), .B(n_8_0_968), .CO(n_8_0_915), .S());
   HA_X1 i_8_0_916 (.A(\out_as[3] [5]), .B(n_8_0_1255), .CO(n_8_0_916), .S());
   HA_X1 i_8_0_917 (.A(\out_as[2] [5]), .B(n_8_0_1263), .CO(n_8_0_917), .S());
   HA_X1 i_8_0_918 (.A(\out_as[1] [5]), .B(n_8_0_1266), .CO(n_8_0_918), .S());
   HA_X1 i_8_0_919 (.A(\out_as[0] [5]), .B(n_8_0_967), .CO(n_8_0_919), .S());
   HA_X1 i_8_0_920 (.A(\out_as[7] [5]), .B(n_8_0_1239), .CO(n_8_0_920), .S());
   HA_X1 i_8_0_921 (.A(\out_as[6] [5]), .B(n_8_0_1246), .CO(n_8_0_921), .S());
   HA_X1 i_8_0_922 (.A(\out_as[5] [5]), .B(n_8_0_1237), .CO(n_8_0_922), .S());
   HA_X1 i_8_0_923 (.A(\out_as[4] [5]), .B(n_8_0_1235), .CO(n_8_0_923), .S());
   HA_X1 i_8_0_924 (.A(\out_as[3] [5]), .B(n_8_0_1249), .CO(n_8_0_924), .S());
   HA_X1 i_8_0_925 (.A(\out_as[2] [5]), .B(n_8_0_1116), .CO(n_8_0_925), .S());
   HA_X1 i_8_0_926 (.A(\out_as[1] [5]), .B(n_8_0_1137), .CO(n_8_0_926), .S());
   HA_X1 i_8_0_927 (.A(\out_as[0] [5]), .B(n_8_0_966), .CO(n_8_0_927), .S());
   HA_X1 i_8_0_928 (.A(\out_as[7] [5]), .B(n_8_0_1225), .CO(n_8_0_928), .S());
   HA_X1 i_8_0_929 (.A(\out_as[6] [5]), .B(n_8_0_1220), .CO(n_8_0_929), .S());
   HA_X1 i_8_0_930 (.A(\out_as[5] [5]), .B(n_8_0_1217), .CO(n_8_0_930), .S());
   HA_X1 i_8_0_931 (.A(\out_as[4] [5]), .B(n_8_0_1232), .CO(n_8_0_931), .S());
   HA_X1 i_8_0_932 (.A(\out_as[3] [5]), .B(n_8_0_1099), .CO(n_8_0_932), .S());
   HA_X1 i_8_0_933 (.A(\out_as[2] [5]), .B(n_8_0_1223), .CO(n_8_0_933), .S());
   HA_X1 i_8_0_934 (.A(\out_as[1] [5]), .B(n_8_0_1140), .CO(n_8_0_934), .S());
   HA_X1 i_8_0_935 (.A(\out_as[0] [5]), .B(n_8_0_1227), .CO(n_8_0_935), .S());
   HA_X1 i_8_0_936 (.A(\out_as[7] [5]), .B(n_8_0_995), .CO(n_8_0_936), .S());
   HA_X1 i_8_0_937 (.A(\out_as[6] [5]), .B(n_8_0_1013), .CO(n_8_0_937), .S());
   HA_X1 i_8_0_938 (.A(\out_as[5] [5]), .B(n_8_0_1044), .CO(n_8_0_938), .S());
   HA_X1 i_8_0_939 (.A(\out_as[4] [5]), .B(n_8_0_1069), .CO(n_8_0_939), .S());
   HA_X1 i_8_0_940 (.A(\out_as[3] [5]), .B(n_8_0_1094), .CO(n_8_0_940), .S());
   HA_X1 i_8_0_941 (.A(\out_as[2] [5]), .B(n_8_0_965), .CO(n_8_0_941), .S());
   HA_X1 i_8_0_942 (.A(\out_as[1] [5]), .B(n_8_0_1139), .CO(n_8_0_942), .S());
   HA_X1 i_8_0_943 (.A(\out_as[0] [5]), .B(n_8_0_1202), .CO(n_8_0_943), .S());
   HA_X1 i_8_0_944 (.A(\out_as[7] [5]), .B(n_8_0_997), .CO(n_8_0_944), .S());
   HA_X1 i_8_0_945 (.A(\out_as[6] [5]), .B(n_8_0_964), .CO(n_8_0_945), .S());
   HA_X1 i_8_0_946 (.A(\out_as[5] [5]), .B(n_8_0_1199), .CO(n_8_0_946), .S());
   HA_X1 i_8_0_947 (.A(\out_as[4] [5]), .B(n_8_0_1071), .CO(n_8_0_947), .S());
   HA_X1 i_8_0_948 (.A(\out_as[3] [5]), .B(n_8_0_1096), .CO(n_8_0_948), .S());
   HA_X1 i_8_0_949 (.A(\out_as[2] [5]), .B(n_8_0_1122), .CO(n_8_0_949), .S());
   HA_X1 i_8_0_950 (.A(\out_as[1] [5]), .B(n_8_0_1143), .CO(n_8_0_950), .S());
   HA_X1 i_8_0_951 (.A(\out_as[0] [5]), .B(n_8_0_1189), .CO(n_8_0_951), .S());
   HA_X1 i_8_0_952 (.A(\out_as[7] [5]), .B(n_8_0_1000), .CO(n_8_0_952), .S());
   HA_X1 i_8_0_953 (.A(\out_as[6] [5]), .B(n_8_0_963), .CO(n_8_0_953), .S());
   HA_X1 i_8_0_954 (.A(\out_as[5] [5]), .B(n_8_0_1046), .CO(n_8_0_954), .S());
   HA_X1 i_8_0_955 (.A(\out_as[4] [5]), .B(n_8_0_1073), .CO(n_8_0_955), .S());
   HA_X1 i_8_0_956 (.A(\out_as[3] [5]), .B(n_8_0_1098), .CO(n_8_0_956), .S());
   HA_X1 i_8_0_957 (.A(\out_as[2] [5]), .B(n_8_0_962), .CO(n_8_0_957), .S());
   HA_X1 i_8_0_958 (.A(\out_as[1] [5]), .B(n_8_0_961), .CO(n_8_0_958), .S());
   HA_X1 i_8_0_959 (.A(\out_as[0] [5]), .B(n_8_0_960), .CO(n_8_0_959), .S());
   NAND2_X1 i_8_0_960 (.A1(n_8_0_2835), .A2(n_8_0_2731), .ZN(n_8_0_960));
   NAND2_X1 i_8_0_961 (.A1(n_8_0_2970), .A2(n_8_0_2727), .ZN(n_8_0_961));
   NAND3_X1 i_8_0_962 (.A1(n_8_0_2829), .A2(n_8_0_2725), .A3(n_8_0_7064), 
      .ZN(n_8_0_962));
   NAND3_X1 i_8_0_963 (.A1(n_8_0_2823), .A2(n_8_0_2734), .A3(n_8_0_7016), 
      .ZN(n_8_0_963));
   NAND3_X1 i_8_0_964 (.A1(n_8_0_2823), .A2(n_8_0_7013), .A3(n_8_0_7016), 
      .ZN(n_8_0_964));
   NAND3_X1 i_8_0_965 (.A1(n_8_0_2829), .A2(n_8_0_6861), .A3(n_8_0_7064), 
      .ZN(n_8_0_965));
   OR2_X1 i_8_0_966 (.A1(n_8_0_1244), .A2(\out_as[0] [4]), .ZN(n_8_0_966));
   OR2_X1 i_8_0_967 (.A1(n_8_0_1251), .A2(\out_as[0] [4]), .ZN(n_8_0_967));
   OR2_X1 i_8_0_968 (.A1(n_8_0_1297), .A2(n_8_0_556), .ZN(n_8_0_968));
   NAND2_X1 i_8_0_969 (.A1(n_8_0_1417), .A2(n_8_0_7027), .ZN(n_8_0_969));
   NAND2_X1 i_8_0_970 (.A1(n_8_0_2747), .A2(n_8_0_7038), .ZN(n_8_0_970));
   NAND2_X1 i_8_0_971 (.A1(n_8_0_2803), .A2(n_8_0_7050), .ZN(n_8_0_971));
   NAND2_X1 i_8_0_972 (.A1(n_8_0_2779), .A2(n_8_0_7038), .ZN(n_8_0_972));
   NAND2_X1 i_8_0_973 (.A1(n_8_0_2731), .A2(n_8_0_7086), .ZN(n_8_0_973));
   NAND2_X1 i_8_0_974 (.A1(n_8_0_2725), .A2(n_8_0_7062), .ZN(n_8_0_974));
   NAND2_X1 i_8_0_975 (.A1(n_8_0_2734), .A2(n_8_0_7014), .ZN(n_8_0_975));
   OR2_X1 i_8_0_976 (.A1(\out_as[7] [5]), .A2(n_8_0_657), .ZN(n_8_0_976));
   OR2_X1 i_8_0_977 (.A1(\out_as[7] [5]), .A2(n_8_0_704), .ZN(n_8_0_977));
   OR2_X1 i_8_0_978 (.A1(\out_as[7] [5]), .A2(n_8_0_736), .ZN(n_8_0_978));
   OR2_X1 i_8_0_979 (.A1(\out_as[7] [5]), .A2(n_8_0_752), .ZN(n_8_0_979));
   OR2_X1 i_8_0_980 (.A1(\out_as[7] [5]), .A2(n_8_0_768), .ZN(n_8_0_980));
   OR2_X1 i_8_0_981 (.A1(\out_as[7] [5]), .A2(n_8_0_784), .ZN(n_8_0_981));
   OR2_X1 i_8_0_982 (.A1(n_8_0_1360), .A2(n_8_0_506), .ZN(n_8_0_982));
   OR2_X1 i_8_0_983 (.A1(n_8_0_1360), .A2(n_8_0_545), .ZN(n_8_0_983));
   OR2_X1 i_8_0_984 (.A1(n_8_0_1336), .A2(\out_as[7] [5]), .ZN(n_8_0_984));
   OR2_X1 i_8_0_985 (.A1(n_8_0_1360), .A2(n_8_0_608), .ZN(n_8_0_985));
   OR2_X1 i_8_0_986 (.A1(n_8_0_1360), .A2(n_8_0_632), .ZN(n_8_0_986));
   OR2_X1 i_8_0_987 (.A1(n_8_0_1360), .A2(n_8_0_656), .ZN(n_8_0_987));
   OR2_X1 i_8_0_988 (.A1(n_8_0_1360), .A2(n_8_0_680), .ZN(n_8_0_988));
   OR2_X1 i_8_0_989 (.A1(n_8_0_1360), .A2(n_8_0_1286), .ZN(n_8_0_989));
   OR2_X1 i_8_0_990 (.A1(n_8_0_1360), .A2(n_8_0_1262), .ZN(n_8_0_990));
   OR2_X1 i_8_0_991 (.A1(n_8_0_1296), .A2(n_8_0_544), .ZN(n_8_0_991));
   OR2_X1 i_8_0_992 (.A1(n_8_0_1360), .A2(n_8_0_1240), .ZN(n_8_0_992));
   NAND2_X1 i_8_0_993 (.A1(n_8_0_1416), .A2(n_8_0_7002), .ZN(n_8_0_993));
   NAND2_X1 i_8_0_994 (.A1(n_8_0_2796), .A2(n_8_0_1416), .ZN(n_8_0_994));
   NAND2_X1 i_8_0_995 (.A1(n_8_0_2983), .A2(n_8_0_2796), .ZN(n_8_0_995));
   NAND2_X1 i_8_0_996 (.A1(n_8_0_2757), .A2(n_8_0_1416), .ZN(n_8_0_996));
   NAND2_X1 i_8_0_997 (.A1(n_8_0_2983), .A2(n_8_0_2757), .ZN(n_8_0_997));
   NAND2_X1 i_8_0_998 (.A1(n_8_0_2736), .A2(n_8_0_1416), .ZN(n_8_0_998));
   INV_X1 i_8_0_999 (.A(n_8_0_1416), .ZN(n_8_0_999));
   NOR2_X1 i_8_0_1000 (.A1(n_8_0_1296), .A2(\out_as[7] [5]), .ZN(n_8_0_1416));
   NAND2_X1 i_8_0_1001 (.A1(n_8_0_2983), .A2(n_8_0_2736), .ZN(n_8_0_1000));
   NAND2_X1 i_8_0_1002 (.A1(n_8_0_2736), .A2(n_8_0_7003), .ZN(n_8_0_1001));
   OR2_X1 i_8_0_1003 (.A1(\out_as[6] [5]), .A2(n_8_0_612), .ZN(n_8_0_1002));
   OR2_X1 i_8_0_1004 (.A1(\out_as[6] [5]), .A2(n_8_0_706), .ZN(n_8_0_1003));
   OR2_X1 i_8_0_1005 (.A1(\out_as[6] [5]), .A2(n_8_0_738), .ZN(n_8_0_1004));
   OR2_X1 i_8_0_1006 (.A1(n_8_0_1358), .A2(n_8_0_511), .ZN(n_8_0_1005));
   OR2_X1 i_8_0_1007 (.A1(n_8_0_1358), .A2(n_8_0_549), .ZN(n_8_0_1006));
   OR2_X1 i_8_0_1008 (.A1(n_8_0_1358), .A2(n_8_0_581), .ZN(n_8_0_1007));
   OR2_X1 i_8_0_1009 (.A1(n_8_0_1358), .A2(n_8_0_635), .ZN(n_8_0_1008));
   NAND2_X1 i_8_0_1010 (.A1(n_8_0_3204), .A2(n_8_0_6855), .ZN(n_8_0_1009));
   NAND2_X1 i_8_0_1011 (.A1(n_8_0_7016), .A2(n_8_0_6855), .ZN(n_8_0_1010));
   OR2_X1 i_8_0_1012 (.A1(n_8_0_1358), .A2(n_8_0_683), .ZN(n_8_0_1011));
   OR2_X1 i_8_0_1013 (.A1(n_8_0_1271), .A2(n_8_0_1206), .ZN(n_8_0_1012));
   OR2_X1 i_8_0_1014 (.A1(n_8_0_1220), .A2(n_8_0_509), .ZN(n_8_0_1013));
   NAND3_X1 i_8_0_1015 (.A1(n_8_0_3204), .A2(n_8_0_2823), .A3(n_8_0_7013), 
      .ZN(n_8_0_1014));
   NAND3_X1 i_8_0_1016 (.A1(n_8_0_3204), .A2(n_8_0_2823), .A3(n_8_0_2734), 
      .ZN(n_8_0_1015));
   OR2_X1 i_8_0_1017 (.A1(\out_as[5] [5]), .A2(n_8_0_517), .ZN(n_8_0_1016));
   OR2_X1 i_8_0_1018 (.A1(\out_as[5] [5]), .A2(n_8_0_554), .ZN(n_8_0_1017));
   OR2_X1 i_8_0_1019 (.A1(\out_as[5] [5]), .A2(n_8_0_586), .ZN(n_8_0_1018));
   OR2_X1 i_8_0_1020 (.A1(\out_as[5] [5]), .A2(n_8_0_615), .ZN(n_8_0_1019));
   OR2_X1 i_8_0_1021 (.A1(\out_as[5] [5]), .A2(n_8_0_639), .ZN(n_8_0_1020));
   OR2_X1 i_8_0_1022 (.A1(\out_as[5] [5]), .A2(n_8_0_687), .ZN(n_8_0_1021));
   OR2_X1 i_8_0_1023 (.A1(\out_as[5] [5]), .A2(n_8_0_708), .ZN(n_8_0_1022));
   OR2_X1 i_8_0_1024 (.A1(\out_as[5] [5]), .A2(n_8_0_724), .ZN(n_8_0_1023));
   OR2_X1 i_8_0_1025 (.A1(\out_as[5] [5]), .A2(n_8_0_740), .ZN(n_8_0_1024));
   OR2_X1 i_8_0_1026 (.A1(\out_as[5] [5]), .A2(n_8_0_756), .ZN(n_8_0_1025));
   OR2_X1 i_8_0_1027 (.A1(\out_as[5] [5]), .A2(n_8_0_772), .ZN(n_8_0_1026));
   OR2_X1 i_8_0_1028 (.A1(\out_as[5] [5]), .A2(n_8_0_788), .ZN(n_8_0_1027));
   OR2_X1 i_8_0_1029 (.A1(\out_as[5] [5]), .A2(n_8_0_804), .ZN(n_8_0_1028));
   OR2_X1 i_8_0_1030 (.A1(\out_as[5] [5]), .A2(n_8_0_820), .ZN(n_8_0_1029));
   OR2_X1 i_8_0_1031 (.A1(n_8_0_1354), .A2(n_8_0_516), .ZN(n_8_0_1030));
   OR2_X1 i_8_0_1032 (.A1(n_8_0_1354), .A2(n_8_0_553), .ZN(n_8_0_1031));
   OR2_X1 i_8_0_1033 (.A1(\out_as[5] [4]), .A2(n_8_0_553), .ZN(n_8_0_1032));
   OR2_X1 i_8_0_1034 (.A1(n_8_0_1354), .A2(n_8_0_585), .ZN(n_8_0_1033));
   OR2_X1 i_8_0_1035 (.A1(\out_as[5] [4]), .A2(n_8_0_585), .ZN(n_8_0_1034));
   OR2_X1 i_8_0_1036 (.A1(n_8_0_1354), .A2(n_8_0_614), .ZN(n_8_0_1035));
   OR2_X1 i_8_0_1037 (.A1(\out_as[5] [4]), .A2(n_8_0_614), .ZN(n_8_0_1036));
   OR2_X1 i_8_0_1038 (.A1(n_8_0_1354), .A2(n_8_0_638), .ZN(n_8_0_1037));
   OR2_X1 i_8_0_1039 (.A1(\out_as[5] [4]), .A2(n_8_0_638), .ZN(n_8_0_1038));
   OR2_X1 i_8_0_1040 (.A1(n_8_0_1354), .A2(n_8_0_662), .ZN(n_8_0_1039));
   OR2_X1 i_8_0_1041 (.A1(n_8_0_1354), .A2(n_8_0_686), .ZN(n_8_0_1040));
   OR2_X1 i_8_0_1042 (.A1(n_8_0_1354), .A2(n_8_0_1258), .ZN(n_8_0_1041));
   NAND3_X1 i_8_0_1043 (.A1(n_8_0_2854), .A2(n_8_0_7028), .A3(n_8_0_7029), 
      .ZN(n_8_0_1042));
   NAND2_X1 i_8_0_1044 (.A1(n_8_0_2816), .A2(n_8_0_2791), .ZN(n_8_0_1043));
   NAND2_X1 i_8_0_1045 (.A1(n_8_0_2958), .A2(n_8_0_2791), .ZN(n_8_0_1044));
   NAND2_X1 i_8_0_1046 (.A1(n_8_0_2816), .A2(n_8_0_1417), .ZN(n_8_0_1045));
   NAND2_X1 i_8_0_1047 (.A1(n_8_0_2958), .A2(n_8_0_1417), .ZN(n_8_0_1046));
   INV_X1 i_8_0_1048 (.A(n_8_0_1417), .ZN(n_8_0_1047));
   NOR2_X1 i_8_0_1049 (.A1(n_8_0_1201), .A2(\out_as[5] [0]), .ZN(n_8_0_1417));
   OR2_X1 i_8_0_1050 (.A1(\out_as[5] [1]), .A2(\out_as[5] [0]), .ZN(n_8_0_1048));
   OR2_X1 i_8_0_1051 (.A1(\out_as[4] [5]), .A2(n_8_0_558), .ZN(n_8_0_1049));
   OR2_X1 i_8_0_1052 (.A1(\out_as[4] [5]), .A2(n_8_0_666), .ZN(n_8_0_1050));
   OR2_X1 i_8_0_1053 (.A1(\out_as[4] [5]), .A2(n_8_0_690), .ZN(n_8_0_1051));
   OR2_X1 i_8_0_1054 (.A1(\out_as[4] [5]), .A2(n_8_0_726), .ZN(n_8_0_1052));
   OR2_X1 i_8_0_1055 (.A1(\out_as[4] [5]), .A2(n_8_0_742), .ZN(n_8_0_1053));
   OR2_X1 i_8_0_1056 (.A1(\out_as[4] [5]), .A2(n_8_0_758), .ZN(n_8_0_1054));
   OR2_X1 i_8_0_1057 (.A1(\out_as[4] [5]), .A2(n_8_0_774), .ZN(n_8_0_1055));
   OR2_X1 i_8_0_1058 (.A1(\out_as[4] [5]), .A2(n_8_0_790), .ZN(n_8_0_1056));
   OR2_X1 i_8_0_1059 (.A1(\out_as[4] [5]), .A2(n_8_0_806), .ZN(n_8_0_1057));
   OR2_X1 i_8_0_1060 (.A1(n_8_0_1357), .A2(n_8_0_521), .ZN(n_8_0_1058));
   OR2_X1 i_8_0_1061 (.A1(n_8_0_1357), .A2(n_8_0_557), .ZN(n_8_0_1059));
   OR2_X1 i_8_0_1062 (.A1(n_8_0_1357), .A2(n_8_0_589), .ZN(n_8_0_1060));
   OR2_X1 i_8_0_1063 (.A1(n_8_0_1357), .A2(n_8_0_617), .ZN(n_8_0_1061));
   OR2_X1 i_8_0_1064 (.A1(n_8_0_1357), .A2(n_8_0_641), .ZN(n_8_0_1062));
   OR2_X1 i_8_0_1065 (.A1(n_8_0_1357), .A2(n_8_0_665), .ZN(n_8_0_1063));
   OR2_X1 i_8_0_1066 (.A1(n_8_0_1357), .A2(n_8_0_689), .ZN(n_8_0_1064));
   OR2_X1 i_8_0_1067 (.A1(n_8_0_1357), .A2(n_8_0_1269), .ZN(n_8_0_1065));
   OR2_X1 i_8_0_1068 (.A1(n_8_0_1357), .A2(n_8_0_1252), .ZN(n_8_0_1066));
   NAND2_X1 i_8_0_1069 (.A1(n_8_0_1418), .A2(n_8_0_7037), .ZN(n_8_0_1067));
   NAND2_X1 i_8_0_1070 (.A1(n_8_0_2779), .A2(n_8_0_1418), .ZN(n_8_0_1068));
   NAND2_X1 i_8_0_1071 (.A1(n_8_0_2988), .A2(n_8_0_2779), .ZN(n_8_0_1069));
   NAND2_X1 i_8_0_1072 (.A1(n_8_0_2747), .A2(n_8_0_1418), .ZN(n_8_0_1070));
   NAND2_X1 i_8_0_1073 (.A1(n_8_0_2988), .A2(n_8_0_2747), .ZN(n_8_0_1071));
   NAND2_X1 i_8_0_1074 (.A1(n_8_0_2730), .A2(n_8_0_1418), .ZN(n_8_0_1072));
   NAND2_X1 i_8_0_1075 (.A1(n_8_0_2988), .A2(n_8_0_2730), .ZN(n_8_0_1073));
   INV_X1 i_8_0_1076 (.A(n_8_0_1418), .ZN(n_8_0_1074));
   NOR2_X1 i_8_0_1077 (.A1(n_8_0_1297), .A2(\out_as[4] [5]), .ZN(n_8_0_1418));
   OR2_X1 i_8_0_1078 (.A1(\out_as[3] [5]), .A2(n_8_0_527), .ZN(n_8_0_1075));
   OR2_X1 i_8_0_1079 (.A1(\out_as[3] [5]), .A2(n_8_0_645), .ZN(n_8_0_1076));
   OR2_X1 i_8_0_1080 (.A1(\out_as[3] [5]), .A2(n_8_0_669), .ZN(n_8_0_1077));
   OR2_X1 i_8_0_1081 (.A1(\out_as[3] [5]), .A2(n_8_0_693), .ZN(n_8_0_1078));
   OR2_X1 i_8_0_1082 (.A1(\out_as[3] [5]), .A2(n_8_0_728), .ZN(n_8_0_1079));
   OR2_X1 i_8_0_1083 (.A1(\out_as[3] [5]), .A2(n_8_0_744), .ZN(n_8_0_1080));
   OR2_X1 i_8_0_1084 (.A1(\out_as[3] [5]), .A2(n_8_0_760), .ZN(n_8_0_1081));
   OR2_X1 i_8_0_1085 (.A1(\out_as[3] [5]), .A2(n_8_0_776), .ZN(n_8_0_1082));
   OR2_X1 i_8_0_1086 (.A1(\out_as[3] [5]), .A2(n_8_0_792), .ZN(n_8_0_1083));
   OR2_X1 i_8_0_1087 (.A1(\out_as[3] [5]), .A2(n_8_0_808), .ZN(n_8_0_1084));
   OR2_X1 i_8_0_1088 (.A1(n_8_0_1353), .A2(n_8_0_526), .ZN(n_8_0_1085));
   OR2_X1 i_8_0_1089 (.A1(n_8_0_1353), .A2(n_8_0_561), .ZN(n_8_0_1086));
   OR2_X1 i_8_0_1090 (.A1(n_8_0_1353), .A2(n_8_0_593), .ZN(n_8_0_1087));
   OR2_X1 i_8_0_1091 (.A1(n_8_0_1353), .A2(n_8_0_620), .ZN(n_8_0_1088));
   OR2_X1 i_8_0_1092 (.A1(n_8_0_1353), .A2(n_8_0_644), .ZN(n_8_0_1089));
   OR2_X1 i_8_0_1093 (.A1(n_8_0_1353), .A2(n_8_0_668), .ZN(n_8_0_1090));
   OR2_X1 i_8_0_1094 (.A1(n_8_0_1353), .A2(n_8_0_1288), .ZN(n_8_0_1091));
   NAND2_X1 i_8_0_1095 (.A1(n_8_0_2893), .A2(n_8_0_7049), .ZN(n_8_0_1092));
   NAND2_X1 i_8_0_1096 (.A1(n_8_0_2893), .A2(n_8_0_2803), .ZN(n_8_0_1093));
   NAND2_X1 i_8_0_1097 (.A1(n_8_0_2963), .A2(n_8_0_2803), .ZN(n_8_0_1094));
   NAND2_X1 i_8_0_1098 (.A1(n_8_0_2893), .A2(n_8_0_2744), .ZN(n_8_0_1095));
   NAND2_X1 i_8_0_1099 (.A1(n_8_0_2963), .A2(n_8_0_2744), .ZN(n_8_0_1096));
   NAND2_X1 i_8_0_1100 (.A1(n_8_0_2893), .A2(n_8_0_2732), .ZN(n_8_0_1097));
   NAND2_X1 i_8_0_1101 (.A1(n_8_0_2963), .A2(n_8_0_2732), .ZN(n_8_0_1098));
   NAND2_X1 i_8_0_1102 (.A1(n_8_0_2963), .A2(n_8_0_7049), .ZN(n_8_0_1099));
   OR2_X1 i_8_0_1103 (.A1(\out_as[2] [5]), .A2(n_8_0_566), .ZN(n_8_0_1100));
   OR2_X1 i_8_0_1104 (.A1(\out_as[2] [5]), .A2(n_8_0_598), .ZN(n_8_0_1101));
   OR2_X1 i_8_0_1105 (.A1(\out_as[2] [5]), .A2(n_8_0_624), .ZN(n_8_0_1102));
   OR2_X1 i_8_0_1106 (.A1(\out_as[2] [5]), .A2(n_8_0_648), .ZN(n_8_0_1103));
   OR2_X1 i_8_0_1107 (.A1(\out_as[2] [5]), .A2(n_8_0_672), .ZN(n_8_0_1104));
   OR2_X1 i_8_0_1108 (.A1(\out_as[2] [5]), .A2(n_8_0_746), .ZN(n_8_0_1105));
   OR2_X1 i_8_0_1109 (.A1(\out_as[2] [5]), .A2(n_8_0_762), .ZN(n_8_0_1106));
   OR2_X1 i_8_0_1110 (.A1(\out_as[2] [5]), .A2(n_8_0_778), .ZN(n_8_0_1107));
   OR2_X1 i_8_0_1111 (.A1(n_8_0_1355), .A2(n_8_0_531), .ZN(n_8_0_1108));
   OR2_X1 i_8_0_1112 (.A1(n_8_0_1355), .A2(n_8_0_565), .ZN(n_8_0_1109));
   NAND2_X1 i_8_0_1113 (.A1(n_8_0_3191), .A2(n_8_0_6857), .ZN(n_8_0_1110));
   OR2_X1 i_8_0_1114 (.A1(n_8_0_1355), .A2(n_8_0_647), .ZN(n_8_0_1111));
   OR2_X1 i_8_0_1115 (.A1(n_8_0_1355), .A2(n_8_0_671), .ZN(n_8_0_1112));
   OR2_X1 i_8_0_1116 (.A1(n_8_0_1355), .A2(n_8_0_695), .ZN(n_8_0_1113));
   NAND2_X1 i_8_0_1117 (.A1(n_8_0_3191), .A2(n_8_0_2911), .ZN(n_8_0_1114));
   NAND2_X1 i_8_0_1118 (.A1(n_8_0_3191), .A2(n_8_0_2862), .ZN(n_8_0_1115));
   NAND2_X1 i_8_0_1119 (.A1(n_8_0_2862), .A2(n_8_0_7064), .ZN(n_8_0_1116));
   NAND3_X1 i_8_0_1120 (.A1(n_8_0_3191), .A2(n_8_0_2829), .A3(n_8_0_6861), 
      .ZN(n_8_0_1117));
   NAND2_X1 i_8_0_1121 (.A1(n_8_0_2829), .A2(n_8_0_6861), .ZN(n_8_0_1118));
   NAND2_X1 i_8_0_1122 (.A1(n_8_0_7062), .A2(n_8_0_6861), .ZN(n_8_0_1119));
   OR2_X1 i_8_0_1123 (.A1(n_8_0_1195), .A2(n_8_0_1121), .ZN(n_8_0_1120));
   NAND2_X1 i_8_0_1124 (.A1(n_8_0_3191), .A2(n_8_0_7063), .ZN(n_8_0_1121));
   NAND3_X1 i_8_0_1125 (.A1(n_8_0_2829), .A2(n_8_0_7061), .A3(n_8_0_7064), 
      .ZN(n_8_0_1122));
   NAND3_X1 i_8_0_1126 (.A1(n_8_0_3191), .A2(n_8_0_2829), .A3(n_8_0_2725), 
      .ZN(n_8_0_1123));
   NAND2_X1 i_8_0_1127 (.A1(n_8_0_7077), .A2(n_8_0_6860), .ZN(n_8_0_1124));
   OR2_X1 i_8_0_1128 (.A1(\out_as[1] [5]), .A2(n_8_0_651), .ZN(n_8_0_1125));
   OR2_X1 i_8_0_1129 (.A1(\out_as[1] [5]), .A2(n_8_0_675), .ZN(n_8_0_1126));
   OR2_X1 i_8_0_1130 (.A1(\out_as[1] [5]), .A2(n_8_0_716), .ZN(n_8_0_1127));
   OR2_X1 i_8_0_1131 (.A1(\out_as[1] [5]), .A2(n_8_0_764), .ZN(n_8_0_1128));
   OR2_X1 i_8_0_1132 (.A1(n_8_0_1356), .A2(n_8_0_536), .ZN(n_8_0_1129));
   OR2_X1 i_8_0_1133 (.A1(n_8_0_1356), .A2(n_8_0_569), .ZN(n_8_0_1130));
   OR2_X1 i_8_0_1134 (.A1(n_8_0_1356), .A2(n_8_0_601), .ZN(n_8_0_1131));
   OR2_X1 i_8_0_1135 (.A1(n_8_0_1356), .A2(n_8_0_626), .ZN(n_8_0_1132));
   OR2_X1 i_8_0_1136 (.A1(n_8_0_1356), .A2(n_8_0_650), .ZN(n_8_0_1133));
   OR2_X1 i_8_0_1137 (.A1(n_8_0_1356), .A2(n_8_0_674), .ZN(n_8_0_1134));
   OR2_X1 i_8_0_1138 (.A1(n_8_0_1356), .A2(n_8_0_698), .ZN(n_8_0_1135));
   OR2_X1 i_8_0_1139 (.A1(n_8_0_1356), .A2(n_8_0_1242), .ZN(n_8_0_1136));
   OR2_X1 i_8_0_1140 (.A1(n_8_0_1292), .A2(n_8_0_600), .ZN(n_8_0_1137));
   NAND2_X1 i_8_0_1141 (.A1(n_8_0_2841), .A2(n_8_0_2787), .ZN(n_8_0_1138));
   NAND2_X1 i_8_0_1142 (.A1(n_8_0_2970), .A2(n_8_0_2787), .ZN(n_8_0_1139));
   NAND2_X1 i_8_0_1143 (.A1(n_8_0_2970), .A2(n_8_0_7075), .ZN(n_8_0_1140));
   NAND2_X1 i_8_0_1144 (.A1(n_8_0_2841), .A2(n_8_0_2727), .ZN(n_8_0_1141));
   NAND2_X1 i_8_0_1145 (.A1(n_8_0_2841), .A2(n_8_0_2764), .ZN(n_8_0_1142));
   NAND2_X1 i_8_0_1146 (.A1(n_8_0_2970), .A2(n_8_0_2764), .ZN(n_8_0_1143));
   OR2_X1 i_8_0_1147 (.A1(\out_as[0] [5]), .A2(n_8_0_542), .ZN(n_8_0_1144));
   OR2_X1 i_8_0_1148 (.A1(\out_as[0] [5]), .A2(n_8_0_574), .ZN(n_8_0_1145));
   OR2_X1 i_8_0_1149 (.A1(\out_as[0] [5]), .A2(n_8_0_630), .ZN(n_8_0_1146));
   OR2_X1 i_8_0_1150 (.A1(\out_as[0] [5]), .A2(n_8_0_678), .ZN(n_8_0_1147));
   OR2_X1 i_8_0_1151 (.A1(\out_as[0] [5]), .A2(n_8_0_702), .ZN(n_8_0_1148));
   OR2_X1 i_8_0_1152 (.A1(\out_as[0] [5]), .A2(n_8_0_718), .ZN(n_8_0_1149));
   OR2_X1 i_8_0_1153 (.A1(\out_as[0] [5]), .A2(n_8_0_734), .ZN(n_8_0_1150));
   OR2_X1 i_8_0_1154 (.A1(\out_as[0] [5]), .A2(n_8_0_750), .ZN(n_8_0_1151));
   OR2_X1 i_8_0_1155 (.A1(\out_as[0] [5]), .A2(n_8_0_798), .ZN(n_8_0_1152));
   OR2_X1 i_8_0_1156 (.A1(\out_as[0] [5]), .A2(n_8_0_830), .ZN(n_8_0_1153));
   OR2_X1 i_8_0_1157 (.A1(n_8_0_1359), .A2(n_8_0_541), .ZN(n_8_0_1154));
   OR2_X1 i_8_0_1158 (.A1(n_8_0_1359), .A2(n_8_0_573), .ZN(n_8_0_1155));
   OR2_X1 i_8_0_1159 (.A1(n_8_0_1359), .A2(n_8_0_605), .ZN(n_8_0_1156));
   OR2_X1 i_8_0_1160 (.A1(n_8_0_1359), .A2(n_8_0_629), .ZN(n_8_0_1157));
   OR2_X1 i_8_0_1161 (.A1(n_8_0_1359), .A2(n_8_0_653), .ZN(n_8_0_1158));
   OR2_X1 i_8_0_1162 (.A1(n_8_0_1359), .A2(n_8_0_677), .ZN(n_8_0_1159));
   NAND2_X1 i_8_0_1163 (.A1(n_8_0_3208), .A2(n_8_0_2934), .ZN(n_8_0_1160));
   NAND2_X1 i_8_0_1164 (.A1(n_8_0_3208), .A2(n_8_0_2885), .ZN(n_8_0_1161));
   NAND2_X1 i_8_0_1165 (.A1(n_8_0_2977), .A2(n_8_0_2775), .ZN(n_8_0_1162));
   NAND2_X1 i_8_0_1166 (.A1(n_8_0_2775), .A2(n_8_0_7087), .ZN(n_8_0_1163));
   NAND2_X1 i_8_0_1167 (.A1(n_8_0_2977), .A2(n_8_0_2751), .ZN(n_8_0_1164));
   NAND3_X1 i_8_0_1168 (.A1(n_8_0_3208), .A2(n_8_0_2836), .A3(n_8_0_2731), 
      .ZN(n_8_0_1165));
   NAND2_X1 i_8_0_1169 (.A1(n_8_0_3208), .A2(n_8_0_2836), .ZN(n_8_0_1166));
   MUX2_X1 i_8_0_1170 (.A(n_8_0_1421), .B(n_8_0_1419), .S(n_8_0_2733), .Z(n_0));
   OAI21_X1 i_8_0_1171 (.A(n_8_0_1420), .B1(n_8_0_2735), .B2(n_8_0_6988), 
      .ZN(n_8_0_1419));
   NAND2_X1 i_8_0_1172 (.A1(in_data[4]), .A2(n_8_0_2735), .ZN(n_8_0_1420));
   MUX2_X1 i_8_0_1173 (.A(n_8_0_1422), .B(in_data[8]), .S(n_8_0_1423), .Z(
      n_8_0_1421));
   MUX2_X1 i_8_0_1174 (.A(n_8_0_1424), .B(in_data[12]), .S(n_8_0_1425), .Z(
      n_8_0_1422));
   OAI21_X1 i_8_0_1175 (.A(n_8_0_6824), .B1(n_8_0_2768), .B2(\out_as[5] [0]), 
      .ZN(n_8_0_1423));
   MUX2_X1 i_8_0_1176 (.A(in_data[16]), .B(n_8_0_1426), .S(n_8_0_1427), .Z(
      n_8_0_1424));
   NAND2_X1 i_8_0_1177 (.A1(n_8_0_6795), .A2(n_8_0_2729), .ZN(n_8_0_1425));
   MUX2_X1 i_8_0_1178 (.A(n_8_0_1428), .B(in_data[20]), .S(n_8_0_1429), .Z(
      n_8_0_1426));
   AOI21_X1 i_8_0_1179 (.A(n_8_0_6838), .B1(n_8_0_2962), .B2(n_8_0_2732), 
      .ZN(n_8_0_1427));
   MUX2_X1 i_8_0_1180 (.A(in_data[24]), .B(in_data[28]), .S(n_8_0_1430), 
      .Z(n_8_0_1428));
   NAND2_X1 i_8_0_1181 (.A1(n_8_0_6772), .A2(n_8_0_2724), .ZN(n_8_0_1429));
   NOR2_X1 i_8_0_1182 (.A1(n_8_0_6781), .A2(n_8_0_2726), .ZN(n_8_0_1430));
   AOI21_X1 i_8_0_1183 (.A(n_8_0_1431), .B1(n_8_0_2753), .B2(n_8_0_6988), 
      .ZN(n_1));
   NOR2_X1 i_8_0_1184 (.A1(n_8_0_2753), .A2(n_8_0_1432), .ZN(n_8_0_1431));
   AOI21_X1 i_8_0_1185 (.A(n_8_0_1433), .B1(n_8_0_1434), .B2(n_8_0_2738), 
      .ZN(n_8_0_1432));
   NOR2_X1 i_8_0_1186 (.A1(n_8_0_2738), .A2(in_data[4]), .ZN(n_8_0_1433));
   OAI21_X1 i_8_0_1187 (.A(n_8_0_1435), .B1(n_8_0_1436), .B2(n_8_0_2765), 
      .ZN(n_8_0_1434));
   NAND2_X1 i_8_0_1188 (.A1(n_8_0_2765), .A2(n_8_0_6990), .ZN(n_8_0_1435));
   MUX2_X1 i_8_0_1189 (.A(in_data[12]), .B(n_8_0_1437), .S(n_8_0_2745), .Z(
      n_8_0_1436));
   OAI21_X1 i_8_0_1190 (.A(n_8_0_1438), .B1(n_8_0_2741), .B2(n_8_0_6992), 
      .ZN(n_8_0_1437));
   OAI211_X1 i_8_0_1191 (.A(n_8_0_2741), .B(n_8_0_1439), .C1(n_8_0_1440), 
      .C2(n_8_0_2758), .ZN(n_8_0_1438));
   NAND2_X1 i_8_0_1192 (.A1(n_8_0_6993), .A2(n_8_0_2758), .ZN(n_8_0_1439));
   MUX2_X1 i_8_0_1193 (.A(in_data[28]), .B(in_data[24]), .S(n_8_0_2761), 
      .Z(n_8_0_1440));
   MUX2_X1 i_8_0_1194 (.A(in_data[0]), .B(n_8_0_1441), .S(n_8_0_1448), .Z(n_2));
   AOI22_X1 i_8_0_1195 (.A1(n_8_0_1442), .A2(n_8_0_1443), .B1(n_8_0_2781), 
      .B2(n_8_0_6989), .ZN(n_8_0_1441));
   AOI21_X1 i_8_0_1196 (.A(n_8_0_2781), .B1(n_8_0_2789), .B2(in_data[8]), 
      .ZN(n_8_0_1442));
   OAI211_X1 i_8_0_1197 (.A(n_8_0_1444), .B(n_8_0_2788), .C1(in_data[12]), 
      .C2(n_8_0_2777), .ZN(n_8_0_1443));
   OAI211_X1 i_8_0_1198 (.A(n_8_0_2777), .B(n_8_0_1445), .C1(n_8_0_6992), 
      .C2(n_8_0_2801), .ZN(n_8_0_1444));
   OAI211_X1 i_8_0_1199 (.A(n_8_0_2801), .B(n_8_0_1446), .C1(n_8_0_1447), 
      .C2(n_8_0_2798), .ZN(n_8_0_1445));
   NAND2_X1 i_8_0_1200 (.A1(n_8_0_2798), .A2(n_8_0_6993), .ZN(n_8_0_1446));
   MUX2_X1 i_8_0_1201 (.A(in_data[28]), .B(in_data[24]), .S(n_8_0_2784), 
      .Z(n_8_0_1447));
   AOI21_X1 i_8_0_1202 (.A(n_8_0_2792), .B1(n_8_0_2794), .B2(n_8_0_6729), 
      .ZN(n_8_0_1448));
   OAI21_X1 i_8_0_1203 (.A(n_8_0_1449), .B1(n_8_0_2830), .B2(n_8_0_6988), 
      .ZN(n_3));
   OAI221_X1 i_8_0_1204 (.A(n_8_0_2830), .B1(n_8_0_2819), .B2(in_data[4]), 
      .C1(n_8_0_1450), .C2(n_8_0_1451), .ZN(n_8_0_1449));
   OAI21_X1 i_8_0_1205 (.A(n_8_0_2819), .B1(n_8_0_2812), .B2(n_8_0_1452), 
      .ZN(n_8_0_1450));
   AND2_X1 i_8_0_1206 (.A1(in_data[8]), .A2(n_8_0_2812), .ZN(n_8_0_1451));
   AOI21_X1 i_8_0_1207 (.A(n_8_0_1453), .B1(n_8_0_1454), .B2(n_8_0_2843), 
      .ZN(n_8_0_1452));
   NOR2_X1 i_8_0_1208 (.A1(n_8_0_6991), .A2(n_8_0_2843), .ZN(n_8_0_1453));
   AOI21_X1 i_8_0_1209 (.A(n_8_0_1455), .B1(n_8_0_2809), .B2(n_8_0_6992), 
      .ZN(n_8_0_1454));
   NOR2_X1 i_8_0_1210 (.A1(n_8_0_2809), .A2(n_8_0_1456), .ZN(n_8_0_1455));
   MUX2_X1 i_8_0_1211 (.A(n_8_0_1457), .B(in_data[20]), .S(n_8_0_2824), .Z(
      n_8_0_1456));
   MUX2_X1 i_8_0_1212 (.A(in_data[28]), .B(in_data[24]), .S(n_8_0_2837), 
      .Z(n_8_0_1457));
   MUX2_X1 i_8_0_1213 (.A(n_8_0_1458), .B(in_data[0]), .S(n_8_0_2855), .Z(n_4));
   OAI21_X1 i_8_0_1214 (.A(n_8_0_1459), .B1(n_8_0_2871), .B2(n_8_0_6989), 
      .ZN(n_8_0_1458));
   OAI211_X1 i_8_0_1215 (.A(n_8_0_2871), .B(n_8_0_1460), .C1(n_8_0_1461), 
      .C2(n_8_0_2852), .ZN(n_8_0_1459));
   NAND2_X1 i_8_0_1216 (.A1(n_8_0_6990), .A2(n_8_0_2852), .ZN(n_8_0_1460));
   OAI22_X1 i_8_0_1217 (.A1(n_8_0_1463), .A2(n_8_0_1462), .B1(n_8_0_6991), 
      .B2(n_8_0_2847), .ZN(n_8_0_1461));
   OAI21_X1 i_8_0_1218 (.A(n_8_0_2847), .B1(n_8_0_2874), .B2(in_data[16]), 
      .ZN(n_8_0_1462));
   AOI211_X1 i_8_0_1219 (.A(n_8_0_2875), .B(n_8_0_1464), .C1(n_8_0_1465), 
      .C2(n_8_0_2860), .ZN(n_8_0_1463));
   NOR2_X1 i_8_0_1220 (.A1(n_8_0_2860), .A2(n_8_0_6993), .ZN(n_8_0_1464));
   MUX2_X1 i_8_0_1221 (.A(in_data[24]), .B(in_data[28]), .S(n_8_0_2864), 
      .Z(n_8_0_1465));
   AOI22_X1 i_8_0_1222 (.A1(n_8_0_1467), .A2(n_8_0_1466), .B1(n_8_0_6988), 
      .B2(n_8_0_2906), .ZN(n_5));
   AOI21_X1 i_8_0_1223 (.A(n_8_0_2906), .B1(n_8_0_2901), .B2(in_data[4]), 
      .ZN(n_8_0_1466));
   OAI211_X1 i_8_0_1224 (.A(n_8_0_2900), .B(n_8_0_1468), .C1(n_8_0_1469), 
      .C2(n_8_0_2896), .ZN(n_8_0_1467));
   NAND2_X1 i_8_0_1225 (.A1(n_8_0_6990), .A2(n_8_0_2896), .ZN(n_8_0_1468));
   MUX2_X1 i_8_0_1226 (.A(in_data[12]), .B(n_8_0_1470), .S(n_8_0_2886), .Z(
      n_8_0_1469));
   AOI21_X1 i_8_0_1227 (.A(n_8_0_1471), .B1(n_8_0_2890), .B2(n_8_0_6992), 
      .ZN(n_8_0_1470));
   AOI211_X1 i_8_0_1228 (.A(n_8_0_2890), .B(n_8_0_1472), .C1(in_data[20]), 
      .C2(n_8_0_2909), .ZN(n_8_0_1471));
   AOI211_X1 i_8_0_1229 (.A(n_8_0_1473), .B(n_8_0_2909), .C1(n_8_0_2913), 
      .C2(n_8_0_6995), .ZN(n_8_0_1472));
   NOR2_X1 i_8_0_1230 (.A1(in_data[24]), .A2(n_8_0_2913), .ZN(n_8_0_1473));
   OAI22_X1 i_8_0_1231 (.A1(n_8_0_1475), .A2(n_8_0_1474), .B1(n_8_0_6988), 
      .B2(n_8_0_2943), .ZN(n_6));
   OAI21_X1 i_8_0_1232 (.A(n_8_0_2943), .B1(n_8_0_2924), .B2(in_data[4]), 
      .ZN(n_8_0_1474));
   AOI21_X1 i_8_0_1233 (.A(n_8_0_1476), .B1(n_8_0_1477), .B2(n_8_0_2928), 
      .ZN(n_8_0_1475));
   OAI21_X1 i_8_0_1234 (.A(n_8_0_2924), .B1(n_8_0_2928), .B2(n_8_0_6990), 
      .ZN(n_8_0_1476));
   AOI21_X1 i_8_0_1235 (.A(n_8_0_1478), .B1(n_8_0_1479), .B2(n_8_0_2921), 
      .ZN(n_8_0_1477));
   NOR2_X1 i_8_0_1236 (.A1(n_8_0_2921), .A2(in_data[12]), .ZN(n_8_0_1478));
   OAI21_X1 i_8_0_1237 (.A(n_8_0_1480), .B1(n_8_0_2947), .B2(in_data[16]), 
      .ZN(n_8_0_1479));
   NAND2_X1 i_8_0_1238 (.A1(n_8_0_2947), .A2(n_8_0_1481), .ZN(n_8_0_1480));
   OAI21_X1 i_8_0_1239 (.A(n_8_0_1483), .B1(n_8_0_1482), .B2(n_8_0_2939), 
      .ZN(n_8_0_1481));
   MUX2_X1 i_8_0_1240 (.A(in_data[24]), .B(in_data[28]), .S(n_8_0_2935), 
      .Z(n_8_0_1482));
   NAND2_X1 i_8_0_1241 (.A1(n_8_0_2939), .A2(n_8_0_6993), .ZN(n_8_0_1483));
   OAI21_X1 i_8_0_1244 (.A(n_8_0_2964), .B1(n_8_0_1487), .B2(n_8_0_1486), 
      .ZN(n_8_0_1485));
   NOR2_X1 i_8_0_1245 (.A1(n_8_0_6990), .A2(n_8_0_2955), .ZN(n_8_0_1486));
   AOI21_X1 i_8_0_1246 (.A(n_8_0_1488), .B1(n_8_0_1489), .B2(n_8_0_2984), 
      .ZN(n_8_0_1487));
   OAI21_X1 i_8_0_1247 (.A(n_8_0_2955), .B1(n_8_0_2984), .B2(in_data[12]), 
      .ZN(n_8_0_1488));
   INV_X1 i_8_0_1248 (.A(n_8_0_1490), .ZN(n_8_0_1489));
   NOR2_X1 i_8_0_1249 (.A1(n_8_0_1492), .A2(n_8_0_1491), .ZN(n_8_0_1490));
   NOR2_X1 i_8_0_1250 (.A1(in_data[16]), .A2(n_8_0_2959), .ZN(n_8_0_1491));
   AOI21_X1 i_8_0_1251 (.A(n_8_0_1493), .B1(n_8_0_1494), .B2(n_8_0_2972), 
      .ZN(n_8_0_1492));
   OAI21_X1 i_8_0_1252 (.A(n_8_0_2959), .B1(n_8_0_2972), .B2(n_8_0_6993), 
      .ZN(n_8_0_1493));
   AOI21_X1 i_8_0_1253 (.A(n_8_0_1495), .B1(n_8_0_2967), .B2(n_8_0_6995), 
      .ZN(n_8_0_1494));
   NOR2_X1 i_8_0_1254 (.A1(in_data[24]), .A2(n_8_0_2967), .ZN(n_8_0_1495));
   AOI21_X1 i_8_0_1255 (.A(n_8_0_1496), .B1(n_8_0_3007), .B2(n_8_0_6988), 
      .ZN(n_7));
   AOI21_X1 i_8_0_1256 (.A(n_8_0_1497), .B1(n_8_0_1498), .B2(n_8_0_3004), 
      .ZN(n_8_0_1496));
   OAI21_X1 i_8_0_1257 (.A(n_8_0_3008), .B1(n_8_0_3004), .B2(n_8_0_6989), 
      .ZN(n_8_0_1497));
   MUX2_X1 i_8_0_1258 (.A(n_8_0_1499), .B(in_data[8]), .S(n_8_0_2992), .Z(
      n_8_0_1498));
   OAI21_X1 i_8_0_1259 (.A(n_8_0_1500), .B1(n_8_0_1501), .B2(n_8_0_2994), 
      .ZN(n_8_0_1499));
   NAND2_X1 i_8_0_1260 (.A1(in_data[12]), .A2(n_8_0_2994), .ZN(n_8_0_1500));
   AOI21_X1 i_8_0_1261 (.A(n_8_0_1502), .B1(n_8_0_1503), .B2(n_8_0_2998), 
      .ZN(n_8_0_1501));
   NOR2_X1 i_8_0_1262 (.A1(n_8_0_2998), .A2(n_8_0_6992), .ZN(n_8_0_1502));
   OAI21_X1 i_8_0_1263 (.A(n_8_0_1504), .B1(n_8_0_3017), .B2(n_8_0_6993), 
      .ZN(n_8_0_1503));
   NAND2_X1 i_8_0_1264 (.A1(n_8_0_3017), .A2(n_8_0_1505), .ZN(n_8_0_1504));
   MUX2_X1 i_8_0_1265 (.A(in_data[24]), .B(in_data[28]), .S(n_8_0_3011), 
      .Z(n_8_0_1505));
   OAI22_X1 i_8_0_1266 (.A1(n_8_0_1507), .A2(n_8_0_1506), .B1(n_8_0_6988), 
      .B2(n_8_0_3035), .ZN(n_8));
   OAI21_X1 i_8_0_1267 (.A(n_8_0_3035), .B1(n_8_0_3045), .B2(in_data[4]), 
      .ZN(n_8_0_1506));
   NOR2_X1 i_8_0_1268 (.A1(n_8_0_1509), .A2(n_8_0_1508), .ZN(n_8_0_1507));
   OAI21_X1 i_8_0_1269 (.A(n_8_0_3045), .B1(n_8_0_3031), .B2(n_8_0_6990), 
      .ZN(n_8_0_1508));
   AOI21_X1 i_8_0_1270 (.A(n_8_0_1510), .B1(n_8_0_1511), .B2(n_8_0_3029), 
      .ZN(n_8_0_1509));
   OAI21_X1 i_8_0_1271 (.A(n_8_0_3031), .B1(n_8_0_3029), .B2(in_data[12]), 
      .ZN(n_8_0_1510));
   OAI21_X1 i_8_0_1272 (.A(n_8_0_1512), .B1(n_8_0_3026), .B2(in_data[16]), 
      .ZN(n_8_0_1511));
   OAI211_X1 i_8_0_1273 (.A(n_8_0_1513), .B(n_8_0_3026), .C1(n_8_0_3038), 
      .C2(n_8_0_6993), .ZN(n_8_0_1512));
   NAND2_X1 i_8_0_1274 (.A1(n_8_0_3038), .A2(n_8_0_1514), .ZN(n_8_0_1513));
   MUX2_X1 i_8_0_1275 (.A(in_data[24]), .B(in_data[28]), .S(n_8_0_3042), 
      .Z(n_8_0_1514));
   OAI21_X1 i_8_0_1276 (.A(n_8_0_1515), .B1(n_8_0_1517), .B2(n_8_0_6988), 
      .ZN(n_9));
   OAI21_X1 i_8_0_1277 (.A(n_8_0_1517), .B1(n_8_0_1516), .B2(n_8_0_1518), 
      .ZN(n_8_0_1515));
   AND2_X1 i_8_0_1278 (.A1(n_8_0_3058), .A2(in_data[4]), .ZN(n_8_0_1516));
   AOI21_X1 i_8_0_1279 (.A(n_8_0_3052), .B1(n_8_0_3051), .B2(n_8_0_6729), 
      .ZN(n_8_0_1517));
   AOI211_X1 i_8_0_1280 (.A(n_8_0_3058), .B(n_8_0_1519), .C1(n_8_0_1520), 
      .C2(n_8_0_3072), .ZN(n_8_0_1518));
   NOR2_X1 i_8_0_1281 (.A1(n_8_0_3072), .A2(in_data[8]), .ZN(n_8_0_1519));
   OAI21_X1 i_8_0_1282 (.A(n_8_0_1523), .B1(n_8_0_1521), .B2(n_8_0_3061), 
      .ZN(n_8_0_1520));
   OAI21_X1 i_8_0_1283 (.A(n_8_0_1522), .B1(n_8_0_3054), .B2(n_8_0_6995), 
      .ZN(n_8_0_1521));
   NAND2_X1 i_8_0_1284 (.A1(n_8_0_3054), .A2(in_data[24]), .ZN(n_8_0_1522));
   OAI21_X1 i_8_0_1285 (.A(n_8_0_1524), .B1(n_8_0_3062), .B2(n_8_0_6991), 
      .ZN(n_8_0_1523));
   NAND2_X1 i_8_0_1286 (.A1(n_8_0_1525), .A2(n_8_0_3062), .ZN(n_8_0_1524));
   OAI21_X1 i_8_0_1287 (.A(n_8_0_1526), .B1(n_8_0_3069), .B2(n_8_0_6992), 
      .ZN(n_8_0_1525));
   OAI21_X1 i_8_0_1288 (.A(n_8_0_3069), .B1(n_8_0_3066), .B2(in_data[20]), 
      .ZN(n_8_0_1526));
   NAND2_X1 i_8_0_1293 (.A1(n_8_0_1531), .A2(n_8_0_3087), .ZN(n_8_0_1530));
   OAI21_X1 i_8_0_1294 (.A(n_8_0_1532), .B1(n_8_0_3093), .B2(n_8_0_6991), 
      .ZN(n_8_0_1531));
   OAI211_X1 i_8_0_1295 (.A(n_8_0_3093), .B(n_8_0_1533), .C1(n_8_0_1534), 
      .C2(n_8_0_3095), .ZN(n_8_0_1532));
   NAND2_X1 i_8_0_1296 (.A1(n_8_0_6992), .A2(n_8_0_3095), .ZN(n_8_0_1533));
   AOI21_X1 i_8_0_1297 (.A(n_8_0_1535), .B1(n_8_0_3085), .B2(n_8_0_6993), 
      .ZN(n_8_0_1534));
   AOI211_X1 i_8_0_1298 (.A(n_8_0_3085), .B(n_8_0_1536), .C1(n_8_0_3082), 
      .C2(in_data[24]), .ZN(n_8_0_1535));
   NOR2_X1 i_8_0_1299 (.A1(n_8_0_6995), .A2(n_8_0_3082), .ZN(n_8_0_1536));
   AOI21_X1 i_8_0_1300 (.A(n_8_0_1537), .B1(n_8_0_3114), .B2(n_8_0_6988), 
      .ZN(n_10));
   NOR2_X1 i_8_0_1301 (.A1(n_8_0_3114), .A2(n_8_0_1538), .ZN(n_8_0_1537));
   AOI22_X1 i_8_0_1302 (.A1(n_8_0_1540), .A2(n_8_0_1539), .B1(n_8_0_6989), 
      .B2(n_8_0_3102), .ZN(n_8_0_1538));
   AOI21_X1 i_8_0_1303 (.A(n_8_0_3102), .B1(n_8_0_3120), .B2(in_data[8]), 
      .ZN(n_8_0_1539));
   OAI221_X1 i_8_0_1304 (.A(n_8_0_3121), .B1(n_8_0_3105), .B2(in_data[12]), 
      .C1(n_8_0_1542), .C2(n_8_0_1541), .ZN(n_8_0_1540));
   OAI21_X1 i_8_0_1305 (.A(n_8_0_3105), .B1(n_8_0_3118), .B2(n_8_0_6992), 
      .ZN(n_8_0_1541));
   AND2_X1 i_8_0_1306 (.A1(n_8_0_3118), .A2(n_8_0_1543), .ZN(n_8_0_1542));
   AOI21_X1 i_8_0_1307 (.A(n_8_0_1544), .B1(n_8_0_1545), .B2(n_8_0_3111), 
      .ZN(n_8_0_1543));
   NOR2_X1 i_8_0_1308 (.A1(n_8_0_3111), .A2(in_data[20]), .ZN(n_8_0_1544));
   OAI21_X1 i_8_0_1309 (.A(n_8_0_1546), .B1(n_8_0_3108), .B2(in_data[24]), 
      .ZN(n_8_0_1545));
   NAND2_X1 i_8_0_1310 (.A1(n_8_0_3108), .A2(n_8_0_6995), .ZN(n_8_0_1546));
   MUX2_X1 i_8_0_1311 (.A(n_8_0_1547), .B(in_data[0]), .S(n_8_0_3139), .Z(n_11));
   MUX2_X1 i_8_0_1312 (.A(in_data[4]), .B(n_8_0_1548), .S(n_8_0_3131), .Z(
      n_8_0_1547));
   OAI22_X1 i_8_0_1313 (.A1(n_8_0_1550), .A2(n_8_0_1549), .B1(n_8_0_6990), 
      .B2(n_8_0_3145), .ZN(n_8_0_1548));
   OAI21_X1 i_8_0_1314 (.A(n_8_0_3145), .B1(n_8_0_3129), .B2(in_data[12]), 
      .ZN(n_8_0_1549));
   AOI21_X1 i_8_0_1315 (.A(n_8_0_1551), .B1(n_8_0_3142), .B2(in_data[16]), 
      .ZN(n_8_0_1550));
   OAI21_X1 i_8_0_1316 (.A(n_8_0_3129), .B1(n_8_0_1552), .B2(n_8_0_3142), 
      .ZN(n_8_0_1551));
   OAI22_X1 i_8_0_1317 (.A1(n_8_0_1553), .A2(n_8_0_1554), .B1(n_8_0_3137), 
      .B2(in_data[20]), .ZN(n_8_0_1552));
   OAI21_X1 i_8_0_1318 (.A(n_8_0_3137), .B1(n_8_0_3134), .B2(n_8_0_6995), 
      .ZN(n_8_0_1553));
   AND2_X1 i_8_0_1319 (.A1(n_8_0_3134), .A2(in_data[24]), .ZN(n_8_0_1554));
   OAI22_X1 i_8_0_1320 (.A1(n_8_0_1556), .A2(n_8_0_1555), .B1(n_8_0_6988), 
      .B2(n_8_0_3171), .ZN(n_12));
   OAI21_X1 i_8_0_1321 (.A(n_8_0_3171), .B1(n_8_0_3163), .B2(in_data[4]), 
      .ZN(n_8_0_1555));
   AOI211_X1 i_8_0_1322 (.A(n_8_0_3162), .B(n_8_0_1557), .C1(n_8_0_3153), 
      .C2(in_data[8]), .ZN(n_8_0_1556));
   AOI211_X1 i_8_0_1323 (.A(n_8_0_3153), .B(n_8_0_1558), .C1(n_8_0_6991), 
      .C2(n_8_0_3155), .ZN(n_8_0_1557));
   AOI211_X1 i_8_0_1324 (.A(n_8_0_3155), .B(n_8_0_1559), .C1(in_data[16]), 
      .C2(n_8_0_3159), .ZN(n_8_0_1558));
   AOI211_X1 i_8_0_1325 (.A(n_8_0_3159), .B(n_8_0_1560), .C1(n_8_0_1561), 
      .C2(n_8_0_3165), .ZN(n_8_0_1559));
   NOR2_X1 i_8_0_1326 (.A1(n_8_0_3165), .A2(in_data[20]), .ZN(n_8_0_1560));
   AOI21_X1 i_8_0_1327 (.A(n_8_0_1562), .B1(n_8_0_3168), .B2(in_data[24]), 
      .ZN(n_8_0_1561));
   NOR2_X1 i_8_0_1328 (.A1(n_8_0_3168), .A2(n_8_0_6995), .ZN(n_8_0_1562));
   OAI21_X1 i_8_0_1329 (.A(n_8_0_1563), .B1(n_8_0_3209), .B2(n_8_0_6988), 
      .ZN(n_13));
   NAND2_X1 i_8_0_1330 (.A1(n_8_0_3209), .A2(n_8_0_1564), .ZN(n_8_0_1563));
   MUX2_X1 i_8_0_1331 (.A(in_data[4]), .B(n_8_0_1565), .S(n_8_0_3200), .Z(
      n_8_0_1564));
   MUX2_X1 i_8_0_1332 (.A(in_data[8]), .B(n_8_0_1566), .S(n_8_0_3182), .Z(
      n_8_0_1565));
   MUX2_X1 i_8_0_1333 (.A(in_data[12]), .B(n_8_0_1567), .S(n_8_0_3196), .Z(
      n_8_0_1566));
   OAI21_X1 i_8_0_1334 (.A(n_8_0_1568), .B1(n_8_0_3177), .B2(n_8_0_6992), 
      .ZN(n_8_0_1567));
   NAND2_X1 i_8_0_1335 (.A1(n_8_0_3177), .A2(n_8_0_1569), .ZN(n_8_0_1568));
   MUX2_X1 i_8_0_1336 (.A(n_8_0_1570), .B(in_data[20]), .S(n_8_0_3187), .Z(
      n_8_0_1569));
   MUX2_X1 i_8_0_1337 (.A(in_data[24]), .B(in_data[28]), .S(n_8_0_3192), 
      .Z(n_8_0_1570));
   OAI21_X1 i_8_0_1338 (.A(n_8_0_1571), .B1(n_8_0_3241), .B2(n_8_0_6988), 
      .ZN(n_14));
   NAND2_X1 i_8_0_1339 (.A1(n_8_0_1572), .A2(n_8_0_3241), .ZN(n_8_0_1571));
   MUX2_X1 i_8_0_1340 (.A(n_8_0_1573), .B(in_data[4]), .S(n_8_0_3235), .Z(
      n_8_0_1572));
   MUX2_X1 i_8_0_1341 (.A(n_8_0_1574), .B(in_data[8]), .S(n_8_0_3224), .Z(
      n_8_0_1573));
   OAI22_X1 i_8_0_1342 (.A1(n_8_0_1576), .A2(n_8_0_1575), .B1(n_8_0_6991), 
      .B2(n_8_0_3219), .ZN(n_8_0_1574));
   OAI21_X1 i_8_0_1343 (.A(n_8_0_3219), .B1(n_8_0_3228), .B2(in_data[16]), 
      .ZN(n_8_0_1575));
   AOI21_X1 i_8_0_1344 (.A(n_8_0_1577), .B1(n_8_0_1578), .B2(n_8_0_3231), 
      .ZN(n_8_0_1576));
   OAI21_X1 i_8_0_1345 (.A(n_8_0_3228), .B1(n_8_0_3231), .B2(n_8_0_6993), 
      .ZN(n_8_0_1577));
   OAI21_X1 i_8_0_1346 (.A(n_8_0_1579), .B1(n_8_0_3216), .B2(n_8_0_6995), 
      .ZN(n_8_0_1578));
   NAND2_X1 i_8_0_1347 (.A1(n_8_0_3216), .A2(in_data[24]), .ZN(n_8_0_1579));
   OAI22_X1 i_8_0_1348 (.A1(n_8_0_1581), .A2(n_8_0_1580), .B1(n_8_0_6988), 
      .B2(n_8_0_3256), .ZN(n_15));
   OAI21_X1 i_8_0_1349 (.A(n_8_0_3256), .B1(n_8_0_3273), .B2(in_data[4]), 
      .ZN(n_8_0_1580));
   AOI211_X1 i_8_0_1350 (.A(n_8_0_3272), .B(n_8_0_1582), .C1(n_8_0_3266), 
      .C2(in_data[8]), .ZN(n_8_0_1581));
   AOI211_X1 i_8_0_1351 (.A(n_8_0_3266), .B(n_8_0_1583), .C1(n_8_0_1584), 
      .C2(n_8_0_3253), .ZN(n_8_0_1582));
   NOR2_X1 i_8_0_1352 (.A1(in_data[12]), .A2(n_8_0_3253), .ZN(n_8_0_1583));
   OAI21_X1 i_8_0_1353 (.A(n_8_0_1585), .B1(n_8_0_1586), .B2(n_8_0_3250), 
      .ZN(n_8_0_1584));
   NAND2_X1 i_8_0_1354 (.A1(n_8_0_6992), .A2(n_8_0_3250), .ZN(n_8_0_1585));
   AOI22_X1 i_8_0_1355 (.A1(n_8_0_1587), .A2(n_8_0_1588), .B1(n_8_0_3263), 
      .B2(n_8_0_6993), .ZN(n_8_0_1586));
   AOI21_X1 i_8_0_1356 (.A(n_8_0_3263), .B1(n_8_0_3260), .B2(in_data[28]), 
      .ZN(n_8_0_1587));
   NAND2_X1 i_8_0_1357 (.A1(n_8_0_3259), .A2(in_data[24]), .ZN(n_8_0_1588));
   AOI21_X1 i_8_0_1361 (.A(n_8_0_3285), .B1(n_8_0_3296), .B2(n_8_0_6990), 
      .ZN(n_8_0_1591));
   MUX2_X1 i_8_0_1362 (.A(in_data[12]), .B(n_8_0_1593), .S(n_8_0_3298), .Z(
      n_8_0_1592));
   AOI21_X1 i_8_0_1363 (.A(n_8_0_1594), .B1(n_8_0_3280), .B2(n_8_0_6992), 
      .ZN(n_8_0_1593));
   NOR2_X1 i_8_0_1364 (.A1(n_8_0_1595), .A2(n_8_0_3280), .ZN(n_8_0_1594));
   AOI21_X1 i_8_0_1365 (.A(n_8_0_1596), .B1(n_8_0_1597), .B2(n_8_0_3293), 
      .ZN(n_8_0_1595));
   NOR2_X1 i_8_0_1366 (.A1(n_8_0_3293), .A2(in_data[20]), .ZN(n_8_0_1596));
   OAI21_X1 i_8_0_1367 (.A(n_8_0_1598), .B1(n_8_0_3290), .B2(in_data[24]), 
      .ZN(n_8_0_1597));
   NAND2_X1 i_8_0_1368 (.A1(n_8_0_3290), .A2(n_8_0_6995), .ZN(n_8_0_1598));
   OAI211_X1 i_8_0_1372 (.A(n_8_0_1602), .B(n_8_0_3306), .C1(n_8_0_3326), 
      .C2(n_8_0_1603), .ZN(n_8_0_1601));
   AOI22_X1 i_8_0_1373 (.A1(n_8_0_1606), .A2(n_8_0_3319), .B1(n_8_0_3326), 
      .B2(in_data[12]), .ZN(n_8_0_1602));
   AOI21_X1 i_8_0_1374 (.A(n_8_0_1604), .B1(n_8_0_3320), .B2(in_data[16]), 
      .ZN(n_8_0_1603));
   NOR2_X1 i_8_0_1375 (.A1(n_8_0_3320), .A2(n_8_0_1605), .ZN(n_8_0_1604));
   NAND2_X1 i_8_0_1376 (.A1(n_8_0_3322), .A2(in_data[20]), .ZN(n_8_0_1605));
   MUX2_X1 i_8_0_1377 (.A(in_data[28]), .B(in_data[24]), .S(n_8_0_3316), 
      .Z(n_8_0_1606));
   OAI21_X1 i_8_0_1380 (.A(n_8_0_1609), .B1(n_8_0_1611), .B2(n_8_0_3352), 
      .ZN(n_8_0_1608));
   AOI21_X1 i_8_0_1381 (.A(n_8_0_3350), .B1(n_8_0_3352), .B2(n_8_0_6991), 
      .ZN(n_8_0_1609));
   AOI21_X1 i_8_0_1382 (.A(n_8_0_3346), .B1(n_8_0_3350), .B2(in_data[8]), 
      .ZN(n_8_0_1610));
   NOR2_X1 i_8_0_1383 (.A1(n_8_0_1613), .A2(n_8_0_1612), .ZN(n_8_0_1611));
   NOR2_X1 i_8_0_1384 (.A1(in_data[16]), .A2(n_8_0_3333), .ZN(n_8_0_1612));
   AOI21_X1 i_8_0_1385 (.A(n_8_0_1614), .B1(n_8_0_1615), .B2(n_8_0_3343), 
      .ZN(n_8_0_1613));
   OAI21_X1 i_8_0_1386 (.A(n_8_0_3333), .B1(n_8_0_3343), .B2(n_8_0_6993), 
      .ZN(n_8_0_1614));
   MUX2_X1 i_8_0_1387 (.A(in_data[24]), .B(in_data[28]), .S(n_8_0_3340), 
      .Z(n_8_0_1615));
   OAI21_X1 i_8_0_1391 (.A(n_8_0_3365), .B1(n_8_0_3372), .B2(n_8_0_6990), 
      .ZN(n_8_0_1618));
   OAI21_X1 i_8_0_1392 (.A(n_8_0_1620), .B1(n_8_0_1621), .B2(n_8_0_3367), 
      .ZN(n_8_0_1619));
   NAND2_X1 i_8_0_1393 (.A1(n_8_0_3367), .A2(in_data[12]), .ZN(n_8_0_1620));
   AOI21_X1 i_8_0_1394 (.A(n_8_0_1622), .B1(n_8_0_1623), .B2(n_8_0_3369), 
      .ZN(n_8_0_1621));
   NOR2_X1 i_8_0_1395 (.A1(n_8_0_3369), .A2(n_8_0_6992), .ZN(n_8_0_1622));
   OAI21_X1 i_8_0_1396 (.A(n_8_0_1624), .B1(n_8_0_3363), .B2(n_8_0_6993), 
      .ZN(n_8_0_1623));
   NAND2_X1 i_8_0_1397 (.A1(n_8_0_3363), .A2(n_8_0_1625), .ZN(n_8_0_1624));
   MUX2_X1 i_8_0_1398 (.A(in_data[24]), .B(in_data[28]), .S(n_8_0_3360), 
      .Z(n_8_0_1625));
   OAI22_X1 i_8_0_1399 (.A1(n_8_0_1627), .A2(n_8_0_1626), .B1(n_8_0_6988), 
      .B2(n_8_0_1637), .ZN(n_16));
   OAI21_X1 i_8_0_1400 (.A(n_8_0_1637), .B1(n_8_0_3385), .B2(in_data[4]), 
      .ZN(n_8_0_1626));
   AOI21_X1 i_8_0_1401 (.A(n_8_0_1628), .B1(n_8_0_1631), .B2(n_8_0_1630), 
      .ZN(n_8_0_1627));
   NAND2_X1 i_8_0_1402 (.A1(n_8_0_1629), .A2(n_8_0_3385), .ZN(n_8_0_1628));
   NAND2_X1 i_8_0_1403 (.A1(in_data[8]), .A2(n_8_0_3388), .ZN(n_8_0_1629));
   AOI21_X1 i_8_0_1404 (.A(n_8_0_3388), .B1(n_8_0_3404), .B2(n_8_0_6991), 
      .ZN(n_8_0_1630));
   OR2_X1 i_8_0_1405 (.A1(n_8_0_1632), .A2(n_8_0_3404), .ZN(n_8_0_1631));
   AOI21_X1 i_8_0_1406 (.A(n_8_0_1633), .B1(n_8_0_3400), .B2(n_8_0_6992), 
      .ZN(n_8_0_1632));
   NOR2_X1 i_8_0_1407 (.A1(n_8_0_3400), .A2(n_8_0_1634), .ZN(n_8_0_1633));
   AOI21_X1 i_8_0_1408 (.A(n_8_0_1635), .B1(n_8_0_3391), .B2(n_8_0_6993), 
      .ZN(n_8_0_1634));
   AOI211_X1 i_8_0_1409 (.A(n_8_0_3391), .B(n_8_0_1636), .C1(in_data[24]), 
      .C2(n_8_0_3394), .ZN(n_8_0_1635));
   NOR2_X1 i_8_0_1410 (.A1(n_8_0_6995), .A2(n_8_0_3394), .ZN(n_8_0_1636));
   OAI21_X1 i_8_0_1411 (.A(n_8_0_3397), .B1(n_8_0_6729), .B2(n_8_0_3398), 
      .ZN(n_8_0_1637));
   MUX2_X1 i_8_0_1412 (.A(n_8_0_1638), .B(in_data[0]), .S(n_8_0_3409), .Z(n_17));
   OAI21_X1 i_8_0_1413 (.A(n_8_0_1639), .B1(n_8_0_3418), .B2(n_8_0_6989), 
      .ZN(n_8_0_1638));
   OAI221_X1 i_8_0_1414 (.A(n_8_0_3418), .B1(n_8_0_3421), .B2(in_data[8]), 
      .C1(n_8_0_1640), .C2(n_8_0_1641), .ZN(n_8_0_1639));
   OAI21_X1 i_8_0_1415 (.A(n_8_0_3421), .B1(n_8_0_1642), .B2(n_8_0_3424), 
      .ZN(n_8_0_1640));
   OAI21_X1 i_8_0_1416 (.A(n_8_0_1645), .B1(n_8_0_3428), .B2(n_8_0_6991), 
      .ZN(n_8_0_1641));
   INV_X1 i_8_0_1417 (.A(n_8_0_1643), .ZN(n_8_0_1642));
   OAI21_X1 i_8_0_1418 (.A(n_8_0_1644), .B1(n_8_0_3413), .B2(n_8_0_6995), 
      .ZN(n_8_0_1643));
   NAND2_X1 i_8_0_1419 (.A1(in_data[24]), .A2(n_8_0_3413), .ZN(n_8_0_1644));
   OAI211_X1 i_8_0_1420 (.A(n_8_0_3428), .B(n_8_0_1646), .C1(in_data[16]), 
      .C2(n_8_0_3431), .ZN(n_8_0_1645));
   OAI21_X1 i_8_0_1421 (.A(n_8_0_3431), .B1(n_8_0_3425), .B2(n_8_0_6993), 
      .ZN(n_8_0_1646));
   OAI21_X1 i_8_0_1422 (.A(n_8_0_1647), .B1(n_8_0_3439), .B2(n_8_0_6988), 
      .ZN(n_18));
   OAI211_X1 i_8_0_1423 (.A(n_8_0_3439), .B(n_8_0_1648), .C1(n_8_0_1649), 
      .C2(n_8_0_3457), .ZN(n_8_0_1647));
   NAND2_X1 i_8_0_1424 (.A1(n_8_0_3457), .A2(n_8_0_6989), .ZN(n_8_0_1648));
   OAI21_X1 i_8_0_1425 (.A(n_8_0_1650), .B1(n_8_0_3455), .B2(n_8_0_6990), 
      .ZN(n_8_0_1649));
   OAI211_X1 i_8_0_1426 (.A(n_8_0_1651), .B(n_8_0_3455), .C1(in_data[12]), 
      .C2(n_8_0_3453), .ZN(n_8_0_1650));
   OAI211_X1 i_8_0_1427 (.A(n_8_0_1652), .B(n_8_0_3453), .C1(n_8_0_6992), 
      .C2(n_8_0_3447), .ZN(n_8_0_1651));
   OAI211_X1 i_8_0_1428 (.A(n_8_0_1653), .B(n_8_0_3447), .C1(in_data[20]), 
      .C2(n_8_0_3442), .ZN(n_8_0_1652));
   NAND2_X1 i_8_0_1429 (.A1(n_8_0_3442), .A2(n_8_0_1654), .ZN(n_8_0_1653));
   OAI21_X1 i_8_0_1430 (.A(n_8_0_1655), .B1(n_8_0_3437), .B2(in_data[24]), 
      .ZN(n_8_0_1654));
   NAND2_X1 i_8_0_1431 (.A1(n_8_0_3437), .A2(n_8_0_6995), .ZN(n_8_0_1655));
   AOI21_X1 i_8_0_1435 (.A(n_8_0_1659), .B1(n_8_0_1660), .B2(n_8_0_3481), 
      .ZN(n_8_0_1658));
   NOR2_X1 i_8_0_1436 (.A1(n_8_0_3481), .A2(n_8_0_6990), .ZN(n_8_0_1659));
   OAI21_X1 i_8_0_1437 (.A(n_8_0_1661), .B1(n_8_0_3479), .B2(n_8_0_6991), 
      .ZN(n_8_0_1660));
   OAI211_X1 i_8_0_1438 (.A(n_8_0_3479), .B(n_8_0_1662), .C1(n_8_0_1663), 
      .C2(n_8_0_3463), .ZN(n_8_0_1661));
   NAND2_X1 i_8_0_1439 (.A1(n_8_0_6992), .A2(n_8_0_3463), .ZN(n_8_0_1662));
   AOI21_X1 i_8_0_1440 (.A(n_8_0_1664), .B1(n_8_0_3468), .B2(n_8_0_6993), 
      .ZN(n_8_0_1663));
   NOR2_X1 i_8_0_1441 (.A1(n_8_0_1665), .A2(n_8_0_3468), .ZN(n_8_0_1664));
   MUX2_X1 i_8_0_1442 (.A(in_data[28]), .B(in_data[24]), .S(n_8_0_3471), 
      .Z(n_8_0_1665));
   AOI22_X1 i_8_0_1443 (.A1(n_8_0_1668), .A2(n_8_0_1666), .B1(n_8_0_1667), 
      .B2(n_8_0_6988), .ZN(n_19));
   AOI21_X1 i_8_0_1444 (.A(n_8_0_1667), .B1(n_8_0_3511), .B2(in_data[4]), 
      .ZN(n_8_0_1666));
   OAI21_X1 i_8_0_1445 (.A(n_8_0_3497), .B1(n_8_0_3496), .B2(n_8_0_6730), 
      .ZN(n_8_0_1667));
   OAI21_X1 i_8_0_1446 (.A(n_8_0_1669), .B1(n_8_0_1670), .B2(n_8_0_3506), 
      .ZN(n_8_0_1668));
   AOI21_X1 i_8_0_1447 (.A(n_8_0_3511), .B1(n_8_0_3506), .B2(n_8_0_6990), 
      .ZN(n_8_0_1669));
   MUX2_X1 i_8_0_1448 (.A(in_data[12]), .B(n_8_0_1671), .S(n_8_0_3503), .Z(
      n_8_0_1670));
   AOI21_X1 i_8_0_1449 (.A(n_8_0_1672), .B1(n_8_0_3514), .B2(n_8_0_6992), 
      .ZN(n_8_0_1671));
   NOR2_X1 i_8_0_1450 (.A1(n_8_0_1673), .A2(n_8_0_3514), .ZN(n_8_0_1672));
   MUX2_X1 i_8_0_1451 (.A(in_data[20]), .B(n_8_0_1674), .S(n_8_0_3491), .Z(
      n_8_0_1673));
   OAI21_X1 i_8_0_1452 (.A(n_8_0_1675), .B1(n_8_0_3500), .B2(n_8_0_6995), 
      .ZN(n_8_0_1674));
   NAND2_X1 i_8_0_1453 (.A1(n_8_0_3500), .A2(in_data[24]), .ZN(n_8_0_1675));
   OAI21_X1 i_8_0_1454 (.A(n_8_0_1676), .B1(n_8_0_3527), .B2(n_8_0_6988), 
      .ZN(n_20));
   OAI211_X1 i_8_0_1455 (.A(n_8_0_3527), .B(n_8_0_1685), .C1(n_8_0_1677), 
      .C2(n_8_0_3541), .ZN(n_8_0_1676));
   AOI21_X1 i_8_0_1456 (.A(n_8_0_1678), .B1(n_8_0_3534), .B2(n_8_0_6990), 
      .ZN(n_8_0_1677));
   AOI21_X1 i_8_0_1457 (.A(n_8_0_3534), .B1(n_8_0_1680), .B2(n_8_0_1679), 
      .ZN(n_8_0_1678));
   OR2_X1 i_8_0_1458 (.A1(in_data[12]), .A2(n_8_0_3536), .ZN(n_8_0_1679));
   OAI211_X1 i_8_0_1459 (.A(n_8_0_1681), .B(n_8_0_3536), .C1(n_8_0_6992), 
      .C2(n_8_0_3530), .ZN(n_8_0_1680));
   OAI221_X1 i_8_0_1460 (.A(n_8_0_3530), .B1(n_8_0_3524), .B2(in_data[20]), 
      .C1(n_8_0_1682), .C2(n_8_0_1684), .ZN(n_8_0_1681));
   NAND2_X1 i_8_0_1461 (.A1(n_8_0_3524), .A2(n_8_0_1683), .ZN(n_8_0_1682));
   NAND2_X1 i_8_0_1462 (.A1(n_8_0_3520), .A2(in_data[24]), .ZN(n_8_0_1683));
   NOR2_X1 i_8_0_1463 (.A1(n_8_0_6995), .A2(n_8_0_3520), .ZN(n_8_0_1684));
   NAND2_X1 i_8_0_1464 (.A1(n_8_0_6989), .A2(n_8_0_3541), .ZN(n_8_0_1685));
   OAI21_X1 i_8_0_1465 (.A(n_8_0_1686), .B1(n_8_0_3554), .B2(n_8_0_6988), 
      .ZN(n_21));
   OAI211_X1 i_8_0_1466 (.A(n_8_0_3554), .B(n_8_0_1687), .C1(n_8_0_1688), 
      .C2(n_8_0_3551), .ZN(n_8_0_1686));
   NAND2_X1 i_8_0_1467 (.A1(n_8_0_3551), .A2(n_8_0_6989), .ZN(n_8_0_1687));
   MUX2_X1 i_8_0_1468 (.A(n_8_0_1689), .B(in_data[8]), .S(n_8_0_3557), .Z(
      n_8_0_1688));
   OAI21_X1 i_8_0_1469 (.A(n_8_0_1690), .B1(n_8_0_3558), .B2(n_8_0_6991), 
      .ZN(n_8_0_1689));
   OAI211_X1 i_8_0_1470 (.A(n_8_0_3558), .B(n_8_0_1691), .C1(n_8_0_1692), 
      .C2(n_8_0_3566), .ZN(n_8_0_1690));
   NAND2_X1 i_8_0_1471 (.A1(n_8_0_6992), .A2(n_8_0_3566), .ZN(n_8_0_1691));
   AOI21_X1 i_8_0_1472 (.A(n_8_0_1693), .B1(n_8_0_3561), .B2(n_8_0_6993), 
      .ZN(n_8_0_1692));
   AOI211_X1 i_8_0_1473 (.A(n_8_0_3561), .B(n_8_0_1694), .C1(n_8_0_3548), 
      .C2(in_data[28]), .ZN(n_8_0_1693));
   NOR2_X1 i_8_0_1474 (.A1(n_8_0_3548), .A2(n_8_0_6994), .ZN(n_8_0_1694));
   OAI22_X1 i_8_0_1475 (.A1(n_8_0_1696), .A2(n_8_0_1695), .B1(n_8_0_6988), 
      .B2(n_8_0_3580), .ZN(n_22));
   OAI21_X1 i_8_0_1476 (.A(n_8_0_3580), .B1(n_8_0_3574), .B2(in_data[4]), 
      .ZN(n_8_0_1695));
   NOR3_X1 i_8_0_1477 (.A1(n_8_0_3576), .A2(n_8_0_3575), .A3(n_8_0_1697), 
      .ZN(n_8_0_1696));
   AOI21_X1 i_8_0_1478 (.A(n_8_0_1698), .B1(n_8_0_3594), .B2(n_8_0_6990), 
      .ZN(n_8_0_1697));
   AOI211_X1 i_8_0_1479 (.A(n_8_0_3594), .B(n_8_0_1699), .C1(n_8_0_3577), 
      .C2(in_data[12]), .ZN(n_8_0_1698));
   AOI211_X1 i_8_0_1480 (.A(n_8_0_3577), .B(n_8_0_1700), .C1(n_8_0_1701), 
      .C2(n_8_0_3591), .ZN(n_8_0_1699));
   NOR2_X1 i_8_0_1481 (.A1(in_data[16]), .A2(n_8_0_3591), .ZN(n_8_0_1700));
   OAI21_X1 i_8_0_1482 (.A(n_8_0_1702), .B1(n_8_0_3587), .B2(in_data[20]), 
      .ZN(n_8_0_1701));
   OAI211_X1 i_8_0_1483 (.A(n_8_0_3587), .B(n_8_0_1703), .C1(n_8_0_3583), 
      .C2(n_8_0_6994), .ZN(n_8_0_1702));
   NAND2_X1 i_8_0_1484 (.A1(n_8_0_3583), .A2(in_data[28]), .ZN(n_8_0_1703));
   OAI22_X1 i_8_0_1485 (.A1(n_8_0_1705), .A2(n_8_0_1704), .B1(n_8_0_6988), 
      .B2(n_8_0_3601), .ZN(n_23));
   OAI21_X1 i_8_0_1486 (.A(n_8_0_3601), .B1(n_8_0_3631), .B2(in_data[4]), 
      .ZN(n_8_0_1704));
   AOI211_X1 i_8_0_1487 (.A(n_8_0_3630), .B(n_8_0_1706), .C1(n_8_0_3615), 
      .C2(in_data[8]), .ZN(n_8_0_1705));
   NOR3_X1 i_8_0_1488 (.A1(n_8_0_1708), .A2(n_8_0_1707), .A3(n_8_0_3615), 
      .ZN(n_8_0_1706));
   NOR2_X1 i_8_0_1489 (.A1(in_data[12]), .A2(n_8_0_3628), .ZN(n_8_0_1707));
   AOI21_X1 i_8_0_1490 (.A(n_8_0_1709), .B1(n_8_0_1710), .B2(n_8_0_3625), 
      .ZN(n_8_0_1708));
   OAI21_X1 i_8_0_1491 (.A(n_8_0_3628), .B1(n_8_0_3625), .B2(n_8_0_6992), 
      .ZN(n_8_0_1709));
   OAI22_X1 i_8_0_1492 (.A1(n_8_0_1712), .A2(n_8_0_1711), .B1(n_8_0_6993), 
      .B2(n_8_0_3612), .ZN(n_8_0_1710));
   OAI21_X1 i_8_0_1493 (.A(n_8_0_3612), .B1(n_8_0_3606), .B2(in_data[28]), 
      .ZN(n_8_0_1711));
   NOR2_X1 i_8_0_1494 (.A1(in_data[24]), .A2(n_8_0_3607), .ZN(n_8_0_1712));
   OAI21_X1 i_8_0_1495 (.A(n_8_0_1713), .B1(n_8_0_1714), .B2(n_8_0_3655), 
      .ZN(n_24));
   NAND2_X1 i_8_0_1496 (.A1(n_8_0_3655), .A2(in_data[0]), .ZN(n_8_0_1713));
   OAI21_X1 i_8_0_1497 (.A(n_8_0_1715), .B1(n_8_0_3644), .B2(in_data[4]), 
      .ZN(n_8_0_1714));
   NAND3_X1 i_8_0_1498 (.A1(n_8_0_1717), .A2(n_8_0_1716), .A3(n_8_0_3644), 
      .ZN(n_8_0_1715));
   NAND2_X1 i_8_0_1499 (.A1(in_data[8]), .A2(n_8_0_3660), .ZN(n_8_0_1716));
   OAI21_X1 i_8_0_1500 (.A(n_8_0_1718), .B1(n_8_0_1722), .B2(n_8_0_3666), 
      .ZN(n_8_0_1717));
   AOI21_X1 i_8_0_1501 (.A(n_8_0_3660), .B1(n_8_0_1719), .B2(n_8_0_3666), 
      .ZN(n_8_0_1718));
   INV_X1 i_8_0_1502 (.A(n_8_0_1720), .ZN(n_8_0_1719));
   OAI21_X1 i_8_0_1503 (.A(n_8_0_1721), .B1(n_8_0_3667), .B2(n_8_0_6991), 
      .ZN(n_8_0_1720));
   NAND2_X1 i_8_0_1504 (.A1(in_data[16]), .A2(n_8_0_3667), .ZN(n_8_0_1721));
   AOI21_X1 i_8_0_1505 (.A(n_8_0_1723), .B1(n_8_0_3636), .B2(n_8_0_6993), 
      .ZN(n_8_0_1722));
   AOI211_X1 i_8_0_1506 (.A(n_8_0_3636), .B(n_8_0_1724), .C1(in_data[24]), 
      .C2(n_8_0_3649), .ZN(n_8_0_1723));
   NOR2_X1 i_8_0_1507 (.A1(n_8_0_3649), .A2(n_8_0_6995), .ZN(n_8_0_1724));
   OAI21_X1 i_8_0_1508 (.A(n_8_0_1725), .B1(n_8_0_3689), .B2(n_8_0_6988), 
      .ZN(n_25));
   OAI211_X1 i_8_0_1509 (.A(n_8_0_1726), .B(n_8_0_3689), .C1(in_data[4]), 
      .C2(n_8_0_3687), .ZN(n_8_0_1725));
   OAI211_X1 i_8_0_1510 (.A(n_8_0_3687), .B(n_8_0_1727), .C1(n_8_0_1728), 
      .C2(n_8_0_3688), .ZN(n_8_0_1726));
   NAND2_X1 i_8_0_1511 (.A1(in_data[8]), .A2(n_8_0_3688), .ZN(n_8_0_1727));
   INV_X1 i_8_0_1512 (.A(n_8_0_1729), .ZN(n_8_0_1728));
   AOI21_X1 i_8_0_1513 (.A(n_8_0_1730), .B1(n_8_0_3681), .B2(n_8_0_6991), 
      .ZN(n_8_0_1729));
   AOI211_X1 i_8_0_1514 (.A(n_8_0_3681), .B(n_8_0_1731), .C1(in_data[16]), 
      .C2(n_8_0_3682), .ZN(n_8_0_1730));
   AOI211_X1 i_8_0_1515 (.A(n_8_0_3682), .B(n_8_0_1732), .C1(n_8_0_6993), 
      .C2(n_8_0_3694), .ZN(n_8_0_1731));
   AOI211_X1 i_8_0_1516 (.A(n_8_0_1733), .B(n_8_0_3694), .C1(in_data[24]), 
      .C2(n_8_0_3693), .ZN(n_8_0_1732));
   NOR2_X1 i_8_0_1517 (.A1(n_8_0_6995), .A2(n_8_0_3693), .ZN(n_8_0_1733));
   AOI21_X1 i_8_0_1523 (.A(n_8_0_3702), .B1(n_8_0_3721), .B2(n_8_0_6991), 
      .ZN(n_8_0_1738));
   OAI21_X1 i_8_0_1524 (.A(n_8_0_1740), .B1(n_8_0_1741), .B2(n_8_0_3705), 
      .ZN(n_8_0_1739));
   NAND2_X1 i_8_0_1525 (.A1(n_8_0_3705), .A2(in_data[16]), .ZN(n_8_0_1740));
   OAI21_X1 i_8_0_1526 (.A(n_8_0_1742), .B1(n_8_0_1743), .B2(n_8_0_3718), 
      .ZN(n_8_0_1741));
   NAND2_X1 i_8_0_1527 (.A1(n_8_0_6993), .A2(n_8_0_3718), .ZN(n_8_0_1742));
   OAI21_X1 i_8_0_1528 (.A(n_8_0_1744), .B1(n_8_0_3714), .B2(n_8_0_6995), 
      .ZN(n_8_0_1743));
   NAND2_X1 i_8_0_1529 (.A1(n_8_0_3714), .A2(in_data[24]), .ZN(n_8_0_1744));
   MUX2_X1 i_8_0_1530 (.A(n_8_0_1745), .B(in_data[0]), .S(n_8_0_3732), .Z(n_26));
   AOI21_X1 i_8_0_1531 (.A(n_8_0_1746), .B1(n_8_0_3736), .B2(n_8_0_6989), 
      .ZN(n_8_0_1745));
   AOI221_X1 i_8_0_1532 (.A(n_8_0_3736), .B1(n_8_0_1748), .B2(n_8_0_1747), 
      .C1(n_8_0_3739), .C2(in_data[8]), .ZN(n_8_0_1746));
   AOI21_X1 i_8_0_1533 (.A(n_8_0_3739), .B1(n_8_0_3726), .B2(n_8_0_6991), 
      .ZN(n_8_0_1747));
   OAI21_X1 i_8_0_1534 (.A(n_8_0_1749), .B1(n_8_0_1750), .B2(n_8_0_3729), 
      .ZN(n_8_0_1748));
   AOI21_X1 i_8_0_1535 (.A(n_8_0_3726), .B1(n_8_0_3729), .B2(in_data[16]), 
      .ZN(n_8_0_1749));
   OAI21_X1 i_8_0_1536 (.A(n_8_0_1751), .B1(n_8_0_3746), .B2(in_data[20]), 
      .ZN(n_8_0_1750));
   OAI211_X1 i_8_0_1537 (.A(n_8_0_3746), .B(n_8_0_1752), .C1(n_8_0_6995), 
      .C2(n_8_0_3749), .ZN(n_8_0_1751));
   NAND2_X1 i_8_0_1538 (.A1(n_8_0_3749), .A2(in_data[24]), .ZN(n_8_0_1752));
   AOI21_X1 i_8_0_1543 (.A(n_8_0_1757), .B1(n_8_0_3752), .B2(n_8_0_6991), 
      .ZN(n_8_0_1756));
   AOI211_X1 i_8_0_1544 (.A(n_8_0_3752), .B(n_8_0_1758), .C1(in_data[16]), 
      .C2(n_8_0_3767), .ZN(n_8_0_1757));
   AOI211_X1 i_8_0_1545 (.A(n_8_0_3767), .B(n_8_0_1759), .C1(n_8_0_1760), 
      .C2(n_8_0_3779), .ZN(n_8_0_1758));
   NOR2_X1 i_8_0_1546 (.A1(in_data[20]), .A2(n_8_0_3779), .ZN(n_8_0_1759));
   OAI21_X1 i_8_0_1547 (.A(n_8_0_1761), .B1(n_8_0_3776), .B2(in_data[28]), 
      .ZN(n_8_0_1760));
   NAND2_X1 i_8_0_1548 (.A1(n_8_0_6994), .A2(n_8_0_3776), .ZN(n_8_0_1761));
   OAI21_X1 i_8_0_1549 (.A(n_8_0_1762), .B1(n_8_0_3795), .B2(n_8_0_6988), 
      .ZN(n_27));
   OAI211_X1 i_8_0_1550 (.A(n_8_0_3795), .B(n_8_0_1763), .C1(n_8_0_1766), 
      .C2(n_8_0_1764), .ZN(n_8_0_1762));
   NAND2_X1 i_8_0_1551 (.A1(n_8_0_6989), .A2(n_8_0_3805), .ZN(n_8_0_1763));
   INV_X1 i_8_0_1552 (.A(n_8_0_1765), .ZN(n_8_0_1764));
   AOI21_X1 i_8_0_1553 (.A(n_8_0_3805), .B1(n_8_0_3800), .B2(in_data[8]), 
      .ZN(n_8_0_1765));
   AOI211_X1 i_8_0_1554 (.A(n_8_0_3800), .B(n_8_0_1767), .C1(n_8_0_1768), 
      .C2(n_8_0_3793), .ZN(n_8_0_1766));
   NOR2_X1 i_8_0_1555 (.A1(in_data[12]), .A2(n_8_0_3793), .ZN(n_8_0_1767));
   INV_X1 i_8_0_1556 (.A(n_8_0_1769), .ZN(n_8_0_1768));
   MUX2_X1 i_8_0_1557 (.A(in_data[16]), .B(n_8_0_1770), .S(n_8_0_3807), .Z(
      n_8_0_1769));
   AOI21_X1 i_8_0_1558 (.A(n_8_0_1771), .B1(n_8_0_1772), .B2(n_8_0_3788), 
      .ZN(n_8_0_1770));
   NOR2_X1 i_8_0_1559 (.A1(in_data[20]), .A2(n_8_0_3788), .ZN(n_8_0_1771));
   OAI21_X1 i_8_0_1560 (.A(n_8_0_1773), .B1(n_8_0_3785), .B2(in_data[28]), 
      .ZN(n_8_0_1772));
   NAND2_X1 i_8_0_1561 (.A1(n_8_0_6994), .A2(n_8_0_3785), .ZN(n_8_0_1773));
   MUX2_X1 i_8_0_1564 (.A(n_8_0_1776), .B(in_data[8]), .S(n_8_0_3822), .Z(
      n_8_0_1775));
   MUX2_X1 i_8_0_1565 (.A(n_8_0_1777), .B(in_data[12]), .S(n_8_0_3835), .Z(
      n_8_0_1776));
   AOI21_X1 i_8_0_1566 (.A(n_8_0_1778), .B1(n_8_0_3816), .B2(n_8_0_6992), 
      .ZN(n_8_0_1777));
   NOR2_X1 i_8_0_1567 (.A1(n_8_0_1779), .A2(n_8_0_3816), .ZN(n_8_0_1778));
   AOI21_X1 i_8_0_1568 (.A(n_8_0_1780), .B1(n_8_0_3827), .B2(n_8_0_6993), 
      .ZN(n_8_0_1779));
   AOI211_X1 i_8_0_1569 (.A(n_8_0_1781), .B(n_8_0_3827), .C1(n_8_0_3832), 
      .C2(in_data[28]), .ZN(n_8_0_1780));
   NOR2_X1 i_8_0_1570 (.A1(n_8_0_3832), .A2(n_8_0_6994), .ZN(n_8_0_1781));
   AOI21_X1 i_8_0_1574 (.A(n_8_0_3855), .B1(n_8_0_3844), .B2(in_data[12]), 
      .ZN(n_8_0_1784));
   NAND2_X1 i_8_0_1575 (.A1(n_8_0_3843), .A2(n_8_0_1786), .ZN(n_8_0_1785));
   MUX2_X1 i_8_0_1576 (.A(in_data[16]), .B(n_8_0_1787), .S(n_8_0_3860), .Z(
      n_8_0_1786));
   AOI21_X1 i_8_0_1577 (.A(n_8_0_1788), .B1(n_8_0_1789), .B2(n_8_0_3849), 
      .ZN(n_8_0_1787));
   NOR2_X1 i_8_0_1578 (.A1(in_data[20]), .A2(n_8_0_3849), .ZN(n_8_0_1788));
   OAI21_X1 i_8_0_1579 (.A(n_8_0_1790), .B1(n_8_0_3851), .B2(in_data[28]), 
      .ZN(n_8_0_1789));
   NAND2_X1 i_8_0_1580 (.A1(n_8_0_6994), .A2(n_8_0_3851), .ZN(n_8_0_1790));
   OAI22_X1 i_8_0_1581 (.A1(n_8_0_1792), .A2(n_8_0_1791), .B1(n_8_0_6988), 
      .B2(n_8_0_3883), .ZN(n_28));
   OAI21_X1 i_8_0_1582 (.A(n_8_0_3883), .B1(n_8_0_3870), .B2(in_data[4]), 
      .ZN(n_8_0_1791));
   AOI211_X1 i_8_0_1583 (.A(n_8_0_3871), .B(n_8_0_1793), .C1(in_data[8]), 
      .C2(n_8_0_3889), .ZN(n_8_0_1792));
   AOI211_X1 i_8_0_1584 (.A(n_8_0_3889), .B(n_8_0_1794), .C1(n_8_0_3867), 
      .C2(n_8_0_6991), .ZN(n_8_0_1793));
   NOR2_X1 i_8_0_1585 (.A1(n_8_0_3867), .A2(n_8_0_1795), .ZN(n_8_0_1794));
   MUX2_X1 i_8_0_1586 (.A(n_8_0_1796), .B(in_data[16]), .S(n_8_0_3874), .Z(
      n_8_0_1795));
   OAI21_X1 i_8_0_1587 (.A(n_8_0_1797), .B1(n_8_0_1798), .B2(n_8_0_3887), 
      .ZN(n_8_0_1796));
   NAND2_X1 i_8_0_1588 (.A1(n_8_0_3887), .A2(in_data[20]), .ZN(n_8_0_1797));
   OAI21_X1 i_8_0_1589 (.A(n_8_0_1799), .B1(n_8_0_3878), .B2(in_data[28]), 
      .ZN(n_8_0_1798));
   NAND2_X1 i_8_0_1590 (.A1(n_8_0_6994), .A2(n_8_0_3878), .ZN(n_8_0_1799));
   OAI22_X1 i_8_0_1591 (.A1(n_8_0_1801), .A2(n_8_0_1800), .B1(n_8_0_6988), 
      .B2(n_8_0_3904), .ZN(n_29));
   OAI21_X1 i_8_0_1592 (.A(n_8_0_3904), .B1(n_8_0_3914), .B2(in_data[4]), 
      .ZN(n_8_0_1800));
   AOI211_X1 i_8_0_1593 (.A(n_8_0_3915), .B(n_8_0_1802), .C1(n_8_0_3899), 
      .C2(in_data[8]), .ZN(n_8_0_1801));
   AOI211_X1 i_8_0_1594 (.A(n_8_0_3899), .B(n_8_0_1803), .C1(n_8_0_3895), 
      .C2(n_8_0_6991), .ZN(n_8_0_1802));
   NOR2_X1 i_8_0_1595 (.A1(n_8_0_1804), .A2(n_8_0_3895), .ZN(n_8_0_1803));
   AOI21_X1 i_8_0_1596 (.A(n_8_0_1805), .B1(n_8_0_3913), .B2(n_8_0_6992), 
      .ZN(n_8_0_1804));
   AOI211_X1 i_8_0_1597 (.A(n_8_0_3913), .B(n_8_0_1806), .C1(n_8_0_3910), 
      .C2(in_data[20]), .ZN(n_8_0_1805));
   AOI211_X1 i_8_0_1598 (.A(n_8_0_1807), .B(n_8_0_3910), .C1(n_8_0_6994), 
      .C2(n_8_0_3893), .ZN(n_8_0_1806));
   NOR2_X1 i_8_0_1599 (.A1(n_8_0_3893), .A2(in_data[28]), .ZN(n_8_0_1807));
   OAI21_X1 i_8_0_1600 (.A(n_8_0_1808), .B1(n_8_0_3939), .B2(n_8_0_6988), 
      .ZN(n_30));
   NAND2_X1 i_8_0_1601 (.A1(n_8_0_3939), .A2(n_8_0_1809), .ZN(n_8_0_1808));
   AOI22_X1 i_8_0_1602 (.A1(n_8_0_1811), .A2(n_8_0_1810), .B1(n_8_0_6989), 
      .B2(n_8_0_3921), .ZN(n_8_0_1809));
   AOI21_X1 i_8_0_1603 (.A(n_8_0_3921), .B1(n_8_0_3931), .B2(in_data[8]), 
      .ZN(n_8_0_1810));
   OAI21_X1 i_8_0_1604 (.A(n_8_0_1812), .B1(n_8_0_1813), .B2(n_8_0_3928), 
      .ZN(n_8_0_1811));
   AOI21_X1 i_8_0_1605 (.A(n_8_0_3931), .B1(n_8_0_3928), .B2(n_8_0_6991), 
      .ZN(n_8_0_1812));
   AOI21_X1 i_8_0_1606 (.A(n_8_0_1814), .B1(n_8_0_3923), .B2(n_8_0_6992), 
      .ZN(n_8_0_1813));
   AOI211_X1 i_8_0_1607 (.A(n_8_0_3923), .B(n_8_0_1815), .C1(in_data[20]), 
      .C2(n_8_0_3934), .ZN(n_8_0_1814));
   AOI211_X1 i_8_0_1608 (.A(n_8_0_1816), .B(n_8_0_3934), .C1(n_8_0_6995), 
      .C2(n_8_0_3925), .ZN(n_8_0_1815));
   NOR2_X1 i_8_0_1609 (.A1(in_data[24]), .A2(n_8_0_3925), .ZN(n_8_0_1816));
   OAI22_X1 i_8_0_1610 (.A1(n_8_0_1818), .A2(n_8_0_1817), .B1(n_8_0_6988), 
      .B2(n_8_0_3967), .ZN(n_31));
   OAI21_X1 i_8_0_1611 (.A(n_8_0_3967), .B1(n_8_0_3958), .B2(in_data[4]), 
      .ZN(n_8_0_1817));
   AOI21_X1 i_8_0_1612 (.A(n_8_0_1819), .B1(n_8_0_1820), .B2(n_8_0_3961), 
      .ZN(n_8_0_1818));
   OAI21_X1 i_8_0_1613 (.A(n_8_0_3958), .B1(n_8_0_3961), .B2(n_8_0_6990), 
      .ZN(n_8_0_1819));
   OAI21_X1 i_8_0_1614 (.A(n_8_0_1821), .B1(n_8_0_3964), .B2(n_8_0_6991), 
      .ZN(n_8_0_1820));
   OAI211_X1 i_8_0_1615 (.A(n_8_0_3964), .B(n_8_0_1822), .C1(n_8_0_1823), 
      .C2(n_8_0_3953), .ZN(n_8_0_1821));
   NAND2_X1 i_8_0_1616 (.A1(n_8_0_6992), .A2(n_8_0_3953), .ZN(n_8_0_1822));
   AOI21_X1 i_8_0_1617 (.A(n_8_0_1824), .B1(n_8_0_3950), .B2(n_8_0_6993), 
      .ZN(n_8_0_1823));
   AOI211_X1 i_8_0_1618 (.A(n_8_0_3950), .B(n_8_0_1825), .C1(n_8_0_3945), 
      .C2(in_data[24]), .ZN(n_8_0_1824));
   NOR2_X1 i_8_0_1619 (.A1(n_8_0_6995), .A2(n_8_0_3945), .ZN(n_8_0_1825));
   MUX2_X1 i_8_0_1620 (.A(n_8_0_1826), .B(in_data[0]), .S(n_8_0_3989), .Z(n_32));
   AOI22_X1 i_8_0_1621 (.A1(n_8_0_1828), .A2(n_8_0_1827), .B1(n_8_0_6989), 
      .B2(n_8_0_3992), .ZN(n_8_0_1826));
   AOI21_X1 i_8_0_1622 (.A(n_8_0_3992), .B1(n_8_0_3976), .B2(in_data[8]), 
      .ZN(n_8_0_1827));
   OAI21_X1 i_8_0_1623 (.A(n_8_0_1833), .B1(n_8_0_1829), .B2(n_8_0_3974), 
      .ZN(n_8_0_1828));
   AOI21_X1 i_8_0_1624 (.A(n_8_0_1830), .B1(n_8_0_3979), .B2(n_8_0_6992), 
      .ZN(n_8_0_1829));
   AOI211_X1 i_8_0_1625 (.A(n_8_0_3979), .B(n_8_0_1831), .C1(in_data[20]), 
      .C2(n_8_0_3986), .ZN(n_8_0_1830));
   AOI211_X1 i_8_0_1626 (.A(n_8_0_1832), .B(n_8_0_3986), .C1(n_8_0_6994), 
      .C2(n_8_0_3981), .ZN(n_8_0_1831));
   NOR2_X1 i_8_0_1627 (.A1(n_8_0_3981), .A2(in_data[28]), .ZN(n_8_0_1832));
   AOI21_X1 i_8_0_1628 (.A(n_8_0_3976), .B1(n_8_0_3974), .B2(n_8_0_6991), 
      .ZN(n_8_0_1833));
   AOI21_X1 i_8_0_1629 (.A(n_8_0_1834), .B1(n_8_0_4001), .B2(n_8_0_6988), 
      .ZN(n_33));
   NOR2_X1 i_8_0_1630 (.A1(n_8_0_1835), .A2(n_8_0_4001), .ZN(n_8_0_1834));
   AOI21_X1 i_8_0_1631 (.A(n_8_0_1836), .B1(n_8_0_4004), .B2(n_8_0_6989), 
      .ZN(n_8_0_1835));
   NOR2_X1 i_8_0_1632 (.A1(n_8_0_4004), .A2(n_8_0_1837), .ZN(n_8_0_1836));
   MUX2_X1 i_8_0_1633 (.A(n_8_0_1838), .B(in_data[8]), .S(n_8_0_4013), .Z(
      n_8_0_1837));
   OAI21_X1 i_8_0_1634 (.A(n_8_0_1839), .B1(n_8_0_1840), .B2(n_8_0_4009), 
      .ZN(n_8_0_1838));
   NAND2_X1 i_8_0_1635 (.A1(in_data[12]), .A2(n_8_0_4009), .ZN(n_8_0_1839));
   MUX2_X1 i_8_0_1636 (.A(n_8_0_1841), .B(n_8_0_6992), .S(n_8_0_3998), .Z(
      n_8_0_1840));
   OAI21_X1 i_8_0_1637 (.A(n_8_0_1842), .B1(n_8_0_1843), .B2(n_8_0_4016), 
      .ZN(n_8_0_1841));
   NAND2_X1 i_8_0_1638 (.A1(n_8_0_6993), .A2(n_8_0_4016), .ZN(n_8_0_1842));
   AOI21_X1 i_8_0_1639 (.A(n_8_0_1844), .B1(n_8_0_4017), .B2(n_8_0_6995), 
      .ZN(n_8_0_1843));
   NOR2_X1 i_8_0_1640 (.A1(in_data[24]), .A2(n_8_0_4017), .ZN(n_8_0_1844));
   OAI21_X1 i_8_0_1641 (.A(n_8_0_1845), .B1(n_8_0_4022), .B2(n_8_0_6988), 
      .ZN(n_34));
   NAND3_X1 i_8_0_1642 (.A1(n_8_0_1847), .A2(n_8_0_1846), .A3(n_8_0_4022), 
      .ZN(n_8_0_1845));
   NAND2_X1 i_8_0_1643 (.A1(n_8_0_6989), .A2(n_8_0_4043), .ZN(n_8_0_1846));
   OAI21_X1 i_8_0_1644 (.A(n_8_0_1848), .B1(n_8_0_1849), .B2(n_8_0_4040), 
      .ZN(n_8_0_1847));
   AOI21_X1 i_8_0_1645 (.A(n_8_0_4043), .B1(n_8_0_4040), .B2(in_data[8]), 
      .ZN(n_8_0_1848));
   AOI221_X1 i_8_0_1646 (.A(n_8_0_1851), .B1(n_8_0_1850), .B2(n_8_0_4026), 
      .C1(n_8_0_1852), .C2(n_8_0_4025), .ZN(n_8_0_1849));
   NOR2_X1 i_8_0_1647 (.A1(n_8_0_4030), .A2(n_8_0_6992), .ZN(n_8_0_1850));
   NOR2_X1 i_8_0_1648 (.A1(n_8_0_4026), .A2(n_8_0_6991), .ZN(n_8_0_1851));
   OAI21_X1 i_8_0_1649 (.A(n_8_0_1853), .B1(n_8_0_4033), .B2(n_8_0_6993), 
      .ZN(n_8_0_1852));
   OAI211_X1 i_8_0_1650 (.A(n_8_0_4033), .B(n_8_0_1854), .C1(in_data[28]), 
      .C2(n_8_0_4035), .ZN(n_8_0_1853));
   NAND2_X1 i_8_0_1651 (.A1(n_8_0_6994), .A2(n_8_0_4035), .ZN(n_8_0_1854));
   OAI22_X1 i_8_0_1652 (.A1(n_8_0_1856), .A2(n_8_0_1855), .B1(n_8_0_6988), 
      .B2(n_8_0_4050), .ZN(n_35));
   OAI21_X1 i_8_0_1653 (.A(n_8_0_4050), .B1(n_8_0_4062), .B2(in_data[4]), 
      .ZN(n_8_0_1855));
   NOR2_X1 i_8_0_1654 (.A1(n_8_0_4063), .A2(n_8_0_1857), .ZN(n_8_0_1856));
   MUX2_X1 i_8_0_1655 (.A(n_8_0_1858), .B(in_data[8]), .S(n_8_0_4067), .Z(
      n_8_0_1857));
   MUX2_X1 i_8_0_1656 (.A(in_data[12]), .B(n_8_0_1859), .S(n_8_0_4056), .Z(
      n_8_0_1858));
   MUX2_X1 i_8_0_1657 (.A(n_8_0_1860), .B(in_data[16]), .S(n_8_0_4053), .Z(
      n_8_0_1859));
   MUX2_X1 i_8_0_1658 (.A(n_8_0_1861), .B(in_data[20]), .S(n_8_0_4065), .Z(
      n_8_0_1860));
   OAI21_X1 i_8_0_1659 (.A(n_8_0_1862), .B1(n_8_0_4070), .B2(n_8_0_6994), 
      .ZN(n_8_0_1861));
   NAND2_X1 i_8_0_1660 (.A1(in_data[28]), .A2(n_8_0_4070), .ZN(n_8_0_1862));
   OAI22_X1 i_8_0_1661 (.A1(n_8_0_1864), .A2(n_8_0_1863), .B1(n_8_0_6988), 
      .B2(n_8_0_4079), .ZN(n_36));
   OAI21_X1 i_8_0_1662 (.A(n_8_0_4079), .B1(n_8_0_4082), .B2(in_data[4]), 
      .ZN(n_8_0_1863));
   AOI211_X1 i_8_0_1663 (.A(n_8_0_4083), .B(n_8_0_1865), .C1(n_8_0_1866), 
      .C2(n_8_0_4100), .ZN(n_8_0_1864));
   NOR2_X1 i_8_0_1664 (.A1(n_8_0_6990), .A2(n_8_0_4100), .ZN(n_8_0_1865));
   MUX2_X1 i_8_0_1665 (.A(in_data[12]), .B(n_8_0_1867), .S(n_8_0_4096), .Z(
      n_8_0_1866));
   OAI21_X1 i_8_0_1666 (.A(n_8_0_1868), .B1(n_8_0_1869), .B2(n_8_0_4090), 
      .ZN(n_8_0_1867));
   NAND2_X1 i_8_0_1667 (.A1(n_8_0_4090), .A2(in_data[16]), .ZN(n_8_0_1868));
   OAI21_X1 i_8_0_1668 (.A(n_8_0_1870), .B1(n_8_0_1871), .B2(n_8_0_4093), 
      .ZN(n_8_0_1869));
   NAND2_X1 i_8_0_1669 (.A1(n_8_0_6993), .A2(n_8_0_4093), .ZN(n_8_0_1870));
   OAI21_X1 i_8_0_1670 (.A(n_8_0_1872), .B1(n_8_0_4086), .B2(n_8_0_6994), 
      .ZN(n_8_0_1871));
   NAND2_X1 i_8_0_1671 (.A1(in_data[28]), .A2(n_8_0_4086), .ZN(n_8_0_1872));
   OAI21_X1 i_8_0_1674 (.A(n_8_0_4117), .B1(n_8_0_1875), .B2(n_8_0_4120), 
      .ZN(n_8_0_1874));
   OAI21_X1 i_8_0_1675 (.A(n_8_0_1876), .B1(n_8_0_4134), .B2(n_8_0_6991), 
      .ZN(n_8_0_1875));
   OAI211_X1 i_8_0_1676 (.A(n_8_0_4134), .B(n_8_0_1877), .C1(n_8_0_1878), 
      .C2(n_8_0_4119), .ZN(n_8_0_1876));
   NAND2_X1 i_8_0_1677 (.A1(n_8_0_6992), .A2(n_8_0_4119), .ZN(n_8_0_1877));
   OAI21_X1 i_8_0_1678 (.A(n_8_0_1879), .B1(n_8_0_1880), .B2(n_8_0_4123), 
      .ZN(n_8_0_1878));
   NAND2_X1 i_8_0_1679 (.A1(n_8_0_4123), .A2(in_data[20]), .ZN(n_8_0_1879));
   OAI21_X1 i_8_0_1680 (.A(n_8_0_1881), .B1(n_8_0_4129), .B2(in_data[24]), 
      .ZN(n_8_0_1880));
   NAND2_X1 i_8_0_1681 (.A1(n_8_0_4129), .A2(n_8_0_6995), .ZN(n_8_0_1881));
   NOR2_X1 i_8_0_1682 (.A1(n_8_0_4121), .A2(in_data[8]), .ZN(n_8_0_1882));
   AOI211_X1 i_8_0_1686 (.A(n_8_0_4150), .B(n_8_0_1886), .C1(n_8_0_1887), 
      .C2(n_8_0_4142), .ZN(n_8_0_1885));
   NOR2_X1 i_8_0_1687 (.A1(in_data[12]), .A2(n_8_0_4142), .ZN(n_8_0_1886));
   INV_X1 i_8_0_1688 (.A(n_8_0_1888), .ZN(n_8_0_1887));
   AOI21_X1 i_8_0_1689 (.A(n_8_0_1889), .B1(n_8_0_1890), .B2(n_8_0_4145), 
      .ZN(n_8_0_1888));
   NOR2_X1 i_8_0_1690 (.A1(in_data[16]), .A2(n_8_0_4145), .ZN(n_8_0_1889));
   OAI22_X1 i_8_0_1691 (.A1(n_8_0_1891), .A2(n_8_0_1892), .B1(n_8_0_4139), 
      .B2(in_data[20]), .ZN(n_8_0_1890));
   OAI21_X1 i_8_0_1692 (.A(n_8_0_4139), .B1(n_8_0_4153), .B2(n_8_0_6995), 
      .ZN(n_8_0_1891));
   AND2_X1 i_8_0_1693 (.A1(n_8_0_4153), .A2(in_data[24]), .ZN(n_8_0_1892));
   OAI21_X1 i_8_0_1694 (.A(n_8_0_1893), .B1(n_8_0_4184), .B2(n_8_0_6988), 
      .ZN(n_37));
   OAI211_X1 i_8_0_1695 (.A(n_8_0_1894), .B(n_8_0_4184), .C1(n_8_0_4187), 
      .C2(in_data[4]), .ZN(n_8_0_1893));
   OAI211_X1 i_8_0_1696 (.A(n_8_0_4187), .B(n_8_0_1895), .C1(n_8_0_1896), 
      .C2(n_8_0_4175), .ZN(n_8_0_1894));
   NAND2_X1 i_8_0_1697 (.A1(n_8_0_4175), .A2(in_data[8]), .ZN(n_8_0_1895));
   INV_X1 i_8_0_1698 (.A(n_8_0_1897), .ZN(n_8_0_1896));
   OAI21_X1 i_8_0_1699 (.A(n_8_0_1898), .B1(n_8_0_4178), .B2(n_8_0_6991), 
      .ZN(n_8_0_1897));
   NAND2_X1 i_8_0_1700 (.A1(n_8_0_1899), .A2(n_8_0_4178), .ZN(n_8_0_1898));
   OAI21_X1 i_8_0_1701 (.A(n_8_0_1900), .B1(n_8_0_4181), .B2(n_8_0_6992), 
      .ZN(n_8_0_1899));
   NAND2_X1 i_8_0_1702 (.A1(n_8_0_1901), .A2(n_8_0_4181), .ZN(n_8_0_1900));
   OAI21_X1 i_8_0_1703 (.A(n_8_0_1902), .B1(n_8_0_4169), .B2(n_8_0_6993), 
      .ZN(n_8_0_1901));
   OAI211_X1 i_8_0_1704 (.A(n_8_0_4169), .B(n_8_0_1903), .C1(n_8_0_4166), 
      .C2(in_data[24]), .ZN(n_8_0_1902));
   NAND2_X1 i_8_0_1705 (.A1(n_8_0_4166), .A2(n_8_0_6995), .ZN(n_8_0_1903));
   NAND2_X1 i_8_0_1709 (.A1(n_8_0_4204), .A2(in_data[8]), .ZN(n_8_0_1906));
   INV_X1 i_8_0_1710 (.A(n_8_0_1908), .ZN(n_8_0_1907));
   AOI22_X1 i_8_0_1711 (.A1(n_8_0_1909), .A2(n_8_0_1910), .B1(n_8_0_4214), 
      .B2(n_8_0_6991), .ZN(n_8_0_1908));
   AOI21_X1 i_8_0_1712 (.A(n_8_0_4214), .B1(n_8_0_4208), .B2(n_8_0_1911), 
      .ZN(n_8_0_1909));
   NAND2_X1 i_8_0_1713 (.A1(n_8_0_4209), .A2(in_data[16]), .ZN(n_8_0_1910));
   OAI21_X1 i_8_0_1714 (.A(n_8_0_1912), .B1(n_8_0_4193), .B2(n_8_0_6993), 
      .ZN(n_8_0_1911));
   OAI211_X1 i_8_0_1715 (.A(n_8_0_4193), .B(n_8_0_1913), .C1(in_data[24]), 
      .C2(n_8_0_4196), .ZN(n_8_0_1912));
   NAND2_X1 i_8_0_1716 (.A1(n_8_0_4196), .A2(n_8_0_6995), .ZN(n_8_0_1913));
   OAI21_X1 i_8_0_1717 (.A(n_8_0_1914), .B1(n_8_0_4233), .B2(n_8_0_6988), 
      .ZN(n_38));
   NAND3_X1 i_8_0_1718 (.A1(n_8_0_1916), .A2(n_8_0_1915), .A3(n_8_0_4233), 
      .ZN(n_8_0_1914));
   NAND2_X1 i_8_0_1719 (.A1(n_8_0_6989), .A2(n_8_0_4236), .ZN(n_8_0_1915));
   OAI21_X1 i_8_0_1720 (.A(n_8_0_1917), .B1(n_8_0_1918), .B2(n_8_0_4223), 
      .ZN(n_8_0_1916));
   AOI21_X1 i_8_0_1721 (.A(n_8_0_4236), .B1(n_8_0_4223), .B2(in_data[8]), 
      .ZN(n_8_0_1917));
   INV_X1 i_8_0_1722 (.A(n_8_0_1919), .ZN(n_8_0_1918));
   MUX2_X1 i_8_0_1723 (.A(n_8_0_1920), .B(in_data[12]), .S(n_8_0_4241), .Z(
      n_8_0_1919));
   MUX2_X1 i_8_0_1724 (.A(n_8_0_1921), .B(in_data[16]), .S(n_8_0_4239), .Z(
      n_8_0_1920));
   AOI21_X1 i_8_0_1725 (.A(n_8_0_1922), .B1(n_8_0_4243), .B2(n_8_0_6993), 
      .ZN(n_8_0_1921));
   AOI211_X1 i_8_0_1726 (.A(n_8_0_4243), .B(n_8_0_1923), .C1(n_8_0_4226), 
      .C2(in_data[24]), .ZN(n_8_0_1922));
   NOR2_X1 i_8_0_1727 (.A1(n_8_0_6995), .A2(n_8_0_4226), .ZN(n_8_0_1923));
   OAI21_X1 i_8_0_1728 (.A(n_8_0_1924), .B1(n_8_0_4257), .B2(n_8_0_6988), 
      .ZN(n_39));
   NAND2_X1 i_8_0_1729 (.A1(n_8_0_4257), .A2(n_8_0_1925), .ZN(n_8_0_1924));
   AOI21_X1 i_8_0_1730 (.A(n_8_0_1926), .B1(n_8_0_4252), .B2(n_8_0_6989), 
      .ZN(n_8_0_1925));
   AOI211_X1 i_8_0_1731 (.A(n_8_0_4252), .B(n_8_0_1927), .C1(n_8_0_4250), 
      .C2(in_data[8]), .ZN(n_8_0_1926));
   AOI221_X1 i_8_0_1732 (.A(n_8_0_4250), .B1(n_8_0_4247), .B2(n_8_0_6991), 
      .C1(n_8_0_1929), .C2(n_8_0_1928), .ZN(n_8_0_1927));
   AOI21_X1 i_8_0_1733 (.A(n_8_0_4247), .B1(n_8_0_4273), .B2(in_data[16]), 
      .ZN(n_8_0_1928));
   NAND2_X1 i_8_0_1734 (.A1(n_8_0_1930), .A2(n_8_0_4272), .ZN(n_8_0_1929));
   OAI22_X1 i_8_0_1735 (.A1(n_8_0_1931), .A2(n_8_0_1932), .B1(n_8_0_4260), 
      .B2(n_8_0_6993), .ZN(n_8_0_1930));
   OAI21_X1 i_8_0_1736 (.A(n_8_0_4260), .B1(n_8_0_4269), .B2(in_data[28]), 
      .ZN(n_8_0_1931));
   AND2_X1 i_8_0_1737 (.A1(n_8_0_6994), .A2(n_8_0_4269), .ZN(n_8_0_1932));
   OAI22_X1 i_8_0_1738 (.A1(n_8_0_1934), .A2(n_8_0_1933), .B1(n_8_0_6988), 
      .B2(n_8_0_4290), .ZN(n_40));
   OAI21_X1 i_8_0_1739 (.A(n_8_0_4290), .B1(n_8_0_4298), .B2(in_data[4]), 
      .ZN(n_8_0_1933));
   NOR2_X1 i_8_0_1740 (.A1(n_8_0_1936), .A2(n_8_0_1935), .ZN(n_8_0_1934));
   OAI21_X1 i_8_0_1741 (.A(n_8_0_4298), .B1(n_8_0_4279), .B2(n_8_0_6990), 
      .ZN(n_8_0_1935));
   AOI21_X1 i_8_0_1742 (.A(n_8_0_1937), .B1(n_8_0_1938), .B2(n_8_0_4295), 
      .ZN(n_8_0_1936));
   OAI21_X1 i_8_0_1743 (.A(n_8_0_4279), .B1(n_8_0_4295), .B2(in_data[12]), 
      .ZN(n_8_0_1937));
   INV_X1 i_8_0_1744 (.A(n_8_0_1939), .ZN(n_8_0_1938));
   AOI21_X1 i_8_0_1745 (.A(n_8_0_1940), .B1(n_8_0_4292), .B2(n_8_0_6992), 
      .ZN(n_8_0_1939));
   AOI211_X1 i_8_0_1746 (.A(n_8_0_4292), .B(n_8_0_1941), .C1(n_8_0_1942), 
      .C2(n_8_0_4287), .ZN(n_8_0_1940));
   NOR2_X1 i_8_0_1747 (.A1(n_8_0_4287), .A2(n_8_0_6993), .ZN(n_8_0_1941));
   AOI21_X1 i_8_0_1748 (.A(n_8_0_1943), .B1(n_8_0_4282), .B2(n_8_0_6995), 
      .ZN(n_8_0_1942));
   NOR2_X1 i_8_0_1749 (.A1(in_data[24]), .A2(n_8_0_4282), .ZN(n_8_0_1943));
   AOI211_X1 i_8_0_1754 (.A(n_8_0_4328), .B(n_8_0_1949), .C1(n_8_0_4303), 
      .C2(in_data[16]), .ZN(n_8_0_1947));
   OAI21_X1 i_8_0_1755 (.A(n_8_0_4314), .B1(n_8_0_4327), .B2(in_data[12]), 
      .ZN(n_8_0_1948));
   AOI211_X1 i_8_0_1756 (.A(n_8_0_4303), .B(n_8_0_1950), .C1(n_8_0_6993), 
      .C2(n_8_0_4330), .ZN(n_8_0_1949));
   AOI211_X1 i_8_0_1757 (.A(n_8_0_1951), .B(n_8_0_4330), .C1(in_data[28]), 
      .C2(n_8_0_4320), .ZN(n_8_0_1950));
   NOR2_X1 i_8_0_1758 (.A1(n_8_0_4320), .A2(n_8_0_6994), .ZN(n_8_0_1951));
   MUX2_X1 i_8_0_1759 (.A(n_8_0_1952), .B(in_data[0]), .S(n_8_0_4336), .Z(n_41));
   AOI22_X1 i_8_0_1760 (.A1(n_8_0_1954), .A2(n_8_0_1953), .B1(n_8_0_6989), 
      .B2(n_8_0_4345), .ZN(n_8_0_1952));
   AOI21_X1 i_8_0_1761 (.A(n_8_0_4345), .B1(n_8_0_4352), .B2(in_data[8]), 
      .ZN(n_8_0_1953));
   NAND3_X1 i_8_0_1762 (.A1(n_8_0_4351), .A2(n_8_0_1956), .A3(n_8_0_1955), 
      .ZN(n_8_0_1954));
   NAND2_X1 i_8_0_1763 (.A1(n_8_0_6991), .A2(n_8_0_4337), .ZN(n_8_0_1955));
   OAI21_X1 i_8_0_1764 (.A(n_8_0_1957), .B1(n_8_0_1958), .B2(n_8_0_4339), 
      .ZN(n_8_0_1956));
   AOI21_X1 i_8_0_1765 (.A(n_8_0_4337), .B1(n_8_0_4339), .B2(in_data[16]), 
      .ZN(n_8_0_1957));
   AOI21_X1 i_8_0_1766 (.A(n_8_0_1959), .B1(n_8_0_1960), .B2(n_8_0_4353), 
      .ZN(n_8_0_1958));
   NOR2_X1 i_8_0_1767 (.A1(n_8_0_4353), .A2(n_8_0_6993), .ZN(n_8_0_1959));
   OAI21_X1 i_8_0_1768 (.A(n_8_0_1961), .B1(n_8_0_4342), .B2(n_8_0_6995), 
      .ZN(n_8_0_1960));
   NAND2_X1 i_8_0_1769 (.A1(n_8_0_4342), .A2(in_data[24]), .ZN(n_8_0_1961));
   OAI21_X1 i_8_0_1770 (.A(n_8_0_1962), .B1(n_8_0_1963), .B2(n_8_0_4370), 
      .ZN(n_42));
   NAND2_X1 i_8_0_1771 (.A1(n_8_0_4370), .A2(in_data[0]), .ZN(n_8_0_1962));
   OAI21_X1 i_8_0_1772 (.A(n_8_0_1964), .B1(n_8_0_4373), .B2(in_data[4]), 
      .ZN(n_8_0_1963));
   OAI211_X1 i_8_0_1773 (.A(n_8_0_4373), .B(n_8_0_1965), .C1(n_8_0_1966), 
      .C2(n_8_0_4375), .ZN(n_8_0_1964));
   NAND2_X1 i_8_0_1774 (.A1(n_8_0_4375), .A2(in_data[8]), .ZN(n_8_0_1965));
   INV_X1 i_8_0_1775 (.A(n_8_0_1967), .ZN(n_8_0_1966));
   MUX2_X1 i_8_0_1776 (.A(n_8_0_1968), .B(in_data[12]), .S(n_8_0_4380), .Z(
      n_8_0_1967));
   MUX2_X1 i_8_0_1777 (.A(n_8_0_1969), .B(in_data[16]), .S(n_8_0_4386), .Z(
      n_8_0_1968));
   MUX2_X1 i_8_0_1778 (.A(n_8_0_1970), .B(in_data[20]), .S(n_8_0_4363), .Z(
      n_8_0_1969));
   OAI21_X1 i_8_0_1779 (.A(n_8_0_1971), .B1(n_8_0_4359), .B2(n_8_0_6995), 
      .ZN(n_8_0_1970));
   NAND2_X1 i_8_0_1780 (.A1(n_8_0_4359), .A2(in_data[24]), .ZN(n_8_0_1971));
   NOR2_X1 i_8_0_1784 (.A1(n_8_0_1975), .A2(n_8_0_4401), .ZN(n_8_0_1974));
   AOI21_X1 i_8_0_1785 (.A(n_8_0_1976), .B1(n_8_0_1977), .B2(n_8_0_4393), 
      .ZN(n_8_0_1975));
   NOR2_X1 i_8_0_1786 (.A1(n_8_0_6991), .A2(n_8_0_4393), .ZN(n_8_0_1976));
   OAI21_X1 i_8_0_1787 (.A(n_8_0_1978), .B1(n_8_0_4411), .B2(n_8_0_6992), 
      .ZN(n_8_0_1977));
   OAI211_X1 i_8_0_1788 (.A(n_8_0_1979), .B(n_8_0_4411), .C1(in_data[20]), 
      .C2(n_8_0_4390), .ZN(n_8_0_1978));
   OAI211_X1 i_8_0_1789 (.A(n_8_0_4390), .B(n_8_0_1980), .C1(n_8_0_6995), 
      .C2(n_8_0_4399), .ZN(n_8_0_1979));
   NAND2_X1 i_8_0_1790 (.A1(n_8_0_4399), .A2(in_data[24]), .ZN(n_8_0_1980));
   INV_X1 i_8_0_1791 (.A(n_8_0_1981), .ZN(n_43));
   AOI21_X1 i_8_0_1792 (.A(n_8_0_1982), .B1(n_8_0_4421), .B2(in_data[0]), 
      .ZN(n_8_0_1981));
   AOI211_X1 i_8_0_1793 (.A(n_8_0_4421), .B(n_8_0_1983), .C1(n_8_0_1984), 
      .C2(n_8_0_4418), .ZN(n_8_0_1982));
   NOR2_X1 i_8_0_1794 (.A1(in_data[4]), .A2(n_8_0_4418), .ZN(n_8_0_1983));
   INV_X1 i_8_0_1795 (.A(n_8_0_1985), .ZN(n_8_0_1984));
   OAI22_X1 i_8_0_1796 (.A1(n_8_0_1987), .A2(n_8_0_1986), .B1(n_8_0_6990), 
      .B2(n_8_0_4434), .ZN(n_8_0_1985));
   OAI21_X1 i_8_0_1797 (.A(n_8_0_4434), .B1(n_8_0_4432), .B2(in_data[12]), 
      .ZN(n_8_0_1986));
   AOI221_X1 i_8_0_1798 (.A(n_8_0_4431), .B1(n_8_0_1989), .B2(n_8_0_1988), 
      .C1(n_8_0_4428), .C2(in_data[16]), .ZN(n_8_0_1987));
   AOI21_X1 i_8_0_1799 (.A(n_8_0_4428), .B1(n_8_0_4437), .B2(n_8_0_6993), 
      .ZN(n_8_0_1988));
   OAI21_X1 i_8_0_1800 (.A(n_8_0_1990), .B1(n_8_0_4440), .B2(n_8_0_6994), 
      .ZN(n_8_0_1989));
   AOI21_X1 i_8_0_1801 (.A(n_8_0_4437), .B1(n_8_0_4440), .B2(in_data[28]), 
      .ZN(n_8_0_1990));
   MUX2_X1 i_8_0_1802 (.A(n_8_0_1991), .B(in_data[0]), .S(n_8_0_4468), .Z(n_44));
   AOI22_X1 i_8_0_1803 (.A1(n_8_0_1993), .A2(n_8_0_1992), .B1(n_8_0_6989), 
      .B2(n_8_0_4455), .ZN(n_8_0_1991));
   AOI21_X1 i_8_0_1804 (.A(n_8_0_4455), .B1(n_8_0_4445), .B2(in_data[8]), 
      .ZN(n_8_0_1992));
   OAI21_X1 i_8_0_1805 (.A(n_8_0_1994), .B1(n_8_0_1995), .B2(n_8_0_4448), 
      .ZN(n_8_0_1993));
   AOI21_X1 i_8_0_1806 (.A(n_8_0_4445), .B1(n_8_0_4448), .B2(n_8_0_6991), 
      .ZN(n_8_0_1994));
   AOI21_X1 i_8_0_1807 (.A(n_8_0_1996), .B1(n_8_0_4471), .B2(n_8_0_6992), 
      .ZN(n_8_0_1995));
   NOR2_X1 i_8_0_1808 (.A1(n_8_0_1997), .A2(n_8_0_4471), .ZN(n_8_0_1996));
   AOI21_X1 i_8_0_1809 (.A(n_8_0_1998), .B1(n_8_0_1999), .B2(n_8_0_4461), 
      .ZN(n_8_0_1997));
   NOR2_X1 i_8_0_1810 (.A1(in_data[20]), .A2(n_8_0_4461), .ZN(n_8_0_1998));
   OAI21_X1 i_8_0_1811 (.A(n_8_0_2000), .B1(n_8_0_4465), .B2(in_data[28]), 
      .ZN(n_8_0_1999));
   NAND2_X1 i_8_0_1812 (.A1(n_8_0_6994), .A2(n_8_0_4465), .ZN(n_8_0_2000));
   OAI21_X1 i_8_0_1813 (.A(n_8_0_2001), .B1(n_8_0_4501), .B2(n_8_0_6988), 
      .ZN(n_45));
   NAND2_X1 i_8_0_1814 (.A1(n_8_0_4501), .A2(n_8_0_2002), .ZN(n_8_0_2001));
   MUX2_X1 i_8_0_1815 (.A(in_data[4]), .B(n_8_0_2003), .S(n_8_0_4504), .Z(
      n_8_0_2002));
   MUX2_X1 i_8_0_1816 (.A(n_8_0_2004), .B(in_data[8]), .S(n_8_0_4488), .Z(
      n_8_0_2003));
   MUX2_X1 i_8_0_1817 (.A(in_data[12]), .B(n_8_0_2005), .S(n_8_0_4481), .Z(
      n_8_0_2004));
   AOI21_X1 i_8_0_1818 (.A(n_8_0_2006), .B1(n_8_0_4491), .B2(n_8_0_6992), 
      .ZN(n_8_0_2005));
   NOR2_X1 i_8_0_1819 (.A1(n_8_0_2007), .A2(n_8_0_4491), .ZN(n_8_0_2006));
   AOI21_X1 i_8_0_1820 (.A(n_8_0_2008), .B1(n_8_0_2009), .B2(n_8_0_4495), 
      .ZN(n_8_0_2007));
   NOR2_X1 i_8_0_1821 (.A1(in_data[20]), .A2(n_8_0_4495), .ZN(n_8_0_2008));
   OAI21_X1 i_8_0_1822 (.A(n_8_0_2010), .B1(n_8_0_4478), .B2(in_data[28]), 
      .ZN(n_8_0_2009));
   NAND2_X1 i_8_0_1823 (.A1(n_8_0_6994), .A2(n_8_0_4478), .ZN(n_8_0_2010));
   OAI21_X1 i_8_0_1824 (.A(n_8_0_2011), .B1(n_8_0_4527), .B2(n_8_0_6988), 
      .ZN(n_46));
   NAND2_X1 i_8_0_1825 (.A1(n_8_0_4527), .A2(n_8_0_2012), .ZN(n_8_0_2011));
   MUX2_X1 i_8_0_1826 (.A(in_data[4]), .B(n_8_0_2013), .S(n_8_0_4554), .Z(
      n_8_0_2012));
   MUX2_X1 i_8_0_1827 (.A(n_8_0_2014), .B(in_data[8]), .S(n_8_0_4546), .Z(
      n_8_0_2013));
   MUX2_X1 i_8_0_1828 (.A(in_data[12]), .B(n_8_0_2015), .S(n_8_0_4536), .Z(
      n_8_0_2014));
   AOI21_X1 i_8_0_1829 (.A(n_8_0_2016), .B1(n_8_0_2017), .B2(n_8_0_4533), 
      .ZN(n_8_0_2015));
   NOR2_X1 i_8_0_1830 (.A1(in_data[16]), .A2(n_8_0_4533), .ZN(n_8_0_2016));
   OAI21_X1 i_8_0_1831 (.A(n_8_0_2018), .B1(n_8_0_4516), .B2(in_data[20]), 
      .ZN(n_8_0_2017));
   NAND2_X1 i_8_0_1832 (.A1(n_8_0_4516), .A2(n_8_0_2019), .ZN(n_8_0_2018));
   OAI21_X1 i_8_0_1833 (.A(n_8_0_2020), .B1(n_8_0_4521), .B2(in_data[28]), 
      .ZN(n_8_0_2019));
   NAND2_X1 i_8_0_1834 (.A1(n_8_0_6994), .A2(n_8_0_4521), .ZN(n_8_0_2020));
   OAI21_X1 i_8_0_1835 (.A(n_8_0_2021), .B1(n_8_0_4594), .B2(n_8_0_6988), 
      .ZN(n_47));
   OAI211_X1 i_8_0_1836 (.A(n_8_0_4594), .B(n_8_0_2022), .C1(n_8_0_2025), 
      .C2(n_8_0_2023), .ZN(n_8_0_2021));
   NAND2_X1 i_8_0_1837 (.A1(n_8_0_6989), .A2(n_8_0_4609), .ZN(n_8_0_2022));
   INV_X1 i_8_0_1838 (.A(n_8_0_2024), .ZN(n_8_0_2023));
   AOI21_X1 i_8_0_1839 (.A(n_8_0_4609), .B1(n_8_0_4570), .B2(in_data[8]), 
      .ZN(n_8_0_2024));
   AOI211_X1 i_8_0_1840 (.A(n_8_0_4570), .B(n_8_0_2026), .C1(n_8_0_6991), 
      .C2(n_8_0_4607), .ZN(n_8_0_2025));
   NOR2_X1 i_8_0_1841 (.A1(n_8_0_4607), .A2(n_8_0_2027), .ZN(n_8_0_2026));
   AOI21_X1 i_8_0_1842 (.A(n_8_0_2028), .B1(n_8_0_4589), .B2(n_8_0_6992), 
      .ZN(n_8_0_2027));
   AOI211_X1 i_8_0_1843 (.A(n_8_0_4589), .B(n_8_0_2029), .C1(n_8_0_2030), 
      .C2(n_8_0_4583), .ZN(n_8_0_2028));
   NOR2_X1 i_8_0_1844 (.A1(n_8_0_4583), .A2(n_8_0_6993), .ZN(n_8_0_2029));
   OAI21_X1 i_8_0_1845 (.A(n_8_0_2031), .B1(n_8_0_4578), .B2(n_8_0_6995), 
      .ZN(n_8_0_2030));
   NAND2_X1 i_8_0_1846 (.A1(n_8_0_4578), .A2(in_data[24]), .ZN(n_8_0_2031));
   AOI21_X1 i_8_0_1847 (.A(n_8_0_2032), .B1(n_8_0_2042), .B2(n_8_0_6988), 
      .ZN(n_48));
   NOR2_X1 i_8_0_1848 (.A1(n_8_0_2042), .A2(n_8_0_2033), .ZN(n_8_0_2032));
   AOI22_X1 i_8_0_1849 (.A1(n_8_0_2035), .A2(n_8_0_2034), .B1(n_8_0_6989), 
      .B2(n_8_0_4625), .ZN(n_8_0_2033));
   AOI21_X1 i_8_0_1850 (.A(n_8_0_4625), .B1(n_8_0_4623), .B2(in_data[8]), 
      .ZN(n_8_0_2034));
   OAI21_X1 i_8_0_1851 (.A(n_8_0_2036), .B1(n_8_0_2037), .B2(n_8_0_4624), 
      .ZN(n_8_0_2035));
   AOI21_X1 i_8_0_1852 (.A(n_8_0_4623), .B1(n_8_0_4624), .B2(n_8_0_6991), 
      .ZN(n_8_0_2036));
   OAI21_X1 i_8_0_1853 (.A(n_8_0_2038), .B1(n_8_0_4619), .B2(n_8_0_6992), 
      .ZN(n_8_0_2037));
   OAI211_X1 i_8_0_1854 (.A(n_8_0_2039), .B(n_8_0_4619), .C1(n_8_0_4617), 
      .C2(n_8_0_2040), .ZN(n_8_0_2038));
   NAND2_X1 i_8_0_1855 (.A1(n_8_0_6993), .A2(n_8_0_4617), .ZN(n_8_0_2039));
   OAI21_X1 i_8_0_1856 (.A(n_8_0_2041), .B1(n_8_0_4618), .B2(n_8_0_6995), 
      .ZN(n_8_0_2040));
   NAND2_X1 i_8_0_1857 (.A1(n_8_0_4618), .A2(in_data[24]), .ZN(n_8_0_2041));
   AOI21_X1 i_8_0_1858 (.A(n_8_0_4597), .B1(n_8_0_6465), .B2(n_8_0_441), 
      .ZN(n_8_0_2042));
   OAI21_X1 i_8_0_1859 (.A(n_8_0_2043), .B1(n_8_0_2044), .B2(n_8_0_6988), 
      .ZN(n_49));
   OAI211_X1 i_8_0_1860 (.A(n_8_0_2045), .B(n_8_0_2044), .C1(in_data[4]), 
      .C2(n_8_0_4650), .ZN(n_8_0_2043));
   OAI21_X1 i_8_0_1861 (.A(n_8_0_4630), .B1(n_8_0_6729), .B2(n_8_0_4631), 
      .ZN(n_8_0_2044));
   OAI211_X1 i_8_0_1862 (.A(n_8_0_4650), .B(n_8_0_2046), .C1(n_8_0_2047), 
      .C2(n_8_0_4636), .ZN(n_8_0_2045));
   NAND2_X1 i_8_0_1863 (.A1(in_data[8]), .A2(n_8_0_4636), .ZN(n_8_0_2046));
   INV_X1 i_8_0_1864 (.A(n_8_0_2048), .ZN(n_8_0_2047));
   OAI21_X1 i_8_0_1865 (.A(n_8_0_2049), .B1(n_8_0_4647), .B2(n_8_0_6991), 
      .ZN(n_8_0_2048));
   NAND2_X1 i_8_0_1866 (.A1(n_8_0_4647), .A2(n_8_0_2050), .ZN(n_8_0_2049));
   MUX2_X1 i_8_0_1867 (.A(n_8_0_2051), .B(in_data[16]), .S(n_8_0_4644), .Z(
      n_8_0_2050));
   MUX2_X1 i_8_0_1868 (.A(n_8_0_2052), .B(in_data[20]), .S(n_8_0_4633), .Z(
      n_8_0_2051));
   OAI21_X1 i_8_0_1869 (.A(n_8_0_2053), .B1(n_8_0_4639), .B2(n_8_0_6994), 
      .ZN(n_8_0_2052));
   NAND2_X1 i_8_0_1870 (.A1(n_8_0_4639), .A2(in_data[28]), .ZN(n_8_0_2053));
   OAI22_X1 i_8_0_1871 (.A1(n_8_0_2056), .A2(n_8_0_2054), .B1(n_8_0_2055), 
      .B2(n_8_0_6988), .ZN(n_50));
   OAI21_X1 i_8_0_1872 (.A(n_8_0_2055), .B1(n_8_0_4674), .B2(in_data[4]), 
      .ZN(n_8_0_2054));
   AOI21_X1 i_8_0_1873 (.A(n_8_0_4658), .B1(n_8_0_4659), .B2(n_8_0_6729), 
      .ZN(n_8_0_2055));
   AOI21_X1 i_8_0_1874 (.A(n_8_0_2057), .B1(n_8_0_2058), .B2(n_8_0_4670), 
      .ZN(n_8_0_2056));
   OAI21_X1 i_8_0_1875 (.A(n_8_0_4674), .B1(n_8_0_4670), .B2(n_8_0_6990), 
      .ZN(n_8_0_2057));
   MUX2_X1 i_8_0_1876 (.A(n_8_0_2059), .B(in_data[12]), .S(n_8_0_4672), .Z(
      n_8_0_2058));
   OAI21_X1 i_8_0_1877 (.A(n_8_0_2060), .B1(n_8_0_2061), .B2(n_8_0_4667), 
      .ZN(n_8_0_2059));
   NAND2_X1 i_8_0_1878 (.A1(in_data[16]), .A2(n_8_0_4667), .ZN(n_8_0_2060));
   AOI21_X1 i_8_0_1879 (.A(n_8_0_2062), .B1(n_8_0_2063), .B2(n_8_0_4661), 
      .ZN(n_8_0_2061));
   NOR2_X1 i_8_0_1880 (.A1(n_8_0_6993), .A2(n_8_0_4661), .ZN(n_8_0_2062));
   AOI21_X1 i_8_0_1881 (.A(n_8_0_2064), .B1(n_8_0_4655), .B2(n_8_0_6994), 
      .ZN(n_8_0_2063));
   NOR2_X1 i_8_0_1882 (.A1(in_data[28]), .A2(n_8_0_4655), .ZN(n_8_0_2064));
   OAI22_X1 i_8_0_1883 (.A1(n_8_0_2066), .A2(n_8_0_2065), .B1(n_8_0_6988), 
      .B2(n_8_0_2075), .ZN(n_51));
   OAI21_X1 i_8_0_1884 (.A(n_8_0_2075), .B1(n_8_0_4701), .B2(in_data[4]), 
      .ZN(n_8_0_2065));
   AOI21_X1 i_8_0_1885 (.A(n_8_0_2067), .B1(n_8_0_2068), .B2(n_8_0_4698), 
      .ZN(n_8_0_2066));
   OAI21_X1 i_8_0_1886 (.A(n_8_0_4701), .B1(n_8_0_4698), .B2(n_8_0_6990), 
      .ZN(n_8_0_2067));
   OAI22_X1 i_8_0_1887 (.A1(n_8_0_2070), .A2(n_8_0_2069), .B1(n_8_0_6991), 
      .B2(n_8_0_4695), .ZN(n_8_0_2068));
   OAI21_X1 i_8_0_1888 (.A(n_8_0_4695), .B1(n_8_0_4688), .B2(in_data[16]), 
      .ZN(n_8_0_2069));
   AOI21_X1 i_8_0_1889 (.A(n_8_0_2071), .B1(n_8_0_4692), .B2(in_data[20]), 
      .ZN(n_8_0_2070));
   OAI21_X1 i_8_0_1890 (.A(n_8_0_4688), .B1(n_8_0_2072), .B2(n_8_0_4692), 
      .ZN(n_8_0_2071));
   INV_X1 i_8_0_1891 (.A(n_8_0_2073), .ZN(n_8_0_2072));
   OAI21_X1 i_8_0_1892 (.A(n_8_0_2074), .B1(n_8_0_4683), .B2(n_8_0_6994), 
      .ZN(n_8_0_2073));
   NAND2_X1 i_8_0_1893 (.A1(n_8_0_4683), .A2(in_data[28]), .ZN(n_8_0_2074));
   AOI21_X1 i_8_0_1894 (.A(n_8_0_2076), .B1(n_8_0_6729), .B2(n_8_0_6875), 
      .ZN(n_8_0_2075));
   AOI21_X1 i_8_0_1895 (.A(n_8_0_4686), .B1(n_8_0_6730), .B2(n_8_0_444), 
      .ZN(n_8_0_2076));
   OAI21_X1 i_8_0_1896 (.A(n_8_0_2077), .B1(n_8_0_4714), .B2(n_8_0_6988), 
      .ZN(n_52));
   OAI211_X1 i_8_0_1897 (.A(n_8_0_4714), .B(n_8_0_2078), .C1(n_8_0_2079), 
      .C2(n_8_0_4726), .ZN(n_8_0_2077));
   NAND2_X1 i_8_0_1898 (.A1(n_8_0_4726), .A2(n_8_0_6989), .ZN(n_8_0_2078));
   MUX2_X1 i_8_0_1899 (.A(n_8_0_2080), .B(in_data[8]), .S(n_8_0_4717), .Z(
      n_8_0_2079));
   AOI21_X1 i_8_0_1900 (.A(n_8_0_2081), .B1(n_8_0_4720), .B2(n_8_0_6991), 
      .ZN(n_8_0_2080));
   AOI211_X1 i_8_0_1901 (.A(n_8_0_4720), .B(n_8_0_2082), .C1(n_8_0_2083), 
      .C2(n_8_0_4706), .ZN(n_8_0_2081));
   NOR2_X1 i_8_0_1902 (.A1(n_8_0_6992), .A2(n_8_0_4706), .ZN(n_8_0_2082));
   AOI21_X1 i_8_0_1903 (.A(n_8_0_2084), .B1(n_8_0_2085), .B2(n_8_0_4723), 
      .ZN(n_8_0_2083));
   NOR2_X1 i_8_0_1904 (.A1(n_8_0_4723), .A2(in_data[20]), .ZN(n_8_0_2084));
   OAI21_X1 i_8_0_1905 (.A(n_8_0_2086), .B1(n_8_0_4711), .B2(in_data[24]), 
      .ZN(n_8_0_2085));
   NAND2_X1 i_8_0_1906 (.A1(n_8_0_6995), .A2(n_8_0_4711), .ZN(n_8_0_2086));
   OAI22_X1 i_8_0_1907 (.A1(n_8_0_2088), .A2(n_8_0_2087), .B1(n_8_0_6988), 
      .B2(n_8_0_2096), .ZN(n_53));
   OAI21_X1 i_8_0_1908 (.A(n_8_0_2096), .B1(n_8_0_4757), .B2(in_data[4]), 
      .ZN(n_8_0_2087));
   AOI211_X1 i_8_0_1909 (.A(n_8_0_4756), .B(n_8_0_2089), .C1(n_8_0_4753), 
      .C2(in_data[8]), .ZN(n_8_0_2088));
   AOI211_X1 i_8_0_1910 (.A(n_8_0_4753), .B(n_8_0_2090), .C1(n_8_0_2091), 
      .C2(n_8_0_4750), .ZN(n_8_0_2089));
   NOR2_X1 i_8_0_1911 (.A1(n_8_0_4750), .A2(in_data[12]), .ZN(n_8_0_2090));
   INV_X1 i_8_0_1912 (.A(n_8_0_2092), .ZN(n_8_0_2091));
   OAI21_X1 i_8_0_1913 (.A(n_8_0_2093), .B1(n_8_0_4747), .B2(n_8_0_6992), 
      .ZN(n_8_0_2092));
   OAI211_X1 i_8_0_1914 (.A(n_8_0_4747), .B(n_8_0_2094), .C1(n_8_0_4738), 
      .C2(in_data[20]), .ZN(n_8_0_2093));
   OAI211_X1 i_8_0_1915 (.A(n_8_0_4738), .B(n_8_0_2095), .C1(n_8_0_6994), 
      .C2(n_8_0_4741), .ZN(n_8_0_2094));
   NAND2_X1 i_8_0_1916 (.A1(n_8_0_4741), .A2(in_data[28]), .ZN(n_8_0_2095));
   OAI21_X1 i_8_0_1917 (.A(n_8_0_4744), .B1(n_8_0_6729), .B2(n_8_0_4745), 
      .ZN(n_8_0_2096));
   AOI22_X1 i_8_0_1918 (.A1(n_8_0_2097), .A2(n_8_0_2099), .B1(n_8_0_6988), 
      .B2(n_8_0_2098), .ZN(n_54));
   AOI21_X1 i_8_0_1919 (.A(n_8_0_2098), .B1(n_8_0_4781), .B2(in_data[4]), 
      .ZN(n_8_0_2097));
   OAI21_X1 i_8_0_1920 (.A(n_8_0_4768), .B1(n_8_0_4769), .B2(n_8_0_6730), 
      .ZN(n_8_0_2098));
   OAI21_X1 i_8_0_1921 (.A(n_8_0_2100), .B1(n_8_0_2101), .B2(n_8_0_4784), 
      .ZN(n_8_0_2099));
   AOI21_X1 i_8_0_1922 (.A(n_8_0_4781), .B1(n_8_0_4784), .B2(n_8_0_6990), 
      .ZN(n_8_0_2100));
   AOI21_X1 i_8_0_1923 (.A(n_8_0_2107), .B1(n_8_0_2102), .B2(n_8_0_4779), 
      .ZN(n_8_0_2101));
   OAI21_X1 i_8_0_1924 (.A(n_8_0_2103), .B1(n_8_0_4774), .B2(in_data[16]), 
      .ZN(n_8_0_2102));
   OAI211_X1 i_8_0_1925 (.A(n_8_0_4774), .B(n_8_0_2104), .C1(n_8_0_2105), 
      .C2(n_8_0_4763), .ZN(n_8_0_2103));
   NAND2_X1 i_8_0_1926 (.A1(in_data[20]), .A2(n_8_0_4763), .ZN(n_8_0_2104));
   OAI21_X1 i_8_0_1927 (.A(n_8_0_2106), .B1(n_8_0_4771), .B2(in_data[24]), 
      .ZN(n_8_0_2105));
   NAND2_X1 i_8_0_1928 (.A1(n_8_0_6995), .A2(n_8_0_4771), .ZN(n_8_0_2106));
   NOR2_X1 i_8_0_1929 (.A1(n_8_0_4779), .A2(in_data[12]), .ZN(n_8_0_2107));
   OAI22_X1 i_8_0_1930 (.A1(n_8_0_2109), .A2(n_8_0_2108), .B1(n_8_0_6988), 
      .B2(n_8_0_2118), .ZN(n_55));
   OAI21_X1 i_8_0_1931 (.A(n_8_0_2118), .B1(n_8_0_4790), .B2(in_data[4]), 
      .ZN(n_8_0_2108));
   AOI21_X1 i_8_0_1932 (.A(n_8_0_2110), .B1(n_8_0_2111), .B2(n_8_0_4811), 
      .ZN(n_8_0_2109));
   OAI21_X1 i_8_0_1933 (.A(n_8_0_4790), .B1(n_8_0_4811), .B2(n_8_0_6990), 
      .ZN(n_8_0_2110));
   MUX2_X1 i_8_0_1934 (.A(n_8_0_2112), .B(in_data[12]), .S(n_8_0_4808), .Z(
      n_8_0_2111));
   OAI21_X1 i_8_0_1935 (.A(n_8_0_2113), .B1(n_8_0_2114), .B2(n_8_0_4796), 
      .ZN(n_8_0_2112));
   NAND2_X1 i_8_0_1936 (.A1(in_data[16]), .A2(n_8_0_4796), .ZN(n_8_0_2113));
   OAI21_X1 i_8_0_1937 (.A(n_8_0_2115), .B1(n_8_0_2116), .B2(n_8_0_4799), 
      .ZN(n_8_0_2114));
   NAND2_X1 i_8_0_1938 (.A1(n_8_0_4799), .A2(n_8_0_6993), .ZN(n_8_0_2115));
   OAI21_X1 i_8_0_1939 (.A(n_8_0_2117), .B1(n_8_0_4805), .B2(n_8_0_6994), 
      .ZN(n_8_0_2116));
   NAND2_X1 i_8_0_1940 (.A1(n_8_0_4805), .A2(in_data[28]), .ZN(n_8_0_2117));
   OAI21_X1 i_8_0_1941 (.A(n_8_0_4802), .B1(n_8_0_6729), .B2(n_8_0_4803), 
      .ZN(n_8_0_2118));
   OAI21_X1 i_8_0_1942 (.A(n_8_0_2119), .B1(n_8_0_4820), .B2(n_8_0_6988), 
      .ZN(n_56));
   NAND2_X1 i_8_0_1943 (.A1(n_8_0_2120), .A2(n_8_0_4820), .ZN(n_8_0_2119));
   MUX2_X1 i_8_0_1944 (.A(n_8_0_2121), .B(in_data[4]), .S(n_8_0_4824), .Z(
      n_8_0_2120));
   OAI21_X1 i_8_0_1945 (.A(n_8_0_2122), .B1(n_8_0_4816), .B2(n_8_0_6990), 
      .ZN(n_8_0_2121));
   NAND2_X1 i_8_0_1946 (.A1(n_8_0_4816), .A2(n_8_0_2123), .ZN(n_8_0_2122));
   MUX2_X1 i_8_0_1947 (.A(n_8_0_2124), .B(in_data[12]), .S(n_8_0_4842), .Z(
      n_8_0_2123));
   OAI21_X1 i_8_0_1948 (.A(n_8_0_2128), .B1(n_8_0_2125), .B2(n_8_0_4827), 
      .ZN(n_8_0_2124));
   OAI22_X1 i_8_0_1949 (.A1(n_8_0_2126), .A2(n_8_0_2127), .B1(n_8_0_4832), 
      .B2(in_data[20]), .ZN(n_8_0_2125));
   OAI21_X1 i_8_0_1950 (.A(n_8_0_4832), .B1(n_8_0_4837), .B2(n_8_0_6995), 
      .ZN(n_8_0_2126));
   AND2_X1 i_8_0_1951 (.A1(in_data[24]), .A2(n_8_0_4837), .ZN(n_8_0_2127));
   NAND2_X1 i_8_0_1952 (.A1(n_8_0_4827), .A2(in_data[16]), .ZN(n_8_0_2128));
   AOI21_X1 i_8_0_1953 (.A(n_8_0_2129), .B1(n_8_0_4848), .B2(n_8_0_6988), 
      .ZN(n_57));
   NOR2_X1 i_8_0_1954 (.A1(n_8_0_4848), .A2(n_8_0_2130), .ZN(n_8_0_2129));
   AOI22_X1 i_8_0_1955 (.A1(n_8_0_2131), .A2(n_8_0_2132), .B1(n_8_0_4857), 
      .B2(n_8_0_6989), .ZN(n_8_0_2130));
   AOI21_X1 i_8_0_1956 (.A(n_8_0_4857), .B1(n_8_0_4867), .B2(in_data[8]), 
      .ZN(n_8_0_2131));
   OR2_X1 i_8_0_1957 (.A1(n_8_0_4867), .A2(n_8_0_2133), .ZN(n_8_0_2132));
   AOI21_X1 i_8_0_1958 (.A(n_8_0_2134), .B1(n_8_0_2135), .B2(n_8_0_4864), 
      .ZN(n_8_0_2133));
   NOR2_X1 i_8_0_1959 (.A1(n_8_0_6991), .A2(n_8_0_4864), .ZN(n_8_0_2134));
   OAI21_X1 i_8_0_1960 (.A(n_8_0_2136), .B1(n_8_0_4860), .B2(n_8_0_6992), 
      .ZN(n_8_0_2135));
   OAI21_X1 i_8_0_1961 (.A(n_8_0_2137), .B1(n_8_0_2138), .B2(n_8_0_4851), 
      .ZN(n_8_0_2136));
   AOI21_X1 i_8_0_1962 (.A(n_8_0_4861), .B1(n_8_0_4851), .B2(n_8_0_6993), 
      .ZN(n_8_0_2137));
   MUX2_X1 i_8_0_1963 (.A(in_data[28]), .B(in_data[24]), .S(n_8_0_4854), 
      .Z(n_8_0_2138));
   OAI21_X1 i_8_0_1964 (.A(n_8_0_2139), .B1(n_8_0_2141), .B2(n_8_0_6988), 
      .ZN(n_58));
   OAI211_X1 i_8_0_1965 (.A(n_8_0_2141), .B(n_8_0_2140), .C1(n_8_0_2142), 
      .C2(n_8_0_4879), .ZN(n_8_0_2139));
   NAND2_X1 i_8_0_1966 (.A1(n_8_0_4879), .A2(n_8_0_6989), .ZN(n_8_0_2140));
   OAI21_X1 i_8_0_1967 (.A(n_8_0_4898), .B1(n_8_0_6729), .B2(n_8_0_4897), 
      .ZN(n_8_0_2141));
   OAI21_X1 i_8_0_1968 (.A(n_8_0_2143), .B1(n_8_0_4885), .B2(n_8_0_6990), 
      .ZN(n_8_0_2142));
   NAND2_X1 i_8_0_1969 (.A1(n_8_0_4885), .A2(n_8_0_2144), .ZN(n_8_0_2143));
   OAI21_X1 i_8_0_1970 (.A(n_8_0_2145), .B1(n_8_0_4882), .B2(n_8_0_6991), 
      .ZN(n_8_0_2144));
   NAND2_X1 i_8_0_1971 (.A1(n_8_0_4882), .A2(n_8_0_2146), .ZN(n_8_0_2145));
   MUX2_X1 i_8_0_1972 (.A(n_8_0_2147), .B(in_data[16]), .S(n_8_0_4888), .Z(
      n_8_0_2146));
   AOI21_X1 i_8_0_1973 (.A(n_8_0_2148), .B1(n_8_0_2149), .B2(n_8_0_4891), 
      .ZN(n_8_0_2147));
   NOR2_X1 i_8_0_1974 (.A1(n_8_0_4891), .A2(in_data[20]), .ZN(n_8_0_2148));
   OAI21_X1 i_8_0_1975 (.A(n_8_0_2150), .B1(n_8_0_4894), .B2(in_data[24]), 
      .ZN(n_8_0_2149));
   NAND2_X1 i_8_0_1976 (.A1(n_8_0_6995), .A2(n_8_0_4894), .ZN(n_8_0_2150));
   MUX2_X1 i_8_0_1977 (.A(in_data[0]), .B(n_8_0_2151), .S(n_8_0_2152), .Z(n_59));
   AOI22_X1 i_8_0_1978 (.A1(n_8_0_2153), .A2(n_8_0_2154), .B1(n_8_0_4920), 
      .B2(n_8_0_6989), .ZN(n_8_0_2151));
   OAI21_X1 i_8_0_1979 (.A(n_8_0_4912), .B1(n_8_0_6729), .B2(n_8_0_4911), 
      .ZN(n_8_0_2152));
   AOI21_X1 i_8_0_1980 (.A(n_8_0_4920), .B1(n_8_0_4923), .B2(in_data[8]), 
      .ZN(n_8_0_2153));
   OAI21_X1 i_8_0_1981 (.A(n_8_0_2155), .B1(n_8_0_2156), .B2(n_8_0_4917), 
      .ZN(n_8_0_2154));
   AOI21_X1 i_8_0_1982 (.A(n_8_0_4923), .B1(n_8_0_4917), .B2(n_8_0_6991), 
      .ZN(n_8_0_2155));
   AOI21_X1 i_8_0_1983 (.A(n_8_0_2157), .B1(n_8_0_4914), .B2(n_8_0_6992), 
      .ZN(n_8_0_2156));
   AOI211_X1 i_8_0_1984 (.A(n_8_0_4914), .B(n_8_0_2158), .C1(n_8_0_2159), 
      .C2(n_8_0_4908), .ZN(n_8_0_2157));
   NOR2_X1 i_8_0_1985 (.A1(n_8_0_6993), .A2(n_8_0_4908), .ZN(n_8_0_2158));
   OAI21_X1 i_8_0_1986 (.A(n_8_0_2160), .B1(n_8_0_4905), .B2(n_8_0_6994), 
      .ZN(n_8_0_2159));
   NAND2_X1 i_8_0_1987 (.A1(n_8_0_4905), .A2(in_data[28]), .ZN(n_8_0_2160));
   OAI21_X1 i_8_0_1988 (.A(n_8_0_2161), .B1(n_8_0_2169), .B2(n_8_0_6988), 
      .ZN(n_60));
   OAI211_X1 i_8_0_1989 (.A(n_8_0_2169), .B(n_8_0_2162), .C1(in_data[4]), 
      .C2(n_8_0_4945), .ZN(n_8_0_2161));
   OAI211_X1 i_8_0_1990 (.A(n_8_0_4945), .B(n_8_0_2163), .C1(n_8_0_4935), 
      .C2(n_8_0_6990), .ZN(n_8_0_2162));
   OAI211_X1 i_8_0_1991 (.A(n_8_0_2164), .B(n_8_0_4935), .C1(n_8_0_4948), 
      .C2(in_data[12]), .ZN(n_8_0_2163));
   OAI211_X1 i_8_0_1992 (.A(n_8_0_4948), .B(n_8_0_2165), .C1(n_8_0_4940), 
      .C2(n_8_0_6992), .ZN(n_8_0_2164));
   NAND2_X1 i_8_0_1993 (.A1(n_8_0_4940), .A2(n_8_0_2166), .ZN(n_8_0_2165));
   OAI21_X1 i_8_0_1994 (.A(n_8_0_2167), .B1(n_8_0_4928), .B2(n_8_0_6993), 
      .ZN(n_8_0_2166));
   NAND2_X1 i_8_0_1995 (.A1(n_8_0_4928), .A2(n_8_0_2168), .ZN(n_8_0_2167));
   MUX2_X1 i_8_0_1996 (.A(in_data[28]), .B(in_data[24]), .S(n_8_0_4938), 
      .Z(n_8_0_2168));
   NAND2_X1 i_8_0_1997 (.A1(n_8_0_4933), .A2(n_8_0_2170), .ZN(n_8_0_2169));
   OAI21_X1 i_8_0_1998 (.A(n_8_0_6730), .B1(n_8_0_4934), .B2(n_8_0_453), 
      .ZN(n_8_0_2170));
   MUX2_X1 i_8_0_1999 (.A(in_data[0]), .B(n_8_0_2171), .S(n_8_0_2180), .Z(n_61));
   AOI22_X1 i_8_0_2000 (.A1(n_8_0_2172), .A2(n_8_0_2173), .B1(n_8_0_4964), 
      .B2(n_8_0_6989), .ZN(n_8_0_2171));
   AOI21_X1 i_8_0_2001 (.A(n_8_0_4964), .B1(n_8_0_4970), .B2(in_data[8]), 
      .ZN(n_8_0_2172));
   OAI21_X1 i_8_0_2002 (.A(n_8_0_2174), .B1(n_8_0_2175), .B2(n_8_0_2177), 
      .ZN(n_8_0_2173));
   AOI21_X1 i_8_0_2003 (.A(n_8_0_4970), .B1(n_8_0_4973), .B2(n_8_0_6991), 
      .ZN(n_8_0_2174));
   AOI21_X1 i_8_0_2004 (.A(n_8_0_2176), .B1(n_8_0_2178), .B2(n_8_0_4961), 
      .ZN(n_8_0_2175));
   OAI21_X1 i_8_0_2005 (.A(n_8_0_4967), .B1(n_8_0_4961), .B2(in_data[20]), 
      .ZN(n_8_0_2176));
   OAI21_X1 i_8_0_2006 (.A(n_8_0_4974), .B1(n_8_0_4967), .B2(n_8_0_6992), 
      .ZN(n_8_0_2177));
   OAI21_X1 i_8_0_2007 (.A(n_8_0_2179), .B1(n_8_0_4959), .B2(in_data[24]), 
      .ZN(n_8_0_2178));
   NAND2_X1 i_8_0_2008 (.A1(n_8_0_6995), .A2(n_8_0_4959), .ZN(n_8_0_2179));
   AOI21_X1 i_8_0_2009 (.A(n_8_0_4957), .B1(n_8_0_4956), .B2(n_8_0_6729), 
      .ZN(n_8_0_2180));
   AOI21_X1 i_8_0_2010 (.A(n_8_0_2181), .B1(n_8_0_2184), .B2(n_8_0_2182), 
      .ZN(n_62));
   NOR2_X1 i_8_0_2011 (.A1(in_data[0]), .A2(n_8_0_2183), .ZN(n_8_0_2181));
   AOI221_X1 i_8_0_2012 (.A(n_8_0_4984), .B1(n_8_0_4985), .B2(n_8_0_6729), 
      .C1(in_data[4]), .C2(n_8_0_4998), .ZN(n_8_0_2182));
   AOI21_X1 i_8_0_2013 (.A(n_8_0_4984), .B1(n_8_0_4985), .B2(n_8_0_6729), 
      .ZN(n_8_0_2183));
   OAI21_X1 i_8_0_2014 (.A(n_8_0_2185), .B1(n_8_0_2186), .B2(n_8_0_4990), 
      .ZN(n_8_0_2184));
   AOI21_X1 i_8_0_2015 (.A(n_8_0_4998), .B1(n_8_0_4990), .B2(n_8_0_6990), 
      .ZN(n_8_0_2185));
   OAI21_X1 i_8_0_2016 (.A(n_8_0_2187), .B1(n_8_0_4995), .B2(n_8_0_6991), 
      .ZN(n_8_0_2186));
   OAI221_X1 i_8_0_2017 (.A(n_8_0_4995), .B1(n_8_0_2188), .B2(n_8_0_2190), 
      .C1(in_data[16]), .C2(n_8_0_4993), .ZN(n_8_0_2187));
   NAND2_X1 i_8_0_2018 (.A1(n_8_0_4993), .A2(n_8_0_2189), .ZN(n_8_0_2188));
   OAI211_X1 i_8_0_2019 (.A(n_8_0_4981), .B(n_8_0_2191), .C1(in_data[28]), 
      .C2(n_8_0_4987), .ZN(n_8_0_2189));
   NOR2_X1 i_8_0_2020 (.A1(n_8_0_4981), .A2(n_8_0_6993), .ZN(n_8_0_2190));
   NAND2_X1 i_8_0_2021 (.A1(n_8_0_4987), .A2(n_8_0_6994), .ZN(n_8_0_2191));
   MUX2_X1 i_8_0_2022 (.A(in_data[0]), .B(n_8_0_2192), .S(n_8_0_2193), .Z(n_63));
   MUX2_X1 i_8_0_2023 (.A(n_8_0_2194), .B(in_data[4]), .S(n_8_0_5027), .Z(
      n_8_0_2192));
   AOI21_X1 i_8_0_2024 (.A(n_8_0_5009), .B1(n_8_0_5008), .B2(n_8_0_6729), 
      .ZN(n_8_0_2193));
   MUX2_X1 i_8_0_2025 (.A(n_8_0_2195), .B(in_data[8]), .S(n_8_0_5014), .Z(
      n_8_0_2194));
   MUX2_X1 i_8_0_2026 (.A(n_8_0_2196), .B(in_data[12]), .S(n_8_0_5021), .Z(
      n_8_0_2195));
   MUX2_X1 i_8_0_2027 (.A(n_8_0_2197), .B(in_data[16]), .S(n_8_0_5017), .Z(
      n_8_0_2196));
   OAI21_X1 i_8_0_2028 (.A(n_8_0_2198), .B1(n_8_0_5012), .B2(n_8_0_6993), 
      .ZN(n_8_0_2197));
   NAND2_X1 i_8_0_2029 (.A1(n_8_0_2199), .A2(n_8_0_5012), .ZN(n_8_0_2198));
   OAI21_X1 i_8_0_2030 (.A(n_8_0_2200), .B1(n_8_0_5004), .B2(n_8_0_6995), 
      .ZN(n_8_0_2199));
   NAND2_X1 i_8_0_2031 (.A1(in_data[24]), .A2(n_8_0_5004), .ZN(n_8_0_2200));
   OAI22_X1 i_8_0_2032 (.A1(n_8_0_2202), .A2(n_8_0_2201), .B1(n_8_0_6988), 
      .B2(n_8_0_5055), .ZN(n_64));
   OAI21_X1 i_8_0_2033 (.A(n_8_0_5055), .B1(n_8_0_5033), .B2(in_data[4]), 
      .ZN(n_8_0_2201));
   AOI211_X1 i_8_0_2034 (.A(n_8_0_5034), .B(n_8_0_2203), .C1(in_data[8]), 
      .C2(n_8_0_5050), .ZN(n_8_0_2202));
   AOI21_X1 i_8_0_2035 (.A(n_8_0_2204), .B1(n_8_0_5058), .B2(n_8_0_6991), 
      .ZN(n_8_0_2203));
   OAI21_X1 i_8_0_2036 (.A(n_8_0_5049), .B1(n_8_0_2205), .B2(n_8_0_5058), 
      .ZN(n_8_0_2204));
   AOI21_X1 i_8_0_2037 (.A(n_8_0_2206), .B1(n_8_0_2207), .B2(n_8_0_5043), 
      .ZN(n_8_0_2205));
   NOR2_X1 i_8_0_2038 (.A1(n_8_0_5043), .A2(in_data[16]), .ZN(n_8_0_2206));
   OAI21_X1 i_8_0_2039 (.A(n_8_0_2208), .B1(n_8_0_2209), .B2(n_8_0_5039), 
      .ZN(n_8_0_2207));
   NAND2_X1 i_8_0_2040 (.A1(n_8_0_5039), .A2(n_8_0_6993), .ZN(n_8_0_2208));
   OAI21_X1 i_8_0_2041 (.A(n_8_0_2210), .B1(n_8_0_5045), .B2(n_8_0_6995), 
      .ZN(n_8_0_2209));
   NAND2_X1 i_8_0_2042 (.A1(in_data[24]), .A2(n_8_0_5045), .ZN(n_8_0_2210));
   MUX2_X1 i_8_0_2043 (.A(in_data[0]), .B(n_8_0_2211), .S(n_8_0_2220), .Z(n_65));
   AOI22_X1 i_8_0_2044 (.A1(n_8_0_2213), .A2(n_8_0_2212), .B1(n_8_0_6989), 
      .B2(n_8_0_5071), .ZN(n_8_0_2211));
   AOI21_X1 i_8_0_2045 (.A(n_8_0_5071), .B1(n_8_0_5069), .B2(in_data[8]), 
      .ZN(n_8_0_2212));
   OAI21_X1 i_8_0_2046 (.A(n_8_0_2214), .B1(n_8_0_2215), .B2(n_8_0_5065), 
      .ZN(n_8_0_2213));
   AOI21_X1 i_8_0_2047 (.A(n_8_0_5069), .B1(n_8_0_5065), .B2(n_8_0_6991), 
      .ZN(n_8_0_2214));
   AOI21_X1 i_8_0_2048 (.A(n_8_0_2216), .B1(n_8_0_5082), .B2(n_8_0_6992), 
      .ZN(n_8_0_2215));
   AOI211_X1 i_8_0_2049 (.A(n_8_0_5082), .B(n_8_0_2217), .C1(n_8_0_2218), 
      .C2(n_8_0_5077), .ZN(n_8_0_2216));
   NOR2_X1 i_8_0_2050 (.A1(n_8_0_6993), .A2(n_8_0_5077), .ZN(n_8_0_2217));
   OAI21_X1 i_8_0_2051 (.A(n_8_0_2219), .B1(n_8_0_5074), .B2(n_8_0_6994), 
      .ZN(n_8_0_2218));
   NAND2_X1 i_8_0_2052 (.A1(n_8_0_5074), .A2(in_data[28]), .ZN(n_8_0_2219));
   OAI21_X1 i_8_0_2053 (.A(n_8_0_2221), .B1(n_8_0_5080), .B2(n_8_0_6729), 
      .ZN(n_8_0_2220));
   OAI21_X1 i_8_0_2054 (.A(n_8_0_458), .B1(n_8_0_6730), .B2(n_8_0_5081), 
      .ZN(n_8_0_2221));
   MUX2_X1 i_8_0_2055 (.A(in_data[0]), .B(n_8_0_2222), .S(n_8_0_2233), .Z(n_66));
   AOI21_X1 i_8_0_2056 (.A(n_8_0_2223), .B1(n_8_0_5101), .B2(n_8_0_6989), 
      .ZN(n_8_0_2222));
   NOR2_X1 i_8_0_2057 (.A1(n_8_0_2224), .A2(n_8_0_5101), .ZN(n_8_0_2223));
   MUX2_X1 i_8_0_2058 (.A(n_8_0_2225), .B(in_data[8]), .S(n_8_0_5103), .Z(
      n_8_0_2224));
   OAI21_X1 i_8_0_2059 (.A(n_8_0_2232), .B1(n_8_0_2226), .B2(n_8_0_5106), 
      .ZN(n_8_0_2225));
   AOI21_X1 i_8_0_2060 (.A(n_8_0_2227), .B1(n_8_0_2228), .B2(n_8_0_5112), 
      .ZN(n_8_0_2226));
   NOR2_X1 i_8_0_2061 (.A1(n_8_0_5112), .A2(n_8_0_6992), .ZN(n_8_0_2227));
   OAI21_X1 i_8_0_2062 (.A(n_8_0_2229), .B1(n_8_0_5095), .B2(n_8_0_6993), 
      .ZN(n_8_0_2228));
   NAND2_X1 i_8_0_2063 (.A1(n_8_0_5095), .A2(n_8_0_2230), .ZN(n_8_0_2229));
   OAI21_X1 i_8_0_2064 (.A(n_8_0_2231), .B1(n_8_0_5110), .B2(n_8_0_6994), 
      .ZN(n_8_0_2230));
   NAND2_X1 i_8_0_2065 (.A1(n_8_0_5110), .A2(in_data[28]), .ZN(n_8_0_2231));
   NAND2_X1 i_8_0_2066 (.A1(in_data[12]), .A2(n_8_0_5106), .ZN(n_8_0_2232));
   OAI21_X1 i_8_0_2067 (.A(n_8_0_5092), .B1(n_8_0_6729), .B2(n_8_0_5093), 
      .ZN(n_8_0_2233));
   OAI22_X1 i_8_0_2068 (.A1(n_8_0_2235), .A2(n_8_0_2234), .B1(n_8_0_6988), 
      .B2(n_8_0_2244), .ZN(n_67));
   OAI21_X1 i_8_0_2069 (.A(n_8_0_2244), .B1(n_8_0_5126), .B2(in_data[4]), 
      .ZN(n_8_0_2234));
   AOI21_X1 i_8_0_2070 (.A(n_8_0_2236), .B1(n_8_0_2237), .B2(n_8_0_5138), 
      .ZN(n_8_0_2235));
   OAI21_X1 i_8_0_2071 (.A(n_8_0_5126), .B1(n_8_0_5138), .B2(n_8_0_6990), 
      .ZN(n_8_0_2236));
   OAI21_X1 i_8_0_2072 (.A(n_8_0_2238), .B1(n_8_0_5123), .B2(n_8_0_6991), 
      .ZN(n_8_0_2237));
   NAND2_X1 i_8_0_2073 (.A1(n_8_0_2239), .A2(n_8_0_5123), .ZN(n_8_0_2238));
   OAI21_X1 i_8_0_2074 (.A(n_8_0_2240), .B1(n_8_0_5141), .B2(n_8_0_6992), 
      .ZN(n_8_0_2239));
   OAI211_X1 i_8_0_2075 (.A(n_8_0_5141), .B(n_8_0_2241), .C1(n_8_0_2242), 
      .C2(n_8_0_5132), .ZN(n_8_0_2240));
   NAND2_X1 i_8_0_2076 (.A1(n_8_0_5132), .A2(n_8_0_6993), .ZN(n_8_0_2241));
   OAI21_X1 i_8_0_2077 (.A(n_8_0_2243), .B1(n_8_0_5129), .B2(n_8_0_6994), 
      .ZN(n_8_0_2242));
   NAND2_X1 i_8_0_2078 (.A1(n_8_0_5129), .A2(in_data[28]), .ZN(n_8_0_2243));
   OAI21_X1 i_8_0_2079 (.A(n_8_0_5136), .B1(n_8_0_6729), .B2(n_8_0_5135), 
      .ZN(n_8_0_2244));
   AOI22_X1 i_8_0_2080 (.A1(n_8_0_2245), .A2(n_8_0_2247), .B1(n_8_0_6988), 
      .B2(n_8_0_2246), .ZN(n_68));
   AOI21_X1 i_8_0_2081 (.A(n_8_0_2246), .B1(n_8_0_5153), .B2(in_data[4]), 
      .ZN(n_8_0_2245));
   OAI21_X1 i_8_0_2082 (.A(n_8_0_5166), .B1(n_8_0_5165), .B2(n_8_0_6730), 
      .ZN(n_8_0_2246));
   NAND2_X1 i_8_0_2083 (.A1(n_8_0_5154), .A2(n_8_0_2248), .ZN(n_8_0_2247));
   OAI21_X1 i_8_0_2084 (.A(n_8_0_2256), .B1(n_8_0_2249), .B2(n_8_0_5157), 
      .ZN(n_8_0_2248));
   AOI21_X1 i_8_0_2085 (.A(n_8_0_2250), .B1(n_8_0_2251), .B2(n_8_0_5150), 
      .ZN(n_8_0_2249));
   NOR2_X1 i_8_0_2086 (.A1(n_8_0_5150), .A2(n_8_0_6991), .ZN(n_8_0_2250));
   OAI21_X1 i_8_0_2087 (.A(n_8_0_2252), .B1(n_8_0_5147), .B2(n_8_0_6992), 
      .ZN(n_8_0_2251));
   NAND2_X1 i_8_0_2088 (.A1(n_8_0_2253), .A2(n_8_0_5147), .ZN(n_8_0_2252));
   MUX2_X1 i_8_0_2089 (.A(n_8_0_2254), .B(in_data[20]), .S(n_8_0_5162), .Z(
      n_8_0_2253));
   OAI21_X1 i_8_0_2090 (.A(n_8_0_2255), .B1(n_8_0_5168), .B2(n_8_0_6995), 
      .ZN(n_8_0_2254));
   NAND2_X1 i_8_0_2091 (.A1(in_data[24]), .A2(n_8_0_5168), .ZN(n_8_0_2255));
   NAND2_X1 i_8_0_2092 (.A1(n_8_0_5157), .A2(in_data[8]), .ZN(n_8_0_2256));
   OAI22_X1 i_8_0_2093 (.A1(n_8_0_2258), .A2(n_8_0_2257), .B1(n_8_0_6988), 
      .B2(n_8_0_2265), .ZN(n_69));
   OAI21_X1 i_8_0_2094 (.A(n_8_0_2265), .B1(n_8_0_5182), .B2(in_data[4]), 
      .ZN(n_8_0_2257));
   AOI221_X1 i_8_0_2095 (.A(n_8_0_5181), .B1(n_8_0_2259), .B2(n_8_0_2260), 
      .C1(in_data[8]), .C2(n_8_0_5176), .ZN(n_8_0_2258));
   NOR2_X1 i_8_0_2096 (.A1(n_8_0_2261), .A2(n_8_0_5176), .ZN(n_8_0_2259));
   NAND2_X1 i_8_0_2097 (.A1(n_8_0_5195), .A2(n_8_0_6991), .ZN(n_8_0_2260));
   AOI221_X1 i_8_0_2098 (.A(n_8_0_5195), .B1(n_8_0_2263), .B2(n_8_0_2262), 
      .C1(n_8_0_5178), .C2(in_data[16]), .ZN(n_8_0_2261));
   AOI21_X1 i_8_0_2099 (.A(n_8_0_5178), .B1(n_8_0_5186), .B2(n_8_0_6993), 
      .ZN(n_8_0_2262));
   OAI21_X1 i_8_0_2100 (.A(n_8_0_2264), .B1(n_8_0_5188), .B2(n_8_0_6994), 
      .ZN(n_8_0_2263));
   AOI21_X1 i_8_0_2101 (.A(n_8_0_5186), .B1(n_8_0_5188), .B2(in_data[28]), 
      .ZN(n_8_0_2264));
   AOI21_X1 i_8_0_2102 (.A(n_8_0_5192), .B1(n_8_0_5193), .B2(n_8_0_6729), 
      .ZN(n_8_0_2265));
   OAI22_X1 i_8_0_2103 (.A1(n_8_0_2267), .A2(n_8_0_2266), .B1(n_8_0_6988), 
      .B2(n_8_0_2277), .ZN(n_70));
   OAI21_X1 i_8_0_2104 (.A(n_8_0_2277), .B1(n_8_0_5204), .B2(in_data[4]), 
      .ZN(n_8_0_2266));
   AOI21_X1 i_8_0_2105 (.A(n_8_0_2268), .B1(n_8_0_2269), .B2(n_8_0_5206), 
      .ZN(n_8_0_2267));
   OAI21_X1 i_8_0_2106 (.A(n_8_0_5204), .B1(n_8_0_5206), .B2(n_8_0_6990), 
      .ZN(n_8_0_2268));
   OAI21_X1 i_8_0_2107 (.A(n_8_0_2270), .B1(n_8_0_2271), .B2(n_8_0_5219), 
      .ZN(n_8_0_2269));
   NAND2_X1 i_8_0_2108 (.A1(in_data[12]), .A2(n_8_0_5219), .ZN(n_8_0_2270));
   AOI21_X1 i_8_0_2109 (.A(n_8_0_2272), .B1(n_8_0_2273), .B2(n_8_0_5225), 
      .ZN(n_8_0_2271));
   NOR2_X1 i_8_0_2110 (.A1(n_8_0_5225), .A2(n_8_0_6992), .ZN(n_8_0_2272));
   OAI21_X1 i_8_0_2111 (.A(n_8_0_2274), .B1(n_8_0_2275), .B2(n_8_0_5213), 
      .ZN(n_8_0_2273));
   NAND2_X1 i_8_0_2112 (.A1(n_8_0_5213), .A2(in_data[20]), .ZN(n_8_0_2274));
   OAI21_X1 i_8_0_2113 (.A(n_8_0_2276), .B1(n_8_0_5209), .B2(in_data[24]), 
      .ZN(n_8_0_2275));
   NAND2_X1 i_8_0_2114 (.A1(n_8_0_6995), .A2(n_8_0_5209), .ZN(n_8_0_2276));
   AOI21_X1 i_8_0_2115 (.A(n_8_0_5216), .B1(n_8_0_5217), .B2(n_8_0_6729), 
      .ZN(n_8_0_2277));
   OAI22_X1 i_8_0_2116 (.A1(n_8_0_2279), .A2(n_8_0_2278), .B1(n_8_0_6988), 
      .B2(n_8_0_5247), .ZN(n_71));
   OAI21_X1 i_8_0_2117 (.A(n_8_0_5247), .B1(n_8_0_5240), .B2(in_data[4]), 
      .ZN(n_8_0_2278));
   AOI221_X1 i_8_0_2118 (.A(n_8_0_5239), .B1(n_8_0_2280), .B2(n_8_0_2281), 
      .C1(in_data[8]), .C2(n_8_0_5234), .ZN(n_8_0_2279));
   AOI21_X1 i_8_0_2119 (.A(n_8_0_5234), .B1(n_8_0_5250), .B2(n_8_0_6991), 
      .ZN(n_8_0_2280));
   OAI21_X1 i_8_0_2120 (.A(n_8_0_2282), .B1(n_8_0_2283), .B2(n_8_0_5236), 
      .ZN(n_8_0_2281));
   AOI21_X1 i_8_0_2121 (.A(n_8_0_5250), .B1(n_8_0_5236), .B2(in_data[16]), 
      .ZN(n_8_0_2282));
   AOI21_X1 i_8_0_2122 (.A(n_8_0_2284), .B1(n_8_0_2285), .B2(n_8_0_5242), 
      .ZN(n_8_0_2283));
   NOR2_X1 i_8_0_2123 (.A1(n_8_0_5242), .A2(n_8_0_6993), .ZN(n_8_0_2284));
   OAI21_X1 i_8_0_2124 (.A(n_8_0_2286), .B1(n_8_0_5244), .B2(n_8_0_6994), 
      .ZN(n_8_0_2285));
   NAND2_X1 i_8_0_2125 (.A1(n_8_0_5244), .A2(in_data[28]), .ZN(n_8_0_2286));
   OAI21_X1 i_8_0_2126 (.A(n_8_0_2287), .B1(n_8_0_2297), .B2(n_8_0_6988), 
      .ZN(n_72));
   OAI211_X1 i_8_0_2127 (.A(n_8_0_2297), .B(n_8_0_2288), .C1(in_data[4]), 
      .C2(n_8_0_5270), .ZN(n_8_0_2287));
   OAI211_X1 i_8_0_2128 (.A(n_8_0_5270), .B(n_8_0_2289), .C1(n_8_0_2290), 
      .C2(n_8_0_5265), .ZN(n_8_0_2288));
   NAND2_X1 i_8_0_2129 (.A1(in_data[8]), .A2(n_8_0_5265), .ZN(n_8_0_2289));
   INV_X1 i_8_0_2130 (.A(n_8_0_2291), .ZN(n_8_0_2290));
   MUX2_X1 i_8_0_2131 (.A(n_8_0_2292), .B(in_data[12]), .S(n_8_0_5276), .Z(
      n_8_0_2291));
   OAI22_X1 i_8_0_2132 (.A1(n_8_0_2295), .A2(n_8_0_2293), .B1(n_8_0_6992), 
      .B2(n_8_0_5268), .ZN(n_8_0_2292));
   NAND2_X1 i_8_0_2133 (.A1(n_8_0_2294), .A2(n_8_0_5268), .ZN(n_8_0_2293));
   OAI211_X1 i_8_0_2134 (.A(n_8_0_5257), .B(n_8_0_2296), .C1(n_8_0_6995), 
      .C2(n_8_0_5261), .ZN(n_8_0_2294));
   NOR2_X1 i_8_0_2135 (.A1(n_8_0_5257), .A2(in_data[20]), .ZN(n_8_0_2295));
   NAND2_X1 i_8_0_2136 (.A1(in_data[24]), .A2(n_8_0_5261), .ZN(n_8_0_2296));
   AOI21_X1 i_8_0_2137 (.A(n_8_0_2298), .B1(n_8_0_5481), .B2(n_8_0_6729), 
      .ZN(n_8_0_2297));
   AOI21_X1 i_8_0_2138 (.A(n_8_0_465), .B1(n_8_0_6730), .B2(n_8_0_5482), 
      .ZN(n_8_0_2298));
   MUX2_X1 i_8_0_2139 (.A(in_data[0]), .B(n_8_0_2299), .S(n_8_0_2300), .Z(n_73));
   AOI21_X1 i_8_0_2140 (.A(n_8_0_2301), .B1(n_8_0_5293), .B2(n_8_0_6989), 
      .ZN(n_8_0_2299));
   AOI21_X1 i_8_0_2141 (.A(n_8_0_5285), .B1(n_8_0_5286), .B2(n_8_0_6729), 
      .ZN(n_8_0_2300));
   AOI211_X1 i_8_0_2142 (.A(n_8_0_5293), .B(n_8_0_2302), .C1(in_data[8]), 
      .C2(n_8_0_5299), .ZN(n_8_0_2301));
   AOI211_X1 i_8_0_2143 (.A(n_8_0_5299), .B(n_8_0_2303), .C1(n_8_0_2304), 
      .C2(n_8_0_5295), .ZN(n_8_0_2302));
   NOR2_X1 i_8_0_2144 (.A1(n_8_0_5295), .A2(in_data[12]), .ZN(n_8_0_2303));
   INV_X1 i_8_0_2145 (.A(n_8_0_2305), .ZN(n_8_0_2304));
   OAI21_X1 i_8_0_2146 (.A(n_8_0_2306), .B1(n_8_0_2307), .B2(n_8_0_5303), 
      .ZN(n_8_0_2305));
   NAND2_X1 i_8_0_2147 (.A1(n_8_0_5303), .A2(in_data[16]), .ZN(n_8_0_2306));
   OAI21_X1 i_8_0_2148 (.A(n_8_0_2308), .B1(n_8_0_2309), .B2(n_8_0_5288), 
      .ZN(n_8_0_2307));
   NAND2_X1 i_8_0_2149 (.A1(n_8_0_5288), .A2(n_8_0_6993), .ZN(n_8_0_2308));
   OAI21_X1 i_8_0_2150 (.A(n_8_0_2310), .B1(n_8_0_5290), .B2(n_8_0_6994), 
      .ZN(n_8_0_2309));
   NAND2_X1 i_8_0_2151 (.A1(n_8_0_5290), .A2(in_data[28]), .ZN(n_8_0_2310));
   AOI21_X1 i_8_0_2152 (.A(n_8_0_2311), .B1(n_8_0_2312), .B2(n_8_0_2313), 
      .ZN(n_74));
   NOR2_X1 i_8_0_2153 (.A1(in_data[0]), .A2(n_8_0_2313), .ZN(n_8_0_2311));
   MUX2_X1 i_8_0_2154 (.A(n_8_0_2314), .B(n_8_0_6989), .S(n_8_0_5318), .Z(
      n_8_0_2312));
   OAI21_X1 i_8_0_2155 (.A(n_8_0_5310), .B1(n_8_0_6729), .B2(n_8_0_5311), 
      .ZN(n_8_0_2313));
   AOI21_X1 i_8_0_2156 (.A(n_8_0_2315), .B1(n_8_0_5321), .B2(in_data[8]), 
      .ZN(n_8_0_2314));
   AOI211_X1 i_8_0_2157 (.A(n_8_0_2316), .B(n_8_0_5321), .C1(n_8_0_5328), 
      .C2(n_8_0_2317), .ZN(n_8_0_2315));
   NOR2_X1 i_8_0_2158 (.A1(n_8_0_5328), .A2(in_data[12]), .ZN(n_8_0_2316));
   AOI21_X1 i_8_0_2159 (.A(n_8_0_2318), .B1(n_8_0_5323), .B2(in_data[16]), 
      .ZN(n_8_0_2317));
   AOI221_X1 i_8_0_2160 (.A(n_8_0_5323), .B1(n_8_0_5312), .B2(n_8_0_6993), 
      .C1(n_8_0_2319), .C2(n_8_0_2320), .ZN(n_8_0_2318));
   AOI21_X1 i_8_0_2161 (.A(n_8_0_5312), .B1(n_8_0_5326), .B2(in_data[24]), 
      .ZN(n_8_0_2319));
   OR2_X1 i_8_0_2162 (.A1(n_8_0_6995), .A2(n_8_0_5326), .ZN(n_8_0_2320));
   AOI22_X1 i_8_0_2163 (.A1(n_8_0_2321), .A2(n_8_0_2323), .B1(n_8_0_6988), 
      .B2(n_8_0_2322), .ZN(n_75));
   AOI21_X1 i_8_0_2164 (.A(n_8_0_2322), .B1(n_8_0_5351), .B2(in_data[4]), 
      .ZN(n_8_0_2321));
   OAI21_X1 i_8_0_2165 (.A(n_8_0_5342), .B1(n_8_0_5343), .B2(n_8_0_6730), 
      .ZN(n_8_0_2322));
   OAI21_X1 i_8_0_2166 (.A(n_8_0_2324), .B1(n_8_0_2325), .B2(n_8_0_5353), 
      .ZN(n_8_0_2323));
   AOI21_X1 i_8_0_2167 (.A(n_8_0_5351), .B1(n_8_0_5353), .B2(n_8_0_6990), 
      .ZN(n_8_0_2324));
   MUX2_X1 i_8_0_2168 (.A(in_data[12]), .B(n_8_0_2326), .S(n_8_0_5348), .Z(
      n_8_0_2325));
   AOI21_X1 i_8_0_2169 (.A(n_8_0_2327), .B1(n_8_0_2328), .B2(n_8_0_5345), 
      .ZN(n_8_0_2326));
   NOR2_X1 i_8_0_2170 (.A1(in_data[16]), .A2(n_8_0_5345), .ZN(n_8_0_2327));
   OAI21_X1 i_8_0_2171 (.A(n_8_0_2329), .B1(n_8_0_5335), .B2(in_data[20]), 
      .ZN(n_8_0_2328));
   OAI211_X1 i_8_0_2172 (.A(n_8_0_5335), .B(n_8_0_2330), .C1(n_8_0_6995), 
      .C2(n_8_0_5339), .ZN(n_8_0_2329));
   NAND2_X1 i_8_0_2173 (.A1(n_8_0_5339), .A2(in_data[24]), .ZN(n_8_0_2330));
   MUX2_X1 i_8_0_2174 (.A(n_8_0_2331), .B(in_data[0]), .S(n_8_0_2333), .Z(n_76));
   OAI21_X1 i_8_0_2175 (.A(n_8_0_2332), .B1(n_8_0_5368), .B2(n_8_0_6989), 
      .ZN(n_8_0_2331));
   NAND3_X1 i_8_0_2176 (.A1(n_8_0_5368), .A2(n_8_0_2337), .A3(n_8_0_2336), 
      .ZN(n_8_0_2332));
   OAI21_X1 i_8_0_2177 (.A(n_8_0_2334), .B1(n_8_0_5480), .B2(n_8_0_6730), 
      .ZN(n_8_0_2333));
   INV_X1 i_8_0_2178 (.A(n_8_0_2335), .ZN(n_8_0_2334));
   AOI21_X1 i_8_0_2179 (.A(n_8_0_469), .B1(n_8_0_6730), .B2(n_8_0_5480), 
      .ZN(n_8_0_2335));
   NAND2_X1 i_8_0_2180 (.A1(n_8_0_6990), .A2(n_8_0_5377), .ZN(n_8_0_2336));
   OAI21_X1 i_8_0_2181 (.A(n_8_0_2338), .B1(n_8_0_2339), .B2(n_8_0_5371), 
      .ZN(n_8_0_2337));
   AOI21_X1 i_8_0_2182 (.A(n_8_0_5377), .B1(n_8_0_5371), .B2(in_data[12]), 
      .ZN(n_8_0_2338));
   INV_X1 i_8_0_2183 (.A(n_8_0_2340), .ZN(n_8_0_2339));
   OAI21_X1 i_8_0_2184 (.A(n_8_0_2341), .B1(n_8_0_2342), .B2(n_8_0_5374), 
      .ZN(n_8_0_2340));
   NAND2_X1 i_8_0_2185 (.A1(in_data[16]), .A2(n_8_0_5374), .ZN(n_8_0_2341));
   OAI21_X1 i_8_0_2186 (.A(n_8_0_2343), .B1(n_8_0_5362), .B2(in_data[20]), 
      .ZN(n_8_0_2342));
   OAI211_X1 i_8_0_2187 (.A(n_8_0_5362), .B(n_8_0_2344), .C1(n_8_0_6995), 
      .C2(n_8_0_5365), .ZN(n_8_0_2343));
   NAND2_X1 i_8_0_2188 (.A1(n_8_0_5365), .A2(in_data[24]), .ZN(n_8_0_2344));
   OAI22_X1 i_8_0_2189 (.A1(n_8_0_2348), .A2(n_8_0_2345), .B1(n_8_0_2346), 
      .B2(n_8_0_6988), .ZN(n_77));
   OAI21_X1 i_8_0_2190 (.A(n_8_0_2346), .B1(n_8_0_5384), .B2(in_data[4]), 
      .ZN(n_8_0_2345));
   OAI21_X1 i_8_0_2191 (.A(n_8_0_2347), .B1(n_8_0_5404), .B2(n_8_0_6729), 
      .ZN(n_8_0_2346));
   OAI21_X1 i_8_0_2192 (.A(n_8_0_470), .B1(n_8_0_6730), .B2(n_8_0_5403), 
      .ZN(n_8_0_2347));
   AOI221_X1 i_8_0_2193 (.A(n_8_0_5383), .B1(n_8_0_2350), .B2(n_8_0_2349), 
      .C1(n_8_0_5405), .C2(in_data[8]), .ZN(n_8_0_2348));
   AOI21_X1 i_8_0_2194 (.A(n_8_0_5405), .B1(n_8_0_5407), .B2(n_8_0_6991), 
      .ZN(n_8_0_2349));
   OAI21_X1 i_8_0_2195 (.A(n_8_0_2351), .B1(n_8_0_2352), .B2(n_8_0_5388), 
      .ZN(n_8_0_2350));
   AOI21_X1 i_8_0_2196 (.A(n_8_0_5407), .B1(n_8_0_5388), .B2(in_data[16]), 
      .ZN(n_8_0_2351));
   AOI22_X1 i_8_0_2197 (.A1(n_8_0_2353), .A2(n_8_0_2355), .B1(n_8_0_5398), 
      .B2(in_data[20]), .ZN(n_8_0_2352));
   NOR2_X1 i_8_0_2198 (.A1(n_8_0_5398), .A2(n_8_0_2354), .ZN(n_8_0_2353));
   NOR2_X1 i_8_0_2199 (.A1(in_data[28]), .A2(n_8_0_5392), .ZN(n_8_0_2354));
   NAND2_X1 i_8_0_2200 (.A1(n_8_0_5392), .A2(n_8_0_6994), .ZN(n_8_0_2355));
   AOI22_X1 i_8_0_2201 (.A1(n_8_0_2356), .A2(n_8_0_2358), .B1(n_8_0_6988), 
      .B2(n_8_0_2357), .ZN(n_78));
   AOI21_X1 i_8_0_2202 (.A(n_8_0_2357), .B1(n_8_0_5419), .B2(in_data[4]), 
      .ZN(n_8_0_2356));
   OAI21_X1 i_8_0_2203 (.A(n_8_0_5433), .B1(n_8_0_5435), .B2(n_8_0_6730), 
      .ZN(n_8_0_2357));
   OAI21_X1 i_8_0_2204 (.A(n_8_0_2359), .B1(n_8_0_2360), .B2(n_8_0_5416), 
      .ZN(n_8_0_2358));
   AOI21_X1 i_8_0_2205 (.A(n_8_0_5419), .B1(n_8_0_5416), .B2(n_8_0_6990), 
      .ZN(n_8_0_2359));
   AOI21_X1 i_8_0_2206 (.A(n_8_0_2361), .B1(n_8_0_5438), .B2(n_8_0_6991), 
      .ZN(n_8_0_2360));
   NOR2_X1 i_8_0_2207 (.A1(n_8_0_5438), .A2(n_8_0_2362), .ZN(n_8_0_2361));
   MUX2_X1 i_8_0_2208 (.A(in_data[16]), .B(n_8_0_2363), .S(n_8_0_5414), .Z(
      n_8_0_2362));
   AOI22_X1 i_8_0_2209 (.A1(n_8_0_2364), .A2(n_8_0_2365), .B1(n_8_0_5423), 
      .B2(n_8_0_6993), .ZN(n_8_0_2363));
   AOI21_X1 i_8_0_2210 (.A(n_8_0_5423), .B1(n_8_0_5429), .B2(in_data[28]), 
      .ZN(n_8_0_2364));
   NAND2_X1 i_8_0_2211 (.A1(n_8_0_5430), .A2(in_data[24]), .ZN(n_8_0_2365));
   OAI22_X1 i_8_0_2212 (.A1(n_8_0_2367), .A2(n_8_0_2366), .B1(n_8_0_6988), 
      .B2(n_8_0_2375), .ZN(n_79));
   OAI21_X1 i_8_0_2213 (.A(n_8_0_2375), .B1(n_8_0_5449), .B2(in_data[4]), 
      .ZN(n_8_0_2366));
   AOI211_X1 i_8_0_2214 (.A(n_8_0_5448), .B(n_8_0_2368), .C1(in_data[8]), 
      .C2(n_8_0_5469), .ZN(n_8_0_2367));
   NOR2_X1 i_8_0_2215 (.A1(n_8_0_5469), .A2(n_8_0_2369), .ZN(n_8_0_2368));
   AOI21_X1 i_8_0_2216 (.A(n_8_0_2370), .B1(n_8_0_2371), .B2(n_8_0_5457), 
      .ZN(n_8_0_2369));
   NOR2_X1 i_8_0_2217 (.A1(n_8_0_6991), .A2(n_8_0_5457), .ZN(n_8_0_2370));
   AOI21_X1 i_8_0_2218 (.A(n_8_0_2372), .B1(n_8_0_5463), .B2(n_8_0_6992), 
      .ZN(n_8_0_2371));
   AOI211_X1 i_8_0_2219 (.A(n_8_0_5463), .B(n_8_0_2373), .C1(in_data[20]), 
      .C2(n_8_0_5473), .ZN(n_8_0_2372));
   AOI211_X1 i_8_0_2220 (.A(n_8_0_2374), .B(n_8_0_5473), .C1(n_8_0_5476), 
      .C2(n_8_0_6994), .ZN(n_8_0_2373));
   NOR2_X1 i_8_0_2221 (.A1(n_8_0_5476), .A2(in_data[28]), .ZN(n_8_0_2374));
   OAI21_X1 i_8_0_2222 (.A(n_8_0_5478), .B1(n_8_0_6729), .B2(n_8_0_5479), 
      .ZN(n_8_0_2375));
   MUX2_X1 i_8_0_2223 (.A(n_8_0_2376), .B(in_data[0]), .S(n_8_0_2386), .Z(n_80));
   AOI22_X1 i_8_0_2224 (.A1(n_8_0_2377), .A2(n_8_0_2378), .B1(n_8_0_5490), 
      .B2(n_8_0_6989), .ZN(n_8_0_2376));
   AOI21_X1 i_8_0_2225 (.A(n_8_0_5490), .B1(n_8_0_5491), .B2(in_data[8]), 
      .ZN(n_8_0_2377));
   NAND2_X1 i_8_0_2226 (.A1(n_8_0_2379), .A2(n_8_0_2380), .ZN(n_8_0_2378));
   AOI21_X1 i_8_0_2227 (.A(n_8_0_5491), .B1(n_8_0_5489), .B2(n_8_0_6991), 
      .ZN(n_8_0_2379));
   OAI21_X1 i_8_0_2228 (.A(n_8_0_2381), .B1(n_8_0_2382), .B2(n_8_0_5496), 
      .ZN(n_8_0_2380));
   AOI21_X1 i_8_0_2229 (.A(n_8_0_5489), .B1(n_8_0_5496), .B2(in_data[16]), 
      .ZN(n_8_0_2381));
   OAI21_X1 i_8_0_2230 (.A(n_8_0_2383), .B1(n_8_0_2384), .B2(n_8_0_5492), 
      .ZN(n_8_0_2382));
   NAND2_X1 i_8_0_2231 (.A1(n_8_0_5492), .A2(n_8_0_6993), .ZN(n_8_0_2383));
   OAI21_X1 i_8_0_2232 (.A(n_8_0_2385), .B1(n_8_0_5495), .B2(n_8_0_6995), 
      .ZN(n_8_0_2384));
   NAND2_X1 i_8_0_2233 (.A1(n_8_0_5495), .A2(in_data[24]), .ZN(n_8_0_2385));
   OAI21_X1 i_8_0_2234 (.A(n_8_0_6464), .B1(n_8_0_6718), .B2(n_8_0_473), 
      .ZN(n_8_0_2386));
   NOR2_X1 i_8_0_2235 (.A1(n_8_0_2395), .A2(n_8_0_2387), .ZN(n_81));
   AOI21_X1 i_8_0_2236 (.A(n_8_0_2388), .B1(n_8_0_2389), .B2(n_8_0_5520), 
      .ZN(n_8_0_2387));
   OAI21_X1 i_8_0_2237 (.A(n_8_0_2396), .B1(n_8_0_5520), .B2(n_8_0_6989), 
      .ZN(n_8_0_2388));
   MUX2_X1 i_8_0_2238 (.A(in_data[8]), .B(n_8_0_2390), .S(n_8_0_5516), .Z(
      n_8_0_2389));
   MUX2_X1 i_8_0_2239 (.A(n_8_0_2391), .B(in_data[12]), .S(n_8_0_5527), .Z(
      n_8_0_2390));
   AOI21_X1 i_8_0_2240 (.A(n_8_0_2392), .B1(n_8_0_5498), .B2(n_8_0_6992), 
      .ZN(n_8_0_2391));
   AOI211_X1 i_8_0_2241 (.A(n_8_0_5498), .B(n_8_0_2393), .C1(in_data[20]), 
      .C2(n_8_0_5512), .ZN(n_8_0_2392));
   AOI21_X1 i_8_0_2242 (.A(n_8_0_2394), .B1(n_8_0_5523), .B2(n_8_0_6995), 
      .ZN(n_8_0_2393));
   OAI21_X1 i_8_0_2243 (.A(n_8_0_5513), .B1(n_8_0_5523), .B2(in_data[24]), 
      .ZN(n_8_0_2394));
   NOR2_X1 i_8_0_2244 (.A1(n_8_0_2396), .A2(in_data[0]), .ZN(n_8_0_2395));
   AOI21_X1 i_8_0_2245 (.A(n_8_0_5509), .B1(n_8_0_5510), .B2(n_8_0_6729), 
      .ZN(n_8_0_2396));
   MUX2_X1 i_8_0_2246 (.A(in_data[0]), .B(n_8_0_2397), .S(n_8_0_2407), .Z(n_82));
   AOI22_X1 i_8_0_2247 (.A1(n_8_0_2398), .A2(n_8_0_2399), .B1(n_8_0_5541), 
      .B2(n_8_0_6989), .ZN(n_8_0_2397));
   AOI21_X1 i_8_0_2248 (.A(n_8_0_5541), .B1(n_8_0_5538), .B2(in_data[8]), 
      .ZN(n_8_0_2398));
   NAND2_X1 i_8_0_2249 (.A1(n_8_0_5537), .A2(n_8_0_2400), .ZN(n_8_0_2399));
   MUX2_X1 i_8_0_2250 (.A(n_8_0_2401), .B(in_data[12]), .S(n_8_0_5534), .Z(
      n_8_0_2400));
   AOI21_X1 i_8_0_2251 (.A(n_8_0_2402), .B1(n_8_0_2403), .B2(n_8_0_5561), 
      .ZN(n_8_0_2401));
   NOR2_X1 i_8_0_2252 (.A1(n_8_0_5561), .A2(in_data[16]), .ZN(n_8_0_2402));
   OAI21_X1 i_8_0_2253 (.A(n_8_0_2404), .B1(n_8_0_2405), .B2(n_8_0_5549), 
      .ZN(n_8_0_2403));
   NAND2_X1 i_8_0_2254 (.A1(n_8_0_5549), .A2(n_8_0_6993), .ZN(n_8_0_2404));
   OAI21_X1 i_8_0_2255 (.A(n_8_0_2406), .B1(n_8_0_5545), .B2(n_8_0_6994), 
      .ZN(n_8_0_2405));
   NAND2_X1 i_8_0_2256 (.A1(n_8_0_5545), .A2(in_data[28]), .ZN(n_8_0_2406));
   AOI21_X1 i_8_0_2257 (.A(n_8_0_5555), .B1(n_8_0_5558), .B2(n_8_0_6729), 
      .ZN(n_8_0_2407));
   MUX2_X1 i_8_0_2258 (.A(in_data[0]), .B(n_8_0_2408), .S(n_8_0_2417), .Z(n_83));
   AOI22_X1 i_8_0_2259 (.A1(n_8_0_2409), .A2(n_8_0_2410), .B1(n_8_0_5582), 
      .B2(n_8_0_6989), .ZN(n_8_0_2408));
   AOI21_X1 i_8_0_2260 (.A(n_8_0_5582), .B1(n_8_0_5574), .B2(in_data[8]), 
      .ZN(n_8_0_2409));
   NAND2_X1 i_8_0_2261 (.A1(n_8_0_2411), .A2(n_8_0_5575), .ZN(n_8_0_2410));
   OAI21_X1 i_8_0_2262 (.A(n_8_0_2412), .B1(n_8_0_5570), .B2(n_8_0_6991), 
      .ZN(n_8_0_2411));
   OAI211_X1 i_8_0_2263 (.A(n_8_0_5570), .B(n_8_0_2413), .C1(in_data[16]), 
      .C2(n_8_0_5578), .ZN(n_8_0_2412));
   NAND2_X1 i_8_0_2264 (.A1(n_8_0_5578), .A2(n_8_0_2414), .ZN(n_8_0_2413));
   OAI21_X1 i_8_0_2265 (.A(n_8_0_2415), .B1(n_8_0_5587), .B2(in_data[20]), 
      .ZN(n_8_0_2414));
   OAI211_X1 i_8_0_2266 (.A(n_8_0_5587), .B(n_8_0_2416), .C1(n_8_0_5584), 
      .C2(n_8_0_6995), .ZN(n_8_0_2415));
   NAND2_X1 i_8_0_2267 (.A1(in_data[24]), .A2(n_8_0_5584), .ZN(n_8_0_2416));
   AOI21_X1 i_8_0_2268 (.A(n_8_0_5591), .B1(n_8_0_5592), .B2(n_8_0_6729), 
      .ZN(n_8_0_2417));
   OAI21_X1 i_8_0_2269 (.A(n_8_0_2418), .B1(n_8_0_2428), .B2(n_8_0_6988), 
      .ZN(n_84));
   OAI211_X1 i_8_0_2270 (.A(n_8_0_2428), .B(n_8_0_2419), .C1(in_data[4]), 
      .C2(n_8_0_5623), .ZN(n_8_0_2418));
   OAI211_X1 i_8_0_2271 (.A(n_8_0_5623), .B(n_8_0_2427), .C1(n_8_0_2420), 
      .C2(n_8_0_5600), .ZN(n_8_0_2419));
   OAI21_X1 i_8_0_2272 (.A(n_8_0_2421), .B1(n_8_0_2422), .B2(n_8_0_5603), 
      .ZN(n_8_0_2420));
   NAND2_X1 i_8_0_2273 (.A1(n_8_0_5603), .A2(n_8_0_6991), .ZN(n_8_0_2421));
   OAI21_X1 i_8_0_2274 (.A(n_8_0_2426), .B1(n_8_0_2423), .B2(n_8_0_5597), 
      .ZN(n_8_0_2422));
   OAI21_X1 i_8_0_2275 (.A(n_8_0_2424), .B1(n_8_0_5613), .B2(in_data[20]), 
      .ZN(n_8_0_2423));
   OAI211_X1 i_8_0_2276 (.A(n_8_0_5613), .B(n_8_0_2425), .C1(n_8_0_6995), 
      .C2(n_8_0_5619), .ZN(n_8_0_2424));
   NAND2_X1 i_8_0_2277 (.A1(in_data[24]), .A2(n_8_0_5619), .ZN(n_8_0_2425));
   NAND2_X1 i_8_0_2278 (.A1(n_8_0_5597), .A2(in_data[16]), .ZN(n_8_0_2426));
   NAND2_X1 i_8_0_2279 (.A1(in_data[8]), .A2(n_8_0_5600), .ZN(n_8_0_2427));
   AOI21_X1 i_8_0_2280 (.A(n_8_0_5611), .B1(n_8_0_5610), .B2(n_8_0_6729), 
      .ZN(n_8_0_2428));
   OAI21_X1 i_8_0_2281 (.A(n_8_0_2429), .B1(n_8_0_2431), .B2(n_8_0_6988), 
      .ZN(n_85));
   OAI211_X1 i_8_0_2282 (.A(n_8_0_2431), .B(n_8_0_2430), .C1(n_8_0_5657), 
      .C2(n_8_0_2432), .ZN(n_8_0_2429));
   NAND2_X1 i_8_0_2283 (.A1(n_8_0_6989), .A2(n_8_0_5657), .ZN(n_8_0_2430));
   AOI21_X1 i_8_0_2284 (.A(n_8_0_5651), .B1(n_8_0_5650), .B2(n_8_0_6729), 
      .ZN(n_8_0_2431));
   OAI22_X1 i_8_0_2285 (.A1(n_8_0_2433), .A2(n_8_0_2434), .B1(n_8_0_5654), 
      .B2(n_8_0_6990), .ZN(n_8_0_2432));
   NOR2_X1 i_8_0_2286 (.A1(n_8_0_2435), .A2(n_8_0_5631), .ZN(n_8_0_2433));
   OAI21_X1 i_8_0_2287 (.A(n_8_0_5654), .B1(n_8_0_5632), .B2(in_data[12]), 
      .ZN(n_8_0_2434));
   MUX2_X1 i_8_0_2288 (.A(n_8_0_2436), .B(in_data[16]), .S(n_8_0_5628), .Z(
      n_8_0_2435));
   OAI22_X1 i_8_0_2289 (.A1(n_8_0_2437), .A2(n_8_0_2438), .B1(n_8_0_5639), 
      .B2(n_8_0_6993), .ZN(n_8_0_2436));
   OAI21_X1 i_8_0_2290 (.A(n_8_0_5639), .B1(n_8_0_5643), .B2(in_data[24]), 
      .ZN(n_8_0_2437));
   NOR2_X1 i_8_0_2291 (.A1(in_data[28]), .A2(n_8_0_5644), .ZN(n_8_0_2438));
   NOR2_X1 i_8_0_2292 (.A1(n_8_0_2449), .A2(n_8_0_2439), .ZN(n_86));
   AOI21_X1 i_8_0_2293 (.A(n_8_0_2440), .B1(n_8_0_2441), .B2(n_8_0_5675), 
      .ZN(n_8_0_2439));
   OAI21_X1 i_8_0_2294 (.A(n_8_0_2450), .B1(n_8_0_5675), .B2(n_8_0_6989), 
      .ZN(n_8_0_2440));
   OAI21_X1 i_8_0_2295 (.A(n_8_0_2442), .B1(n_8_0_5679), .B2(n_8_0_6990), 
      .ZN(n_8_0_2441));
   OAI211_X1 i_8_0_2296 (.A(n_8_0_5679), .B(n_8_0_2443), .C1(n_8_0_2444), 
      .C2(n_8_0_5688), .ZN(n_8_0_2442));
   NAND2_X1 i_8_0_2297 (.A1(n_8_0_5688), .A2(n_8_0_6991), .ZN(n_8_0_2443));
   AOI21_X1 i_8_0_2298 (.A(n_8_0_2445), .B1(n_8_0_2446), .B2(n_8_0_5684), 
      .ZN(n_8_0_2444));
   NOR2_X1 i_8_0_2299 (.A1(n_8_0_5684), .A2(in_data[16]), .ZN(n_8_0_2445));
   OAI22_X1 i_8_0_2300 (.A1(n_8_0_2447), .A2(n_8_0_2448), .B1(n_8_0_5662), 
      .B2(in_data[20]), .ZN(n_8_0_2446));
   OAI21_X1 i_8_0_2301 (.A(n_8_0_5662), .B1(n_8_0_5666), .B2(n_8_0_6995), 
      .ZN(n_8_0_2447));
   AND2_X1 i_8_0_2302 (.A1(in_data[24]), .A2(n_8_0_5666), .ZN(n_8_0_2448));
   NOR2_X1 i_8_0_2303 (.A1(n_8_0_2450), .A2(in_data[0]), .ZN(n_8_0_2449));
   AOI21_X1 i_8_0_2304 (.A(n_8_0_5672), .B1(n_8_0_5671), .B2(n_8_0_6729), 
      .ZN(n_8_0_2450));
   OAI22_X1 i_8_0_2305 (.A1(n_8_0_2452), .A2(n_8_0_2451), .B1(n_8_0_6988), 
      .B2(n_8_0_2461), .ZN(n_87));
   OAI21_X1 i_8_0_2306 (.A(n_8_0_2461), .B1(n_8_0_5720), .B2(in_data[4]), 
      .ZN(n_8_0_2451));
   AOI211_X1 i_8_0_2307 (.A(n_8_0_5719), .B(n_8_0_2453), .C1(n_8_0_5699), 
      .C2(in_data[8]), .ZN(n_8_0_2452));
   AOI211_X1 i_8_0_2308 (.A(n_8_0_5699), .B(n_8_0_2454), .C1(n_8_0_2455), 
      .C2(n_8_0_5725), .ZN(n_8_0_2453));
   NOR2_X1 i_8_0_2309 (.A1(n_8_0_5725), .A2(in_data[12]), .ZN(n_8_0_2454));
   INV_X1 i_8_0_2310 (.A(n_8_0_2456), .ZN(n_8_0_2455));
   AOI21_X1 i_8_0_2311 (.A(n_8_0_2457), .B1(n_8_0_5693), .B2(n_8_0_6992), 
      .ZN(n_8_0_2456));
   AOI211_X1 i_8_0_2312 (.A(n_8_0_5693), .B(n_8_0_2458), .C1(n_8_0_2459), 
      .C2(n_8_0_5704), .ZN(n_8_0_2457));
   NOR2_X1 i_8_0_2313 (.A1(n_8_0_6993), .A2(n_8_0_5704), .ZN(n_8_0_2458));
   OAI21_X1 i_8_0_2314 (.A(n_8_0_2460), .B1(n_8_0_5708), .B2(n_8_0_6994), 
      .ZN(n_8_0_2459));
   NAND2_X1 i_8_0_2315 (.A1(n_8_0_5708), .A2(in_data[28]), .ZN(n_8_0_2460));
   OAI21_X1 i_8_0_2316 (.A(n_8_0_5713), .B1(n_8_0_6729), .B2(n_8_0_5714), 
      .ZN(n_8_0_2461));
   AOI21_X1 i_8_0_2317 (.A(n_8_0_2462), .B1(n_8_0_5735), .B2(n_8_0_6988), 
      .ZN(n_88));
   AOI21_X1 i_8_0_2318 (.A(n_8_0_5735), .B1(n_8_0_2464), .B2(n_8_0_2463), 
      .ZN(n_8_0_2462));
   NAND2_X1 i_8_0_2319 (.A1(n_8_0_5749), .A2(n_8_0_6989), .ZN(n_8_0_2463));
   OAI21_X1 i_8_0_2320 (.A(n_8_0_2465), .B1(n_8_0_2466), .B2(n_8_0_5746), 
      .ZN(n_8_0_2464));
   AOI21_X1 i_8_0_2321 (.A(n_8_0_5749), .B1(n_8_0_5746), .B2(in_data[8]), 
      .ZN(n_8_0_2465));
   INV_X1 i_8_0_2322 (.A(n_8_0_2467), .ZN(n_8_0_2466));
   MUX2_X1 i_8_0_2323 (.A(n_8_0_2468), .B(in_data[12]), .S(n_8_0_5742), .Z(
      n_8_0_2467));
   AOI21_X1 i_8_0_2324 (.A(n_8_0_2469), .B1(n_8_0_5738), .B2(n_8_0_6992), 
      .ZN(n_8_0_2468));
   AOI211_X1 i_8_0_2325 (.A(n_8_0_5738), .B(n_8_0_2470), .C1(n_8_0_2471), 
      .C2(n_8_0_5733), .ZN(n_8_0_2469));
   NOR2_X1 i_8_0_2326 (.A1(n_8_0_6993), .A2(n_8_0_5733), .ZN(n_8_0_2470));
   OAI21_X1 i_8_0_2327 (.A(n_8_0_2472), .B1(n_8_0_5731), .B2(n_8_0_6994), 
      .ZN(n_8_0_2471));
   NAND2_X1 i_8_0_2328 (.A1(n_8_0_5731), .A2(in_data[28]), .ZN(n_8_0_2472));
   MUX2_X1 i_8_0_2329 (.A(in_data[0]), .B(n_8_0_2473), .S(n_8_0_2483), .Z(n_89));
   OAI21_X1 i_8_0_2330 (.A(n_8_0_2474), .B1(n_8_0_5765), .B2(n_8_0_6989), 
      .ZN(n_8_0_2473));
   NAND2_X1 i_8_0_2331 (.A1(n_8_0_5765), .A2(n_8_0_2475), .ZN(n_8_0_2474));
   OAI21_X1 i_8_0_2332 (.A(n_8_0_2476), .B1(n_8_0_5772), .B2(n_8_0_6990), 
      .ZN(n_8_0_2475));
   NAND2_X1 i_8_0_2333 (.A1(n_8_0_5772), .A2(n_8_0_2477), .ZN(n_8_0_2476));
   OAI221_X1 i_8_0_2334 (.A(n_8_0_2481), .B1(n_8_0_2478), .B2(n_8_0_5776), 
      .C1(n_8_0_5780), .C2(n_8_0_6991), .ZN(n_8_0_2477));
   INV_X1 i_8_0_2335 (.A(n_8_0_2479), .ZN(n_8_0_2478));
   OAI21_X1 i_8_0_2336 (.A(n_8_0_2480), .B1(n_8_0_5755), .B2(n_8_0_6994), 
      .ZN(n_8_0_2479));
   NAND2_X1 i_8_0_2337 (.A1(n_8_0_5755), .A2(in_data[28]), .ZN(n_8_0_2480));
   OAI211_X1 i_8_0_2338 (.A(n_8_0_5780), .B(n_8_0_2482), .C1(in_data[16]), 
      .C2(n_8_0_5784), .ZN(n_8_0_2481));
   OAI21_X1 i_8_0_2339 (.A(n_8_0_5784), .B1(n_8_0_5777), .B2(n_8_0_6993), 
      .ZN(n_8_0_2482));
   OAI21_X1 i_8_0_2340 (.A(n_8_0_2484), .B1(n_8_0_5762), .B2(n_8_0_6729), 
      .ZN(n_8_0_2483));
   OAI21_X1 i_8_0_2341 (.A(n_8_0_482), .B1(n_8_0_6730), .B2(n_8_0_5761), 
      .ZN(n_8_0_2484));
   AOI21_X1 i_8_0_2342 (.A(n_8_0_2485), .B1(n_8_0_2495), .B2(n_8_0_6988), 
      .ZN(n_90));
   NOR2_X1 i_8_0_2343 (.A1(n_8_0_2495), .A2(n_8_0_2486), .ZN(n_8_0_2485));
   AOI22_X1 i_8_0_2344 (.A1(n_8_0_2487), .A2(n_8_0_2488), .B1(n_8_0_5820), 
      .B2(n_8_0_6989), .ZN(n_8_0_2486));
   AOI21_X1 i_8_0_2345 (.A(n_8_0_5820), .B1(n_8_0_5794), .B2(in_data[8]), 
      .ZN(n_8_0_2487));
   OAI21_X1 i_8_0_2346 (.A(n_8_0_2489), .B1(n_8_0_2490), .B2(n_8_0_5797), 
      .ZN(n_8_0_2488));
   AOI21_X1 i_8_0_2347 (.A(n_8_0_5794), .B1(n_8_0_5797), .B2(n_8_0_6991), 
      .ZN(n_8_0_2489));
   AOI22_X1 i_8_0_2348 (.A1(n_8_0_2491), .A2(n_8_0_2492), .B1(n_8_0_5791), 
      .B2(n_8_0_6992), .ZN(n_8_0_2490));
   AOI21_X1 i_8_0_2349 (.A(n_8_0_5791), .B1(n_8_0_5811), .B2(in_data[20]), 
      .ZN(n_8_0_2491));
   NAND2_X1 i_8_0_2350 (.A1(n_8_0_5810), .A2(n_8_0_2493), .ZN(n_8_0_2492));
   OAI21_X1 i_8_0_2351 (.A(n_8_0_2494), .B1(n_8_0_5816), .B2(n_8_0_6995), 
      .ZN(n_8_0_2493));
   NAND2_X1 i_8_0_2352 (.A1(in_data[24]), .A2(n_8_0_5816), .ZN(n_8_0_2494));
   OAI21_X1 i_8_0_2353 (.A(n_8_0_5808), .B1(n_8_0_5807), .B2(n_8_0_6730), 
      .ZN(n_8_0_2495));
   OAI21_X1 i_8_0_2354 (.A(n_8_0_2496), .B1(n_8_0_2507), .B2(n_8_0_6988), 
      .ZN(n_91));
   NAND3_X1 i_8_0_2355 (.A1(n_8_0_2498), .A2(n_8_0_2497), .A3(n_8_0_2507), 
      .ZN(n_8_0_2496));
   NAND2_X1 i_8_0_2356 (.A1(n_8_0_5825), .A2(n_8_0_6989), .ZN(n_8_0_2497));
   OAI21_X1 i_8_0_2357 (.A(n_8_0_2499), .B1(n_8_0_2500), .B2(n_8_0_5829), 
      .ZN(n_8_0_2498));
   AOI21_X1 i_8_0_2358 (.A(n_8_0_5825), .B1(n_8_0_5829), .B2(in_data[8]), 
      .ZN(n_8_0_2499));
   INV_X1 i_8_0_2359 (.A(n_8_0_2501), .ZN(n_8_0_2500));
   AOI21_X1 i_8_0_2360 (.A(n_8_0_2502), .B1(n_8_0_5832), .B2(n_8_0_6991), 
      .ZN(n_8_0_2501));
   AOI211_X1 i_8_0_2361 (.A(n_8_0_5832), .B(n_8_0_2503), .C1(n_8_0_2504), 
      .C2(n_8_0_5855), .ZN(n_8_0_2502));
   NOR2_X1 i_8_0_2362 (.A1(n_8_0_6992), .A2(n_8_0_5855), .ZN(n_8_0_2503));
   MUX2_X1 i_8_0_2363 (.A(n_8_0_2505), .B(in_data[20]), .S(n_8_0_5843), .Z(
      n_8_0_2504));
   OAI21_X1 i_8_0_2364 (.A(n_8_0_2506), .B1(n_8_0_5847), .B2(n_8_0_6994), 
      .ZN(n_8_0_2505));
   NAND2_X1 i_8_0_2365 (.A1(n_8_0_5847), .A2(in_data[28]), .ZN(n_8_0_2506));
   AOI21_X1 i_8_0_2366 (.A(n_8_0_5840), .B1(n_8_0_5839), .B2(n_8_0_6729), 
      .ZN(n_8_0_2507));
   OAI21_X1 i_8_0_2367 (.A(n_8_0_2508), .B1(n_8_0_2519), .B2(n_8_0_6988), 
      .ZN(n_92));
   OAI211_X1 i_8_0_2368 (.A(n_8_0_2519), .B(n_8_0_2509), .C1(in_data[4]), 
      .C2(n_8_0_5872), .ZN(n_8_0_2508));
   OAI211_X1 i_8_0_2369 (.A(n_8_0_5872), .B(n_8_0_2510), .C1(n_8_0_2511), 
      .C2(n_8_0_5866), .ZN(n_8_0_2509));
   NAND2_X1 i_8_0_2370 (.A1(in_data[8]), .A2(n_8_0_5866), .ZN(n_8_0_2510));
   INV_X1 i_8_0_2371 (.A(n_8_0_2512), .ZN(n_8_0_2511));
   OAI21_X1 i_8_0_2372 (.A(n_8_0_2513), .B1(n_8_0_5869), .B2(n_8_0_6991), 
      .ZN(n_8_0_2512));
   NAND2_X1 i_8_0_2373 (.A1(n_8_0_5869), .A2(n_8_0_2514), .ZN(n_8_0_2513));
   MUX2_X1 i_8_0_2374 (.A(n_8_0_2515), .B(in_data[16]), .S(n_8_0_5862), .Z(
      n_8_0_2514));
   OAI21_X1 i_8_0_2375 (.A(n_8_0_2516), .B1(n_8_0_5879), .B2(n_8_0_6993), 
      .ZN(n_8_0_2515));
   NAND2_X1 i_8_0_2376 (.A1(n_8_0_5879), .A2(n_8_0_2517), .ZN(n_8_0_2516));
   OAI21_X1 i_8_0_2377 (.A(n_8_0_2518), .B1(n_8_0_5875), .B2(n_8_0_6995), 
      .ZN(n_8_0_2517));
   NAND2_X1 i_8_0_2378 (.A1(in_data[24]), .A2(n_8_0_5875), .ZN(n_8_0_2518));
   AOI21_X1 i_8_0_2379 (.A(n_8_0_5877), .B1(n_8_0_5878), .B2(n_8_0_6729), 
      .ZN(n_8_0_2519));
   MUX2_X1 i_8_0_2380 (.A(in_data[0]), .B(n_8_0_2520), .S(n_8_0_2529), .Z(n_93));
   AOI21_X1 i_8_0_2381 (.A(n_8_0_2521), .B1(n_8_0_5888), .B2(n_8_0_6989), 
      .ZN(n_8_0_2520));
   AOI221_X1 i_8_0_2382 (.A(n_8_0_5888), .B1(n_8_0_5919), .B2(in_data[8]), 
      .C1(n_8_0_2522), .C2(n_8_0_2523), .ZN(n_8_0_2521));
   AOI21_X1 i_8_0_2383 (.A(n_8_0_5919), .B1(n_8_0_5895), .B2(n_8_0_6991), 
      .ZN(n_8_0_2522));
   OAI21_X1 i_8_0_2384 (.A(n_8_0_2526), .B1(n_8_0_2524), .B2(n_8_0_5915), 
      .ZN(n_8_0_2523));
   OAI21_X1 i_8_0_2385 (.A(n_8_0_2525), .B1(n_8_0_2527), .B2(n_8_0_5903), 
      .ZN(n_8_0_2524));
   NAND2_X1 i_8_0_2386 (.A1(n_8_0_5903), .A2(n_8_0_6993), .ZN(n_8_0_2525));
   AOI21_X1 i_8_0_2387 (.A(n_8_0_5895), .B1(n_8_0_5915), .B2(in_data[16]), 
      .ZN(n_8_0_2526));
   OAI21_X1 i_8_0_2388 (.A(n_8_0_2528), .B1(n_8_0_5898), .B2(n_8_0_6994), 
      .ZN(n_8_0_2527));
   NAND2_X1 i_8_0_2389 (.A1(n_8_0_5898), .A2(in_data[28]), .ZN(n_8_0_2528));
   AOI21_X1 i_8_0_2390 (.A(n_8_0_5912), .B1(n_8_0_5911), .B2(n_8_0_6729), 
      .ZN(n_8_0_2529));
   OAI21_X1 i_8_0_2391 (.A(n_8_0_2530), .B1(n_8_0_2540), .B2(n_8_0_6988), 
      .ZN(n_94));
   NAND2_X1 i_8_0_2392 (.A1(n_8_0_2531), .A2(n_8_0_2540), .ZN(n_8_0_2530));
   AOI21_X1 i_8_0_2393 (.A(n_8_0_2532), .B1(n_8_0_5933), .B2(n_8_0_6989), 
      .ZN(n_8_0_2531));
   AOI211_X1 i_8_0_2394 (.A(n_8_0_5933), .B(n_8_0_2533), .C1(n_8_0_2534), 
      .C2(n_8_0_5955), .ZN(n_8_0_2532));
   NOR2_X1 i_8_0_2395 (.A1(n_8_0_5955), .A2(n_8_0_6990), .ZN(n_8_0_2533));
   MUX2_X1 i_8_0_2396 (.A(n_8_0_2535), .B(in_data[12]), .S(n_8_0_5925), .Z(
      n_8_0_2534));
   OAI22_X1 i_8_0_2397 (.A1(n_8_0_2536), .A2(n_8_0_2537), .B1(n_8_0_5930), 
      .B2(n_8_0_6992), .ZN(n_8_0_2535));
   OAI21_X1 i_8_0_2398 (.A(n_8_0_5930), .B1(n_8_0_2538), .B2(n_8_0_5945), 
      .ZN(n_8_0_2536));
   AND2_X1 i_8_0_2399 (.A1(n_8_0_5945), .A2(n_8_0_6993), .ZN(n_8_0_2537));
   OAI21_X1 i_8_0_2400 (.A(n_8_0_2539), .B1(n_8_0_5958), .B2(n_8_0_6994), 
      .ZN(n_8_0_2538));
   NAND2_X1 i_8_0_2401 (.A1(n_8_0_5958), .A2(in_data[28]), .ZN(n_8_0_2539));
   AOI21_X1 i_8_0_2402 (.A(n_8_0_5949), .B1(n_8_0_5950), .B2(n_8_0_6729), 
      .ZN(n_8_0_2540));
   NAND2_X1 i_8_0_2406 (.A1(n_8_0_6989), .A2(n_8_0_5971), .ZN(n_8_0_2543));
   AOI21_X1 i_8_0_2409 (.A(n_8_0_5993), .B1(n_8_0_6001), .B2(in_data[16]), 
      .ZN(n_8_0_2546));
   OAI211_X1 i_8_0_2410 (.A(n_8_0_6002), .B(n_8_0_2548), .C1(n_8_0_2549), 
      .C2(n_8_0_5985), .ZN(n_8_0_2547));
   NAND2_X1 i_8_0_2411 (.A1(n_8_0_5985), .A2(n_8_0_6993), .ZN(n_8_0_2548));
   OAI21_X1 i_8_0_2412 (.A(n_8_0_2550), .B1(n_8_0_5977), .B2(n_8_0_6994), 
      .ZN(n_8_0_2549));
   NAND2_X1 i_8_0_2413 (.A1(n_8_0_5977), .A2(in_data[28]), .ZN(n_8_0_2550));
   MUX2_X1 i_8_0_2414 (.A(in_data[0]), .B(n_8_0_2551), .S(n_8_0_2560), .Z(n_95));
   AOI21_X1 i_8_0_2415 (.A(n_8_0_2552), .B1(n_8_0_6011), .B2(n_8_0_6989), 
      .ZN(n_8_0_2551));
   AOI211_X1 i_8_0_2416 (.A(n_8_0_6011), .B(n_8_0_2553), .C1(in_data[8]), 
      .C2(n_8_0_6013), .ZN(n_8_0_2552));
   AOI211_X1 i_8_0_2417 (.A(n_8_0_6013), .B(n_8_0_2554), .C1(n_8_0_6991), 
      .C2(n_8_0_6014), .ZN(n_8_0_2553));
   AOI211_X1 i_8_0_2418 (.A(n_8_0_6014), .B(n_8_0_2555), .C1(n_8_0_6012), 
      .C2(in_data[16]), .ZN(n_8_0_2554));
   AOI211_X1 i_8_0_2419 (.A(n_8_0_6012), .B(n_8_0_2556), .C1(n_8_0_2557), 
      .C2(n_8_0_6018), .ZN(n_8_0_2555));
   NOR2_X1 i_8_0_2420 (.A1(n_8_0_6018), .A2(in_data[20]), .ZN(n_8_0_2556));
   INV_X1 i_8_0_2421 (.A(n_8_0_2558), .ZN(n_8_0_2557));
   OAI21_X1 i_8_0_2422 (.A(n_8_0_2559), .B1(n_8_0_6022), .B2(n_8_0_6994), 
      .ZN(n_8_0_2558));
   NAND2_X1 i_8_0_2423 (.A1(in_data[28]), .A2(n_8_0_6022), .ZN(n_8_0_2559));
   OAI21_X1 i_8_0_2424 (.A(n_8_0_6020), .B1(n_8_0_6729), .B2(n_8_0_6021), 
      .ZN(n_8_0_2560));
   AOI21_X1 i_8_0_2425 (.A(n_8_0_2561), .B1(n_8_0_2563), .B2(n_8_0_6988), 
      .ZN(n_96));
   NOR2_X1 i_8_0_2426 (.A1(n_8_0_2563), .A2(n_8_0_2562), .ZN(n_8_0_2561));
   AOI21_X1 i_8_0_2427 (.A(n_8_0_2564), .B1(n_8_0_6032), .B2(n_8_0_6989), 
      .ZN(n_8_0_2562));
   OAI21_X1 i_8_0_2428 (.A(n_8_0_6039), .B1(n_8_0_6038), .B2(n_8_0_6730), 
      .ZN(n_8_0_2563));
   AOI211_X1 i_8_0_2429 (.A(n_8_0_6032), .B(n_8_0_2565), .C1(in_data[8]), 
      .C2(n_8_0_6055), .ZN(n_8_0_2564));
   AOI221_X1 i_8_0_2430 (.A(n_8_0_6055), .B1(n_8_0_2566), .B2(n_8_0_2567), 
      .C1(n_8_0_6991), .C2(n_8_0_6028), .ZN(n_8_0_2565));
   AOI21_X1 i_8_0_2431 (.A(n_8_0_6028), .B1(n_8_0_2568), .B2(n_8_0_6060), 
      .ZN(n_8_0_2566));
   NAND2_X1 i_8_0_2432 (.A1(n_8_0_6061), .A2(in_data[16]), .ZN(n_8_0_2567));
   AOI21_X1 i_8_0_2433 (.A(n_8_0_2569), .B1(n_8_0_6043), .B2(n_8_0_6993), 
      .ZN(n_8_0_2568));
   AOI211_X1 i_8_0_2434 (.A(n_8_0_6043), .B(n_8_0_2570), .C1(in_data[28]), 
      .C2(n_8_0_6047), .ZN(n_8_0_2569));
   NOR2_X1 i_8_0_2435 (.A1(n_8_0_6994), .A2(n_8_0_6047), .ZN(n_8_0_2570));
   OAI21_X1 i_8_0_2436 (.A(n_8_0_2571), .B1(n_8_0_2582), .B2(n_8_0_6988), 
      .ZN(n_97));
   OAI211_X1 i_8_0_2437 (.A(n_8_0_2582), .B(n_8_0_2572), .C1(in_data[4]), 
      .C2(n_8_0_6083), .ZN(n_8_0_2571));
   OAI211_X1 i_8_0_2438 (.A(n_8_0_6083), .B(n_8_0_2573), .C1(n_8_0_2574), 
      .C2(n_8_0_6094), .ZN(n_8_0_2572));
   NAND2_X1 i_8_0_2439 (.A1(in_data[8]), .A2(n_8_0_6094), .ZN(n_8_0_2573));
   INV_X1 i_8_0_2440 (.A(n_8_0_2575), .ZN(n_8_0_2574));
   OAI21_X1 i_8_0_2441 (.A(n_8_0_2576), .B1(n_8_0_6089), .B2(n_8_0_6991), 
      .ZN(n_8_0_2575));
   NAND2_X1 i_8_0_2442 (.A1(n_8_0_6089), .A2(n_8_0_2577), .ZN(n_8_0_2576));
   OAI21_X1 i_8_0_2443 (.A(n_8_0_2578), .B1(n_8_0_6099), .B2(n_8_0_6992), 
      .ZN(n_8_0_2577));
   OAI211_X1 i_8_0_2444 (.A(n_8_0_2579), .B(n_8_0_6099), .C1(n_8_0_6067), 
      .C2(n_8_0_2580), .ZN(n_8_0_2578));
   NAND2_X1 i_8_0_2445 (.A1(n_8_0_6067), .A2(n_8_0_6993), .ZN(n_8_0_2579));
   OAI21_X1 i_8_0_2446 (.A(n_8_0_2581), .B1(n_8_0_6072), .B2(n_8_0_6994), 
      .ZN(n_8_0_2580));
   NAND2_X1 i_8_0_2447 (.A1(n_8_0_6072), .A2(in_data[28]), .ZN(n_8_0_2581));
   AOI21_X1 i_8_0_2448 (.A(n_8_0_6077), .B1(n_8_0_6078), .B2(n_8_0_6729), 
      .ZN(n_8_0_2582));
   OAI21_X1 i_8_0_2449 (.A(n_8_0_2583), .B1(n_8_0_6115), .B2(n_8_0_6988), 
      .ZN(n_98));
   NAND2_X1 i_8_0_2450 (.A1(n_8_0_2584), .A2(n_8_0_6115), .ZN(n_8_0_2583));
   MUX2_X1 i_8_0_2451 (.A(in_data[4]), .B(n_8_0_2585), .S(n_8_0_6120), .Z(
      n_8_0_2584));
   OAI21_X1 i_8_0_2452 (.A(n_8_0_2586), .B1(n_8_0_6132), .B2(n_8_0_6990), 
      .ZN(n_8_0_2585));
   OAI21_X1 i_8_0_2453 (.A(n_8_0_2587), .B1(n_8_0_6110), .B2(in_data[12]), 
      .ZN(n_8_0_2586));
   AOI21_X1 i_8_0_2454 (.A(n_8_0_6133), .B1(n_8_0_6110), .B2(n_8_0_2588), 
      .ZN(n_8_0_2587));
   INV_X1 i_8_0_2455 (.A(n_8_0_2589), .ZN(n_8_0_2588));
   AOI22_X1 i_8_0_2456 (.A1(n_8_0_2590), .A2(n_8_0_2591), .B1(n_8_0_6105), 
      .B2(n_8_0_6992), .ZN(n_8_0_2589));
   AOI21_X1 i_8_0_2457 (.A(n_8_0_6105), .B1(n_8_0_6129), .B2(in_data[20]), 
      .ZN(n_8_0_2590));
   NAND2_X1 i_8_0_2458 (.A1(n_8_0_6128), .A2(n_8_0_2592), .ZN(n_8_0_2591));
   OAI21_X1 i_8_0_2459 (.A(n_8_0_2593), .B1(n_8_0_6124), .B2(n_8_0_6994), 
      .ZN(n_8_0_2592));
   NAND2_X1 i_8_0_2460 (.A1(n_8_0_6124), .A2(in_data[28]), .ZN(n_8_0_2593));
   OAI21_X1 i_8_0_2461 (.A(n_8_0_2594), .B1(n_8_0_6155), .B2(n_8_0_6988), 
      .ZN(n_99));
   OAI211_X1 i_8_0_2462 (.A(n_8_0_6155), .B(n_8_0_2595), .C1(n_8_0_2596), 
      .C2(n_8_0_2597), .ZN(n_8_0_2594));
   NAND2_X1 i_8_0_2463 (.A1(n_8_0_6152), .A2(n_8_0_6989), .ZN(n_8_0_2595));
   AOI211_X1 i_8_0_2464 (.A(n_8_0_6163), .B(n_8_0_2599), .C1(n_8_0_6991), 
      .C2(n_8_0_6167), .ZN(n_8_0_2596));
   INV_X1 i_8_0_2465 (.A(n_8_0_2598), .ZN(n_8_0_2597));
   AOI21_X1 i_8_0_2466 (.A(n_8_0_6152), .B1(n_8_0_6163), .B2(in_data[8]), 
      .ZN(n_8_0_2598));
   AOI211_X1 i_8_0_2467 (.A(n_8_0_6167), .B(n_8_0_2601), .C1(n_8_0_2600), 
      .C2(n_8_0_2602), .ZN(n_8_0_2599));
   AOI21_X1 i_8_0_2468 (.A(n_8_0_6158), .B1(n_8_0_6148), .B2(n_8_0_2603), 
      .ZN(n_8_0_2600));
   AND2_X1 i_8_0_2469 (.A1(in_data[16]), .A2(n_8_0_6158), .ZN(n_8_0_2601));
   OR2_X1 i_8_0_2470 (.A1(n_8_0_6148), .A2(in_data[20]), .ZN(n_8_0_2602));
   OAI21_X1 i_8_0_2471 (.A(n_8_0_2604), .B1(n_8_0_6144), .B2(in_data[28]), 
      .ZN(n_8_0_2603));
   NAND2_X1 i_8_0_2472 (.A1(n_8_0_6144), .A2(n_8_0_6994), .ZN(n_8_0_2604));
   OAI21_X1 i_8_0_2473 (.A(n_8_0_2605), .B1(n_8_0_6199), .B2(n_8_0_6988), 
      .ZN(n_100));
   OAI211_X1 i_8_0_2474 (.A(n_8_0_6199), .B(n_8_0_2606), .C1(n_8_0_2607), 
      .C2(n_8_0_6193), .ZN(n_8_0_2605));
   NAND2_X1 i_8_0_2475 (.A1(n_8_0_6989), .A2(n_8_0_6193), .ZN(n_8_0_2606));
   MUX2_X1 i_8_0_2476 (.A(n_8_0_2608), .B(in_data[8]), .S(n_8_0_6207), .Z(
      n_8_0_2607));
   AOI21_X1 i_8_0_2477 (.A(n_8_0_2609), .B1(n_8_0_6186), .B2(n_8_0_6991), 
      .ZN(n_8_0_2608));
   AOI211_X1 i_8_0_2478 (.A(n_8_0_6186), .B(n_8_0_2610), .C1(n_8_0_2611), 
      .C2(n_8_0_6212), .ZN(n_8_0_2609));
   NOR2_X1 i_8_0_2479 (.A1(n_8_0_6992), .A2(n_8_0_6212), .ZN(n_8_0_2610));
   OAI21_X1 i_8_0_2480 (.A(n_8_0_2612), .B1(n_8_0_6179), .B2(n_8_0_6993), 
      .ZN(n_8_0_2611));
   OAI211_X1 i_8_0_2481 (.A(n_8_0_6179), .B(n_8_0_2613), .C1(in_data[24]), 
      .C2(n_8_0_6203), .ZN(n_8_0_2612));
   NAND2_X1 i_8_0_2482 (.A1(n_8_0_6995), .A2(n_8_0_6203), .ZN(n_8_0_2613));
   OAI21_X1 i_8_0_2483 (.A(n_8_0_2614), .B1(n_8_0_2616), .B2(n_8_0_6988), 
      .ZN(n_101));
   OAI211_X1 i_8_0_2484 (.A(n_8_0_2615), .B(n_8_0_2616), .C1(n_8_0_2617), 
      .C2(n_8_0_6223), .ZN(n_8_0_2614));
   NAND2_X1 i_8_0_2485 (.A1(n_8_0_6223), .A2(n_8_0_6989), .ZN(n_8_0_2615));
   OAI21_X1 i_8_0_2486 (.A(n_8_0_6234), .B1(n_8_0_6729), .B2(n_8_0_6235), 
      .ZN(n_8_0_2616));
   AOI21_X1 i_8_0_2487 (.A(n_8_0_2618), .B1(n_8_0_6227), .B2(n_8_0_6990), 
      .ZN(n_8_0_2617));
   NOR2_X1 i_8_0_2488 (.A1(n_8_0_6227), .A2(n_8_0_2619), .ZN(n_8_0_2618));
   AOI22_X1 i_8_0_2489 (.A1(n_8_0_2620), .A2(n_8_0_2621), .B1(n_8_0_6241), 
      .B2(n_8_0_6991), .ZN(n_8_0_2619));
   AOI21_X1 i_8_0_2490 (.A(n_8_0_6241), .B1(n_8_0_6254), .B2(in_data[16]), 
      .ZN(n_8_0_2620));
   OR2_X1 i_8_0_2491 (.A1(n_8_0_2622), .A2(n_8_0_6254), .ZN(n_8_0_2621));
   AOI21_X1 i_8_0_2492 (.A(n_8_0_2623), .B1(n_8_0_2624), .B2(n_8_0_6229), 
      .ZN(n_8_0_2622));
   NOR2_X1 i_8_0_2493 (.A1(n_8_0_6993), .A2(n_8_0_6229), .ZN(n_8_0_2623));
   OAI21_X1 i_8_0_2494 (.A(n_8_0_2625), .B1(n_8_0_6239), .B2(n_8_0_6994), 
      .ZN(n_8_0_2624));
   NAND2_X1 i_8_0_2495 (.A1(n_8_0_6239), .A2(in_data[28]), .ZN(n_8_0_2625));
   OAI22_X1 i_8_0_2496 (.A1(n_8_0_2627), .A2(n_8_0_2626), .B1(n_8_0_6988), 
      .B2(n_8_0_6276), .ZN(n_102));
   OAI21_X1 i_8_0_2497 (.A(n_8_0_6276), .B1(n_8_0_6289), .B2(in_data[4]), 
      .ZN(n_8_0_2626));
   AOI21_X1 i_8_0_2498 (.A(n_8_0_2628), .B1(n_8_0_2629), .B2(n_8_0_6295), 
      .ZN(n_8_0_2627));
   OAI21_X1 i_8_0_2499 (.A(n_8_0_6289), .B1(n_8_0_6295), .B2(n_8_0_6990), 
      .ZN(n_8_0_2628));
   MUX2_X1 i_8_0_2500 (.A(in_data[12]), .B(n_8_0_2630), .S(n_8_0_6272), .Z(
      n_8_0_2629));
   MUX2_X1 i_8_0_2501 (.A(in_data[16]), .B(n_8_0_2631), .S(n_8_0_6302), .Z(
      n_8_0_2630));
   OAI21_X1 i_8_0_2502 (.A(n_8_0_2632), .B1(n_8_0_6280), .B2(n_8_0_6993), 
      .ZN(n_8_0_2631));
   NAND2_X1 i_8_0_2503 (.A1(n_8_0_6280), .A2(n_8_0_2633), .ZN(n_8_0_2632));
   OAI21_X1 i_8_0_2504 (.A(n_8_0_2634), .B1(n_8_0_6263), .B2(n_8_0_6994), 
      .ZN(n_8_0_2633));
   NAND2_X1 i_8_0_2505 (.A1(n_8_0_6263), .A2(in_data[28]), .ZN(n_8_0_2634));
   OAI22_X1 i_8_0_2506 (.A1(n_8_0_2636), .A2(n_8_0_2635), .B1(n_8_0_6988), 
      .B2(n_8_0_2637), .ZN(n_103));
   OAI21_X1 i_8_0_2507 (.A(n_8_0_2637), .B1(n_8_0_6309), .B2(in_data[4]), 
      .ZN(n_8_0_2635));
   NOR2_X1 i_8_0_2508 (.A1(n_8_0_6310), .A2(n_8_0_2638), .ZN(n_8_0_2636));
   OAI21_X1 i_8_0_2509 (.A(n_8_0_6316), .B1(n_8_0_6729), .B2(n_8_0_6317), 
      .ZN(n_8_0_2637));
   OAI21_X1 i_8_0_2510 (.A(n_8_0_2639), .B1(n_8_0_6312), .B2(n_8_0_6990), 
      .ZN(n_8_0_2638));
   OAI211_X1 i_8_0_2511 (.A(n_8_0_6312), .B(n_8_0_2640), .C1(n_8_0_2641), 
      .C2(n_8_0_6307), .ZN(n_8_0_2639));
   NAND2_X1 i_8_0_2512 (.A1(n_8_0_6991), .A2(n_8_0_6307), .ZN(n_8_0_2640));
   OAI21_X1 i_8_0_2513 (.A(n_8_0_2642), .B1(n_8_0_6323), .B2(n_8_0_6992), 
      .ZN(n_8_0_2641));
   OAI211_X1 i_8_0_2514 (.A(n_8_0_2643), .B(n_8_0_6323), .C1(in_data[20]), 
      .C2(n_8_0_6318), .ZN(n_8_0_2642));
   OAI211_X1 i_8_0_2515 (.A(n_8_0_6318), .B(n_8_0_2644), .C1(n_8_0_6994), 
      .C2(n_8_0_6320), .ZN(n_8_0_2643));
   NAND2_X1 i_8_0_2516 (.A1(in_data[28]), .A2(n_8_0_6320), .ZN(n_8_0_2644));
   INV_X1 i_8_0_2517 (.A(n_8_0_2645), .ZN(n_104));
   OAI21_X1 i_8_0_2518 (.A(n_8_0_2646), .B1(n_8_0_2649), .B2(n_8_0_6358), 
      .ZN(n_8_0_2645));
   OAI21_X1 i_8_0_2519 (.A(n_8_0_2647), .B1(n_8_0_6359), .B2(n_8_0_6988), 
      .ZN(n_8_0_2646));
   OAI221_X1 i_8_0_2520 (.A(n_8_0_6359), .B1(n_8_0_6364), .B2(in_data[4]), 
      .C1(n_8_0_6370), .C2(n_8_0_2648), .ZN(n_8_0_2647));
   NAND2_X1 i_8_0_2521 (.A1(n_8_0_6990), .A2(n_8_0_6364), .ZN(n_8_0_2648));
   OAI21_X1 i_8_0_2522 (.A(n_8_0_2650), .B1(n_8_0_2651), .B2(n_8_0_6346), 
      .ZN(n_8_0_2649));
   NAND2_X1 i_8_0_2523 (.A1(n_8_0_6346), .A2(in_data[12]), .ZN(n_8_0_2650));
   OAI21_X1 i_8_0_2524 (.A(n_8_0_2652), .B1(n_8_0_6353), .B2(in_data[16]), 
      .ZN(n_8_0_2651));
   OAI211_X1 i_8_0_2525 (.A(n_8_0_6353), .B(n_8_0_2653), .C1(n_8_0_2654), 
      .C2(n_8_0_6331), .ZN(n_8_0_2652));
   NAND2_X1 i_8_0_2526 (.A1(in_data[20]), .A2(n_8_0_6331), .ZN(n_8_0_2653));
   INV_X1 i_8_0_2527 (.A(n_8_0_2655), .ZN(n_8_0_2654));
   MUX2_X1 i_8_0_2528 (.A(in_data[28]), .B(in_data[24]), .S(n_8_0_6337), 
      .Z(n_8_0_2655));
   OAI21_X1 i_8_0_2529 (.A(n_8_0_2656), .B1(n_8_0_6401), .B2(n_8_0_6988), 
      .ZN(n_105));
   OAI211_X1 i_8_0_2530 (.A(n_8_0_6401), .B(n_8_0_2657), .C1(n_8_0_2658), 
      .C2(n_8_0_6383), .ZN(n_8_0_2656));
   NAND2_X1 i_8_0_2531 (.A1(n_8_0_6383), .A2(n_8_0_6989), .ZN(n_8_0_2657));
   AOI21_X1 i_8_0_2532 (.A(n_8_0_2659), .B1(n_8_0_2660), .B2(n_8_0_6406), 
      .ZN(n_8_0_2658));
   NOR2_X1 i_8_0_2533 (.A1(in_data[8]), .A2(n_8_0_6406), .ZN(n_8_0_2659));
   MUX2_X1 i_8_0_2534 (.A(n_8_0_2661), .B(n_8_0_6991), .S(n_8_0_6378), .Z(
      n_8_0_2660));
   OAI21_X1 i_8_0_2535 (.A(n_8_0_2662), .B1(n_8_0_2663), .B2(n_8_0_6410), 
      .ZN(n_8_0_2661));
   NAND2_X1 i_8_0_2536 (.A1(n_8_0_6992), .A2(n_8_0_6410), .ZN(n_8_0_2662));
   AOI21_X1 i_8_0_2537 (.A(n_8_0_2664), .B1(n_8_0_2665), .B2(n_8_0_6396), 
      .ZN(n_8_0_2663));
   NOR2_X1 i_8_0_2538 (.A1(n_8_0_6396), .A2(in_data[20]), .ZN(n_8_0_2664));
   OAI21_X1 i_8_0_2539 (.A(n_8_0_2666), .B1(n_8_0_6389), .B2(in_data[24]), 
      .ZN(n_8_0_2665));
   NAND2_X1 i_8_0_2540 (.A1(n_8_0_6389), .A2(n_8_0_6995), .ZN(n_8_0_2666));
   AOI21_X1 i_8_0_2541 (.A(n_8_0_2667), .B1(n_8_0_6462), .B2(n_8_0_6988), 
      .ZN(n_106));
   AOI21_X1 i_8_0_2542 (.A(n_8_0_2668), .B1(n_8_0_2669), .B2(n_8_0_6476), 
      .ZN(n_8_0_2667));
   OAI21_X1 i_8_0_2543 (.A(n_8_0_6463), .B1(n_8_0_6476), .B2(n_8_0_6989), 
      .ZN(n_8_0_2668));
   OAI22_X1 i_8_0_2544 (.A1(n_8_0_2670), .A2(n_8_0_2672), .B1(n_8_0_6454), 
      .B2(n_8_0_6990), .ZN(n_8_0_2669));
   OAI21_X1 i_8_0_2545 (.A(n_8_0_6454), .B1(n_8_0_2673), .B2(n_8_0_2671), 
      .ZN(n_8_0_2670));
   OAI21_X1 i_8_0_2546 (.A(n_8_0_6430), .B1(n_8_0_6425), .B2(n_8_0_6992), 
      .ZN(n_8_0_2671));
   NOR2_X1 i_8_0_2547 (.A1(n_8_0_6430), .A2(in_data[12]), .ZN(n_8_0_2672));
   AOI21_X1 i_8_0_2548 (.A(n_8_0_2674), .B1(n_8_0_2675), .B2(n_8_0_6449), 
      .ZN(n_8_0_2673));
   OAI21_X1 i_8_0_2549 (.A(n_8_0_6425), .B1(n_8_0_6449), .B2(in_data[20]), 
      .ZN(n_8_0_2674));
   OAI21_X1 i_8_0_2550 (.A(n_8_0_2676), .B1(n_8_0_6443), .B2(in_data[28]), 
      .ZN(n_8_0_2675));
   NAND2_X1 i_8_0_2551 (.A1(n_8_0_6443), .A2(n_8_0_6994), .ZN(n_8_0_2676));
   AOI21_X1 i_8_0_2552 (.A(n_8_0_2687), .B1(n_8_0_2677), .B2(n_8_0_6488), 
      .ZN(n_107));
   AOI21_X1 i_8_0_2553 (.A(n_8_0_2678), .B1(n_8_0_2679), .B2(n_8_0_6490), 
      .ZN(n_8_0_2677));
   MUX2_X1 i_8_0_2554 (.A(n_8_0_2681), .B(in_data[4]), .S(n_8_0_6501), .Z(
      n_8_0_2678));
   OAI21_X1 i_8_0_2555 (.A(n_8_0_2680), .B1(n_8_0_6483), .B2(n_8_0_6994), 
      .ZN(n_8_0_2679));
   NAND2_X1 i_8_0_2556 (.A1(n_8_0_6483), .A2(in_data[28]), .ZN(n_8_0_2680));
   OAI22_X1 i_8_0_2557 (.A1(n_8_0_2682), .A2(n_8_0_2683), .B1(n_8_0_6492), 
      .B2(n_8_0_6990), .ZN(n_8_0_2681));
   OAI21_X1 i_8_0_2558 (.A(n_8_0_6492), .B1(n_8_0_6497), .B2(in_data[12]), 
      .ZN(n_8_0_2682));
   AND2_X1 i_8_0_2559 (.A1(n_8_0_2684), .A2(n_8_0_6497), .ZN(n_8_0_2683));
   OAI21_X1 i_8_0_2560 (.A(n_8_0_2685), .B1(n_8_0_6495), .B2(in_data[16]), 
      .ZN(n_8_0_2684));
   NAND2_X1 i_8_0_2561 (.A1(n_8_0_2686), .A2(n_8_0_6495), .ZN(n_8_0_2685));
   NAND3_X1 i_8_0_2562 (.A1(n_8_0_6500), .A2(n_8_0_6499), .A3(in_data[20]), 
      .ZN(n_8_0_2686));
   NOR2_X1 i_8_0_2563 (.A1(in_data[0]), .A2(n_8_0_6488), .ZN(n_8_0_2687));
   OAI22_X1 i_8_0_2564 (.A1(n_8_0_2689), .A2(n_8_0_2688), .B1(n_8_0_6988), 
      .B2(n_8_0_6538), .ZN(n_108));
   OAI21_X1 i_8_0_2565 (.A(n_8_0_6538), .B1(n_8_0_6546), .B2(in_data[4]), 
      .ZN(n_8_0_2688));
   NOR2_X1 i_8_0_2566 (.A1(n_8_0_6545), .A2(n_8_0_2690), .ZN(n_8_0_2689));
   AOI21_X1 i_8_0_2567 (.A(n_8_0_2691), .B1(n_8_0_6506), .B2(n_8_0_6990), 
      .ZN(n_8_0_2690));
   NOR2_X1 i_8_0_2568 (.A1(n_8_0_6506), .A2(n_8_0_2692), .ZN(n_8_0_2691));
   AOI21_X1 i_8_0_2569 (.A(n_8_0_2693), .B1(n_8_0_6552), .B2(n_8_0_6991), 
      .ZN(n_8_0_2692));
   NOR2_X1 i_8_0_2570 (.A1(n_8_0_6552), .A2(n_8_0_2694), .ZN(n_8_0_2693));
   AOI21_X1 i_8_0_2571 (.A(n_8_0_2695), .B1(n_8_0_6561), .B2(n_8_0_6992), 
      .ZN(n_8_0_2694));
   NOR2_X1 i_8_0_2572 (.A1(n_8_0_6561), .A2(n_8_0_2696), .ZN(n_8_0_2695));
   AOI21_X1 i_8_0_2573 (.A(n_8_0_2697), .B1(n_8_0_2698), .B2(n_8_0_6533), 
      .ZN(n_8_0_2696));
   NOR2_X1 i_8_0_2574 (.A1(n_8_0_6533), .A2(in_data[20]), .ZN(n_8_0_2697));
   OAI21_X1 i_8_0_2575 (.A(n_8_0_2699), .B1(n_8_0_6524), .B2(in_data[28]), 
      .ZN(n_8_0_2698));
   NAND2_X1 i_8_0_2576 (.A1(n_8_0_6524), .A2(n_8_0_6994), .ZN(n_8_0_2699));
   AOI22_X1 i_8_0_2577 (.A1(n_8_0_2700), .A2(n_8_0_2701), .B1(n_8_0_6614), 
      .B2(n_8_0_6988), .ZN(n_109));
   AOI21_X1 i_8_0_2578 (.A(n_8_0_6614), .B1(n_8_0_6582), .B2(in_data[4]), 
      .ZN(n_8_0_2700));
   OAI211_X1 i_8_0_2579 (.A(n_8_0_6581), .B(n_8_0_2702), .C1(in_data[8]), 
      .C2(n_8_0_6617), .ZN(n_8_0_2701));
   OAI211_X1 i_8_0_2580 (.A(n_8_0_6617), .B(n_8_0_2703), .C1(n_8_0_2704), 
      .C2(n_8_0_6620), .ZN(n_8_0_2702));
   NAND2_X1 i_8_0_2581 (.A1(n_8_0_6620), .A2(in_data[12]), .ZN(n_8_0_2703));
   INV_X1 i_8_0_2582 (.A(n_8_0_2705), .ZN(n_8_0_2704));
   OAI21_X1 i_8_0_2583 (.A(n_8_0_2706), .B1(n_8_0_6570), .B2(n_8_0_6992), 
      .ZN(n_8_0_2705));
   OAI211_X1 i_8_0_2584 (.A(n_8_0_6570), .B(n_8_0_2707), .C1(n_8_0_2708), 
      .C2(n_8_0_6602), .ZN(n_8_0_2706));
   NAND2_X1 i_8_0_2585 (.A1(n_8_0_6602), .A2(n_8_0_6993), .ZN(n_8_0_2707));
   AOI21_X1 i_8_0_2586 (.A(n_8_0_2709), .B1(n_8_0_6600), .B2(n_8_0_6995), 
      .ZN(n_8_0_2708));
   NOR2_X1 i_8_0_2587 (.A1(n_8_0_6600), .A2(in_data[24]), .ZN(n_8_0_2709));
   AOI21_X1 i_8_0_2588 (.A(n_8_0_2710), .B1(n_8_0_6713), .B2(n_8_0_6988), 
      .ZN(n_110));
   AOI21_X1 i_8_0_2589 (.A(n_8_0_2711), .B1(n_8_0_2712), .B2(n_8_0_6739), 
      .ZN(n_8_0_2710));
   OAI221_X1 i_8_0_2590 (.A(n_8_0_6730), .B1(n_8_0_6722), .B2(n_8_0_6714), 
      .C1(n_8_0_6739), .C2(n_8_0_6989), .ZN(n_8_0_2711));
   MUX2_X1 i_8_0_2591 (.A(n_8_0_2713), .B(in_data[8]), .S(n_8_0_2714), .Z(
      n_8_0_2712));
   MUX2_X1 i_8_0_2592 (.A(n_8_0_2715), .B(in_data[12]), .S(n_8_0_2716), .Z(
      n_8_0_2713));
   NAND2_X1 i_8_0_2593 (.A1(n_8_0_6824), .A2(n_8_0_6672), .ZN(n_8_0_2714));
   MUX2_X1 i_8_0_2594 (.A(in_data[16]), .B(n_8_0_2717), .S(n_8_0_2718), .Z(
      n_8_0_2715));
   NAND2_X1 i_8_0_2595 (.A1(n_8_0_6795), .A2(n_8_0_6627), .ZN(n_8_0_2716));
   MUX2_X1 i_8_0_2596 (.A(n_8_0_2719), .B(in_data[20]), .S(n_8_0_2720), .Z(
      n_8_0_2717));
   AOI21_X1 i_8_0_2597 (.A(n_8_0_6838), .B1(n_8_0_6650), .B2(n_8_0_6646), 
      .ZN(n_8_0_2718));
   MUX2_X1 i_8_0_2598 (.A(in_data[24]), .B(in_data[28]), .S(n_8_0_2721), 
      .Z(n_8_0_2719));
   NAND2_X1 i_8_0_2599 (.A1(n_8_0_6772), .A2(n_8_0_6701), .ZN(n_8_0_2720));
   NOR2_X1 i_8_0_2600 (.A1(n_8_0_6781), .A2(n_8_0_6687), .ZN(n_8_0_2721));
   AOI21_X1 i_8_0_2601 (.A(n_8_0_6853), .B1(n_8_0_6770), .B2(n_8_0_2722), 
      .ZN(n_111));
   NOR4_X1 i_8_0_2602 (.A1(n_8_0_2733), .A2(n_8_0_2728), .A3(n_8_0_2726), 
      .A4(n_8_0_2723), .ZN(n_8_0_2722));
   OAI21_X1 i_8_0_2603 (.A(n_8_0_2724), .B1(n_8_0_2768), .B2(\out_as[5] [0]), 
      .ZN(n_8_0_2723));
   NAND2_X1 i_8_0_2604 (.A1(n_8_0_2828), .A2(n_8_0_2725), .ZN(n_8_0_2724));
   NAND2_X1 i_8_0_2605 (.A1(n_8_0_2829), .A2(n_8_0_2725), .ZN(n_8_0_1167));
   INV_X1 i_8_0_2606 (.A(n_8_0_2725), .ZN(n_8_0_1168));
   NOR2_X1 i_8_0_2607 (.A1(\out_as[2] [1]), .A2(\out_as[2] [0]), .ZN(n_8_0_2725));
   NOR2_X1 i_8_0_2608 (.A1(n_8_0_3194), .A2(n_8_0_1169), .ZN(n_8_0_2726));
   NAND3_X1 i_8_0_2609 (.A1(n_8_0_2842), .A2(n_8_0_7073), .A3(n_8_0_7074), 
      .ZN(n_8_0_1169));
   INV_X1 i_8_0_2610 (.A(n_8_0_2727), .ZN(n_8_0_1170));
   NOR2_X1 i_8_0_2611 (.A1(n_8_0_1171), .A2(\out_as[1] [2]), .ZN(n_8_0_2727));
   NAND2_X1 i_8_0_2612 (.A1(n_8_0_7074), .A2(n_8_0_7073), .ZN(n_8_0_1171));
   OAI221_X1 i_8_0_2613 (.A(n_8_0_2729), .B1(n_8_0_1178), .B2(n_8_0_2961), 
      .C1(n_8_0_3206), .C2(n_8_0_1175), .ZN(n_8_0_2728));
   NAND2_X1 i_8_0_2614 (.A1(n_8_0_2987), .A2(n_8_0_2730), .ZN(n_8_0_2729));
   NAND2_X1 i_8_0_2615 (.A1(n_8_0_2730), .A2(n_8_0_7038), .ZN(n_8_0_1172));
   INV_X1 i_8_0_2616 (.A(n_8_0_2730), .ZN(n_8_0_1173));
   NOR2_X1 i_8_0_2617 (.A1(n_8_0_1188), .A2(\out_as[4] [0]), .ZN(n_8_0_2730));
   OR2_X1 i_8_0_2618 (.A1(\out_as[4] [1]), .A2(\out_as[4] [0]), .ZN(n_8_0_1174));
   NAND2_X1 i_8_0_2619 (.A1(n_8_0_2836), .A2(n_8_0_2731), .ZN(n_8_0_1175));
   INV_X1 i_8_0_2620 (.A(n_8_0_2731), .ZN(n_8_0_1176));
   NOR2_X1 i_8_0_2621 (.A1(\out_as[0] [1]), .A2(\out_as[0] [0]), .ZN(n_8_0_2731));
   NAND2_X1 i_8_0_2622 (.A1(n_8_0_2732), .A2(n_8_0_7050), .ZN(n_8_0_1177));
   INV_X1 i_8_0_2623 (.A(n_8_0_2732), .ZN(n_8_0_1178));
   NOR2_X1 i_8_0_2624 (.A1(n_8_0_1187), .A2(\out_as[3] [0]), .ZN(n_8_0_2732));
   OR2_X1 i_8_0_2625 (.A1(\out_as[3] [1]), .A2(\out_as[3] [0]), .ZN(n_8_0_1179));
   OAI211_X1 i_8_0_2626 (.A(n_8_0_6755), .B(n_8_0_2735), .C1(n_8_0_1180), 
      .C2(n_8_0_3203), .ZN(n_8_0_2733));
   NAND2_X1 i_8_0_2627 (.A1(n_8_0_2823), .A2(n_8_0_2734), .ZN(n_8_0_1180));
   INV_X1 i_8_0_2628 (.A(n_8_0_2734), .ZN(n_8_0_1181));
   NOR2_X1 i_8_0_2629 (.A1(\out_as[6] [1]), .A2(\out_as[6] [0]), .ZN(n_8_0_2734));
   AOI21_X1 i_8_0_2630 (.A(n_8_0_6729), .B1(n_8_0_2982), .B2(n_8_0_2736), 
      .ZN(n_8_0_2735));
   INV_X1 i_8_0_2631 (.A(n_8_0_2736), .ZN(n_8_0_1182));
   NOR2_X1 i_8_0_2632 (.A1(n_8_0_1193), .A2(\out_as[7] [0]), .ZN(n_8_0_2736));
   OR2_X1 i_8_0_2633 (.A1(\out_as[7] [1]), .A2(\out_as[7] [0]), .ZN(n_8_0_1183));
   OAI21_X1 i_8_0_2636 (.A(n_8_0_2739), .B1(n_8_0_4560), .B2(n_8_0_5522), 
      .ZN(n_8_0_2738));
   OAI21_X1 i_8_0_2637 (.A(n_8_0_2740), .B1(n_8_0_2822), .B2(\out_as[6] [1]), 
      .ZN(n_8_0_2739));
   OAI21_X1 i_8_0_2638 (.A(n_8_0_6754), .B1(n_8_0_5522), .B2(n_8_0_4562), 
      .ZN(n_8_0_2740));
   NAND2_X1 i_8_0_2639 (.A1(n_8_0_2823), .A2(n_8_0_7013), .ZN(n_8_0_1184));
   NAND2_X1 i_8_0_2640 (.A1(n_8_0_7014), .A2(n_8_0_7013), .ZN(n_8_0_1185));
   AOI21_X1 i_8_0_2641 (.A(n_8_0_2742), .B1(n_8_0_6838), .B2(n_8_0_2743), 
      .ZN(n_8_0_2741));
   AOI211_X1 i_8_0_2642 (.A(n_8_0_2961), .B(n_8_0_1187), .C1(n_8_0_5501), 
      .C2(n_8_0_3686), .ZN(n_8_0_2742));
   OAI211_X1 i_8_0_2643 (.A(n_8_0_5501), .B(n_8_0_3686), .C1(n_8_0_2961), 
      .C2(n_8_0_1187), .ZN(n_8_0_2743));
   NAND2_X1 i_8_0_2644 (.A1(n_8_0_2744), .A2(n_8_0_7050), .ZN(n_8_0_1186));
   INV_X1 i_8_0_2645 (.A(n_8_0_2744), .ZN(n_8_0_1187));
   NOR2_X1 i_8_0_2646 (.A1(\out_as[3] [2]), .A2(\out_as[3] [1]), .ZN(n_8_0_2744));
   OAI21_X1 i_8_0_2647 (.A(n_8_0_2746), .B1(n_8_0_3221), .B2(n_8_0_6031), 
      .ZN(n_8_0_2745));
   OAI21_X1 i_8_0_2648 (.A(n_8_0_2748), .B1(n_8_0_1188), .B2(n_8_0_2986), 
      .ZN(n_8_0_2746));
   INV_X1 i_8_0_2649 (.A(n_8_0_2747), .ZN(n_8_0_1188));
   NOR2_X1 i_8_0_2650 (.A1(\out_as[4] [2]), .A2(\out_as[4] [1]), .ZN(n_8_0_2747));
   OAI21_X1 i_8_0_2651 (.A(n_8_0_6794), .B1(n_8_0_6031), .B2(n_8_0_3222), 
      .ZN(n_8_0_2748));
   OAI21_X1 i_8_0_2652 (.A(n_8_0_2750), .B1(n_8_0_3003), .B2(n_8_0_6344), 
      .ZN(n_8_0_2749));
   OAI221_X1 i_8_0_2653 (.A(n_8_0_4132), .B1(n_8_0_2834), .B2(\out_as[0] [1]), 
      .C1(n_8_0_6811), .C2(n_8_0_5506), .ZN(n_8_0_2750));
   NAND2_X1 i_8_0_2654 (.A1(n_8_0_2978), .A2(n_8_0_2751), .ZN(n_8_0_1189));
   NAND2_X1 i_8_0_2655 (.A1(n_8_0_2751), .A2(n_8_0_7087), .ZN(n_8_0_1190));
   INV_X1 i_8_0_2656 (.A(n_8_0_2751), .ZN(n_8_0_1191));
   NOR2_X1 i_8_0_2657 (.A1(\out_as[0] [2]), .A2(\out_as[0] [1]), .ZN(n_8_0_2751));
   NAND2_X1 i_8_0_2663 (.A1(n_8_0_2757), .A2(n_8_0_7003), .ZN(n_8_0_1192));
   INV_X1 i_8_0_2664 (.A(n_8_0_2757), .ZN(n_8_0_1193));
   NOR2_X1 i_8_0_2665 (.A1(\out_as[7] [2]), .A2(\out_as[7] [1]), .ZN(n_8_0_2757));
   AOI21_X1 i_8_0_2667 (.A(n_8_0_2760), .B1(n_8_0_2828), .B2(n_8_0_7061), 
      .ZN(n_8_0_2759));
   NAND2_X1 i_8_0_2668 (.A1(n_8_0_2829), .A2(n_8_0_7061), .ZN(n_8_0_1194));
   NAND2_X1 i_8_0_2669 (.A1(n_8_0_7062), .A2(n_8_0_7061), .ZN(n_8_0_1195));
   AOI21_X1 i_8_0_2670 (.A(n_8_0_6772), .B1(n_8_0_5515), .B2(n_8_0_4367), 
      .ZN(n_8_0_2760));
   INV_X1 i_8_0_2672 (.A(n_8_0_2763), .ZN(n_8_0_2762));
   AOI211_X1 i_8_0_2673 (.A(\out_as[1] [1]), .B(n_8_0_2840), .C1(n_8_0_4199), 
      .C2(n_8_0_5526), .ZN(n_8_0_2763));
   NAND2_X1 i_8_0_2674 (.A1(n_8_0_2842), .A2(n_8_0_7074), .ZN(n_8_0_1196));
   INV_X1 i_8_0_2675 (.A(n_8_0_2764), .ZN(n_8_0_1197));
   NOR2_X1 i_8_0_2676 (.A1(\out_as[1] [2]), .A2(\out_as[1] [1]), .ZN(n_8_0_2764));
   AOI21_X1 i_8_0_2678 (.A(n_8_0_4109), .B1(n_8_0_6830), .B2(n_8_0_2767), 
      .ZN(n_8_0_2766));
   NAND2_X1 i_8_0_2679 (.A1(n_8_0_2816), .A2(n_8_0_2769), .ZN(n_8_0_1198));
   INV_X1 i_8_0_2680 (.A(n_8_0_2768), .ZN(n_8_0_2767));
   NAND2_X1 i_8_0_2681 (.A1(n_8_0_2957), .A2(n_8_0_2769), .ZN(n_8_0_2768));
   NAND2_X1 i_8_0_2682 (.A1(n_8_0_2958), .A2(n_8_0_2769), .ZN(n_8_0_1199));
   NAND2_X1 i_8_0_2683 (.A1(n_8_0_2817), .A2(n_8_0_7025), .ZN(n_8_0_1200));
   INV_X1 i_8_0_2684 (.A(n_8_0_2769), .ZN(n_8_0_1201));
   NOR2_X1 i_8_0_2685 (.A1(\out_as[5] [2]), .A2(\out_as[5] [1]), .ZN(n_8_0_2769));
   AOI21_X1 i_8_0_2686 (.A(n_8_0_6853), .B1(n_8_0_2788), .B2(n_8_0_2770), 
      .ZN(n_112));
   NOR4_X1 i_8_0_2687 (.A1(n_8_0_2771), .A2(n_8_0_2774), .A3(n_8_0_2792), 
      .A4(n_8_0_2793), .ZN(n_8_0_2770));
   OR4_X1 i_8_0_2688 (.A1(n_8_0_2784), .A2(n_8_0_2772), .A3(n_8_0_2781), 
      .A4(n_8_0_2798), .ZN(n_8_0_2771));
   NAND3_X1 i_8_0_2689 (.A1(n_8_0_2801), .A2(n_8_0_2777), .A3(n_8_0_2773), 
      .ZN(n_8_0_2772));
   OAI21_X1 i_8_0_2690 (.A(n_8_0_6810), .B1(n_8_0_5554), .B2(n_8_0_4603), 
      .ZN(n_8_0_2773));
   NOR3_X1 i_8_0_2691 (.A1(n_8_0_2776), .A2(n_8_0_1202), .A3(n_8_0_3643), 
      .ZN(n_8_0_2774));
   NAND2_X1 i_8_0_2692 (.A1(n_8_0_2978), .A2(n_8_0_2775), .ZN(n_8_0_1202));
   INV_X1 i_8_0_2693 (.A(n_8_0_2775), .ZN(n_8_0_1203));
   NOR2_X1 i_8_0_2694 (.A1(\out_as[0] [2]), .A2(n_8_0_539), .ZN(n_8_0_2775));
   NOR2_X1 i_8_0_2695 (.A1(n_8_0_6420), .A2(n_8_0_3003), .ZN(n_8_0_2776));
   OAI22_X1 i_8_0_2696 (.A1(n_8_0_2780), .A2(n_8_0_2778), .B1(n_8_0_6092), 
      .B2(n_8_0_3221), .ZN(n_8_0_2777));
   NOR2_X1 i_8_0_2697 (.A1(n_8_0_2986), .A2(n_8_0_1204), .ZN(n_8_0_2778));
   INV_X1 i_8_0_2698 (.A(n_8_0_2779), .ZN(n_8_0_1204));
   NOR2_X1 i_8_0_2699 (.A1(\out_as[4] [2]), .A2(n_8_0_519), .ZN(n_8_0_2779));
   AOI21_X1 i_8_0_2700 (.A(n_8_0_6795), .B1(n_8_0_6093), .B2(n_8_0_3223), 
      .ZN(n_8_0_2780));
   AOI22_X1 i_8_0_2701 (.A1(n_8_0_5543), .A2(n_8_0_4561), .B1(n_8_0_4347), 
      .B2(n_8_0_2782), .ZN(n_8_0_2781));
   AOI21_X1 i_8_0_2702 (.A(n_8_0_2783), .B1(n_8_0_5544), .B2(n_8_0_6754), 
      .ZN(n_8_0_2782));
   NOR2_X1 i_8_0_2703 (.A1(n_8_0_2822), .A2(n_8_0_509), .ZN(n_8_0_2783));
   OR2_X1 i_8_0_2704 (.A1(n_8_0_1221), .A2(n_8_0_509), .ZN(n_8_0_1205));
   OR2_X1 i_8_0_2705 (.A1(\out_as[6] [2]), .A2(n_8_0_509), .ZN(n_8_0_1206));
   OAI21_X1 i_8_0_2706 (.A(n_8_0_2785), .B1(n_8_0_5548), .B2(n_8_0_6782), 
      .ZN(n_8_0_2784));
   OAI21_X1 i_8_0_2707 (.A(n_8_0_2786), .B1(n_8_0_4198), .B2(n_8_0_5547), 
      .ZN(n_8_0_2785));
   OAI21_X1 i_8_0_2708 (.A(n_8_0_4231), .B1(n_8_0_3194), .B2(n_8_0_1207), 
      .ZN(n_8_0_2786));
   OR2_X1 i_8_0_2709 (.A1(n_8_0_1208), .A2(\out_as[1] [3]), .ZN(n_8_0_1207));
   INV_X1 i_8_0_2710 (.A(n_8_0_2787), .ZN(n_8_0_1208));
   NOR2_X1 i_8_0_2711 (.A1(\out_as[1] [2]), .A2(n_8_0_534), .ZN(n_8_0_2787));
   INV_X1 i_8_0_2712 (.A(n_8_0_2789), .ZN(n_8_0_2788));
   OAI211_X1 i_8_0_2713 (.A(n_8_0_2790), .B(n_8_0_3227), .C1(n_8_0_6098), 
      .C2(n_8_0_6824), .ZN(n_8_0_2789));
   OAI211_X1 i_8_0_2714 (.A(n_8_0_2957), .B(n_8_0_2791), .C1(n_8_0_6097), 
      .C2(n_8_0_3226), .ZN(n_8_0_2790));
   NAND2_X1 i_8_0_2715 (.A1(n_8_0_2791), .A2(n_8_0_7027), .ZN(n_8_0_1209));
   INV_X1 i_8_0_2716 (.A(n_8_0_2791), .ZN(n_8_0_1210));
   NOR2_X1 i_8_0_2717 (.A1(\out_as[5] [2]), .A2(n_8_0_514), .ZN(n_8_0_2791));
   NOR2_X1 i_8_0_2718 (.A1(n_8_0_2795), .A2(n_8_0_2797), .ZN(n_8_0_2792));
   AOI21_X1 i_8_0_2719 (.A(n_8_0_6232), .B1(n_8_0_2797), .B2(n_8_0_2795), 
      .ZN(n_8_0_2793));
   NAND2_X1 i_8_0_2720 (.A1(n_8_0_2795), .A2(n_8_0_2797), .ZN(n_8_0_2794));
   NAND2_X1 i_8_0_2721 (.A1(n_8_0_2982), .A2(n_8_0_2796), .ZN(n_8_0_2795));
   NAND2_X1 i_8_0_2722 (.A1(n_8_0_2796), .A2(n_8_0_7003), .ZN(n_8_0_1211));
   INV_X1 i_8_0_2723 (.A(n_8_0_2796), .ZN(n_8_0_1212));
   NOR2_X1 i_8_0_2724 (.A1(\out_as[7] [2]), .A2(n_8_0_504), .ZN(n_8_0_2796));
   NOR2_X1 i_8_0_2725 (.A1(n_8_0_5560), .A2(n_8_0_4423), .ZN(n_8_0_2797));
   AOI21_X1 i_8_0_2726 (.A(n_8_0_2799), .B1(n_8_0_4127), .B2(n_8_0_5552), 
      .ZN(n_8_0_2798));
   AOI21_X1 i_8_0_2727 (.A(n_8_0_2800), .B1(n_8_0_2828), .B2(n_8_0_6861), 
      .ZN(n_8_0_2799));
   AOI21_X1 i_8_0_2728 (.A(n_8_0_6772), .B1(n_8_0_6400), .B2(n_8_0_3020), 
      .ZN(n_8_0_2800));
   OAI21_X1 i_8_0_2729 (.A(n_8_0_2804), .B1(n_8_0_2802), .B2(n_8_0_3684), 
      .ZN(n_8_0_2801));
   OAI22_X1 i_8_0_2730 (.A1(n_8_0_6837), .A2(n_8_0_5564), .B1(n_8_0_2961), 
      .B2(n_8_0_1213), .ZN(n_8_0_2802));
   INV_X1 i_8_0_2731 (.A(n_8_0_2803), .ZN(n_8_0_1213));
   NOR2_X1 i_8_0_2732 (.A1(\out_as[3] [2]), .A2(n_8_0_524), .ZN(n_8_0_2803));
   NAND2_X1 i_8_0_2733 (.A1(n_8_0_6414), .A2(n_8_0_3000), .ZN(n_8_0_2804));
   AOI21_X1 i_8_0_2734 (.A(n_8_0_6853), .B1(n_8_0_2805), .B2(n_8_0_2830), 
      .ZN(n_113));
   AND4_X1 i_8_0_2735 (.A1(n_8_0_2819), .A2(n_8_0_2806), .A3(n_8_0_2807), 
      .A4(n_8_0_2843), .ZN(n_8_0_2805));
   NOR4_X1 i_8_0_2736 (.A1(n_8_0_2837), .A2(n_8_0_2812), .A3(n_8_0_2809), 
      .A4(n_8_0_2824), .ZN(n_8_0_2806));
   OAI21_X1 i_8_0_2737 (.A(n_8_0_2818), .B1(n_8_0_2808), .B2(n_8_0_5595), 
      .ZN(n_8_0_2807));
   AOI21_X1 i_8_0_2738 (.A(n_8_0_3697), .B1(n_8_0_2834), .B2(n_8_0_4132), 
      .ZN(n_8_0_2808));
   OAI221_X1 i_8_0_2739 (.A(n_8_0_3683), .B1(n_8_0_2810), .B2(\out_as[3] [2]), 
      .C1(n_8_0_6837), .C2(n_8_0_5581), .ZN(n_8_0_2809));
   INV_X1 i_8_0_2740 (.A(n_8_0_2811), .ZN(n_8_0_2810));
   AOI21_X1 i_8_0_2741 (.A(n_8_0_2961), .B1(n_8_0_3452), .B2(n_8_0_5581), 
      .ZN(n_8_0_2811));
   NAND2_X1 i_8_0_2742 (.A1(n_8_0_7050), .A2(n_8_0_7049), .ZN(n_8_0_1214));
   AOI21_X1 i_8_0_2743 (.A(n_8_0_2813), .B1(n_8_0_2814), .B2(n_8_0_2815), 
      .ZN(n_8_0_2812));
   NOR2_X1 i_8_0_2744 (.A1(n_8_0_6136), .A2(n_8_0_3226), .ZN(n_8_0_2813));
   OAI21_X1 i_8_0_2745 (.A(n_8_0_6825), .B1(n_8_0_6136), .B2(n_8_0_3270), 
      .ZN(n_8_0_2814));
   NAND2_X1 i_8_0_2746 (.A1(n_8_0_3186), .A2(n_8_0_2817), .ZN(n_8_0_2815));
   NAND2_X1 i_8_0_2747 (.A1(n_8_0_2816), .A2(n_8_0_7026), .ZN(n_8_0_1215));
   INV_X1 i_8_0_2748 (.A(n_8_0_2816), .ZN(n_8_0_1216));
   NOR2_X1 i_8_0_2749 (.A1(n_8_0_1354), .A2(\out_as[5] [3]), .ZN(n_8_0_2816));
   NAND2_X1 i_8_0_2750 (.A1(n_8_0_2958), .A2(n_8_0_7026), .ZN(n_8_0_1217));
   INV_X1 i_8_0_2751 (.A(n_8_0_2817), .ZN(n_8_0_1218));
   NOR2_X1 i_8_0_2752 (.A1(\out_as[5] [3]), .A2(\out_as[5] [2]), .ZN(n_8_0_2817));
   NAND2_X1 i_8_0_2753 (.A1(n_8_0_6811), .A2(n_8_0_2834), .ZN(n_8_0_2818));
   OAI22_X1 i_8_0_2754 (.A1(n_8_0_6754), .A2(n_8_0_2821), .B1(n_8_0_2820), 
      .B2(n_8_0_6746), .ZN(n_8_0_2819));
   OAI211_X1 i_8_0_2755 (.A(n_8_0_5626), .B(n_8_0_4563), .C1(n_8_0_6763), 
      .C2(n_8_0_2822), .ZN(n_8_0_2820));
   INV_X1 i_8_0_2756 (.A(n_8_0_2822), .ZN(n_8_0_2821));
   NAND3_X1 i_8_0_2757 (.A1(n_8_0_3647), .A2(n_8_0_2823), .A3(n_8_0_7016), 
      .ZN(n_8_0_2822));
   NAND2_X1 i_8_0_2758 (.A1(n_8_0_3204), .A2(n_8_0_2823), .ZN(n_8_0_1219));
   NAND2_X1 i_8_0_2759 (.A1(n_8_0_2823), .A2(n_8_0_7016), .ZN(n_8_0_1220));
   INV_X1 i_8_0_2760 (.A(n_8_0_2823), .ZN(n_8_0_1221));
   NOR2_X1 i_8_0_2761 (.A1(\out_as[6] [3]), .A2(\out_as[6] [2]), .ZN(n_8_0_2823));
   NAND2_X1 i_8_0_2762 (.A1(n_8_0_2827), .A2(n_8_0_2825), .ZN(n_8_0_2824));
   OAI21_X1 i_8_0_2763 (.A(n_8_0_2826), .B1(n_8_0_2828), .B2(n_8_0_6773), 
      .ZN(n_8_0_2825));
   NAND2_X1 i_8_0_2764 (.A1(n_8_0_6453), .A2(n_8_0_3020), .ZN(n_8_0_2826));
   NAND2_X1 i_8_0_2765 (.A1(n_8_0_6773), .A2(n_8_0_2828), .ZN(n_8_0_2827));
   NOR2_X1 i_8_0_2766 (.A1(n_8_0_3190), .A2(n_8_0_1224), .ZN(n_8_0_2828));
   NAND2_X1 i_8_0_2767 (.A1(n_8_0_3191), .A2(n_8_0_2829), .ZN(n_8_0_1222));
   NAND2_X1 i_8_0_2768 (.A1(n_8_0_2829), .A2(n_8_0_7064), .ZN(n_8_0_1223));
   INV_X1 i_8_0_2769 (.A(n_8_0_2829), .ZN(n_8_0_1224));
   NOR2_X1 i_8_0_2770 (.A1(\out_as[2] [3]), .A2(\out_as[2] [2]), .ZN(n_8_0_2829));
   AOI21_X1 i_8_0_2771 (.A(n_8_0_2831), .B1(n_8_0_2832), .B2(n_8_0_6729), 
      .ZN(n_8_0_2830));
   NOR3_X1 i_8_0_2772 (.A1(n_8_0_2833), .A2(n_8_0_1226), .A3(n_8_0_3211), 
      .ZN(n_8_0_2831));
   OAI21_X1 i_8_0_2773 (.A(n_8_0_2833), .B1(n_8_0_2981), .B2(\out_as[7] [2]), 
      .ZN(n_8_0_2832));
   NAND2_X1 i_8_0_2774 (.A1(n_8_0_2983), .A2(n_8_0_7002), .ZN(n_8_0_1225));
   NAND2_X1 i_8_0_2775 (.A1(n_8_0_7003), .A2(n_8_0_7002), .ZN(n_8_0_1226));
   NOR2_X1 i_8_0_2776 (.A1(n_8_0_6118), .A2(n_8_0_3243), .ZN(n_8_0_2833));
   NAND3_X1 i_8_0_2777 (.A1(n_8_0_2835), .A2(n_8_0_7088), .A3(n_8_0_7089), 
      .ZN(n_8_0_2834));
   INV_X1 i_8_0_2778 (.A(n_8_0_2835), .ZN(n_8_0_1227));
   NOR2_X1 i_8_0_2779 (.A1(n_8_0_1228), .A2(\out_as[0] [4]), .ZN(n_8_0_2835));
   INV_X1 i_8_0_2780 (.A(n_8_0_2836), .ZN(n_8_0_1228));
   NOR2_X1 i_8_0_2781 (.A1(\out_as[0] [3]), .A2(\out_as[0] [2]), .ZN(n_8_0_2836));
   AOI22_X1 i_8_0_2782 (.A1(n_8_0_6782), .A2(n_8_0_2840), .B1(n_8_0_2839), 
      .B2(n_8_0_2838), .ZN(n_8_0_2837));
   NAND3_X1 i_8_0_2783 (.A1(n_8_0_6785), .A2(n_8_0_3195), .A3(n_8_0_2842), 
      .ZN(n_8_0_2838));
   NOR2_X1 i_8_0_2784 (.A1(n_8_0_5586), .A2(n_8_0_4324), .ZN(n_8_0_2839));
   NAND2_X1 i_8_0_2785 (.A1(n_8_0_3195), .A2(n_8_0_2842), .ZN(n_8_0_2840));
   NAND2_X1 i_8_0_2786 (.A1(n_8_0_2841), .A2(n_8_0_7075), .ZN(n_8_0_1229));
   INV_X1 i_8_0_2787 (.A(n_8_0_2841), .ZN(n_8_0_1230));
   NOR2_X1 i_8_0_2788 (.A1(n_8_0_1356), .A2(\out_as[1] [3]), .ZN(n_8_0_2841));
   INV_X1 i_8_0_2789 (.A(n_8_0_2842), .ZN(n_8_0_1231));
   NOR2_X1 i_8_0_2790 (.A1(\out_as[1] [3]), .A2(\out_as[1] [2]), .ZN(n_8_0_2842));
   OAI21_X1 i_8_0_2791 (.A(n_8_0_2844), .B1(n_8_0_3221), .B2(n_8_0_6113), 
      .ZN(n_8_0_2843));
   OAI221_X1 i_8_0_2792 (.A(n_8_0_4058), .B1(n_8_0_2986), .B2(\out_as[4] [2]), 
      .C1(n_8_0_6795), .C2(n_8_0_5573), .ZN(n_8_0_2844));
   NAND2_X1 i_8_0_2793 (.A1(n_8_0_2988), .A2(n_8_0_7037), .ZN(n_8_0_1232));
   NAND2_X1 i_8_0_2794 (.A1(n_8_0_7038), .A2(n_8_0_7037), .ZN(n_8_0_1233));
   AOI21_X1 i_8_0_2795 (.A(n_8_0_6853), .B1(n_8_0_2846), .B2(n_8_0_2845), 
      .ZN(n_114));
   NOR4_X1 i_8_0_2796 (.A1(n_8_0_2863), .A2(n_8_0_2855), .A3(n_8_0_2852), 
      .A4(n_8_0_2875), .ZN(n_8_0_2845));
   AND3_X1 i_8_0_2797 (.A1(n_8_0_2871), .A2(n_8_0_2860), .A3(n_8_0_2847), 
      .ZN(n_8_0_2846));
   OAI22_X1 i_8_0_2798 (.A1(n_8_0_6794), .A2(n_8_0_2850), .B1(n_8_0_2848), 
      .B2(n_8_0_6170), .ZN(n_8_0_2847));
   INV_X1 i_8_0_2799 (.A(n_8_0_2849), .ZN(n_8_0_2848));
   AOI21_X1 i_8_0_2800 (.A(n_8_0_3222), .B1(n_8_0_6800), .B2(n_8_0_2850), 
      .ZN(n_8_0_2849));
   NOR2_X1 i_8_0_2801 (.A1(n_8_0_3199), .A2(n_8_0_1236), .ZN(n_8_0_2850));
   OR2_X1 i_8_0_2802 (.A1(n_8_0_1357), .A2(n_8_0_1236), .ZN(n_8_0_1234));
   NAND2_X1 i_8_0_2803 (.A1(n_8_0_2851), .A2(n_8_0_7039), .ZN(n_8_0_1235));
   INV_X1 i_8_0_2804 (.A(n_8_0_2851), .ZN(n_8_0_1236));
   NOR2_X1 i_8_0_2805 (.A1(\out_as[4] [3]), .A2(n_8_0_588), .ZN(n_8_0_2851));
   OAI211_X1 i_8_0_2806 (.A(n_8_0_2853), .B(n_8_0_3227), .C1(n_8_0_6166), 
      .C2(n_8_0_6824), .ZN(n_8_0_2852));
   OAI211_X1 i_8_0_2807 (.A(n_8_0_3186), .B(n_8_0_2854), .C1(n_8_0_6165), 
      .C2(n_8_0_3226), .ZN(n_8_0_2853));
   NAND2_X1 i_8_0_2808 (.A1(n_8_0_2854), .A2(n_8_0_7028), .ZN(n_8_0_1237));
   INV_X1 i_8_0_2809 (.A(n_8_0_2854), .ZN(n_8_0_1238));
   NOR2_X1 i_8_0_2810 (.A1(\out_as[5] [3]), .A2(n_8_0_584), .ZN(n_8_0_2854));
   AOI21_X1 i_8_0_2811 (.A(n_8_0_2856), .B1(n_8_0_6730), .B2(n_8_0_2857), 
      .ZN(n_8_0_2855));
   NOR2_X1 i_8_0_2812 (.A1(n_8_0_2858), .A2(n_8_0_2859), .ZN(n_8_0_2856));
   NAND2_X1 i_8_0_2813 (.A1(n_8_0_2858), .A2(n_8_0_2859), .ZN(n_8_0_2857));
   NAND2_X1 i_8_0_2814 (.A1(n_8_0_6157), .A2(n_8_0_3244), .ZN(n_8_0_2858));
   NOR2_X1 i_8_0_2815 (.A1(n_8_0_3211), .A2(n_8_0_1240), .ZN(n_8_0_2859));
   OR2_X1 i_8_0_2816 (.A1(n_8_0_1296), .A2(n_8_0_576), .ZN(n_8_0_1239));
   OR2_X1 i_8_0_2817 (.A1(\out_as[7] [3]), .A2(n_8_0_576), .ZN(n_8_0_1240));
   AOI22_X1 i_8_0_2818 (.A1(n_8_0_2861), .A2(n_8_0_2974), .B1(n_8_0_3189), 
      .B2(n_8_0_2862), .ZN(n_8_0_2860));
   AOI22_X1 i_8_0_2819 (.A1(n_8_0_596), .A2(n_8_0_6772), .B1(n_8_0_3020), 
      .B2(n_8_0_7056), .ZN(n_8_0_2861));
   INV_X1 i_8_0_2820 (.A(n_8_0_2862), .ZN(n_8_0_1241));
   NOR2_X1 i_8_0_2821 (.A1(\out_as[2] [3]), .A2(n_8_0_596), .ZN(n_8_0_2862));
   OAI211_X1 i_8_0_2822 (.A(n_8_0_2864), .B(n_8_0_2868), .C1(n_8_0_2869), 
      .C2(n_8_0_6811), .ZN(n_8_0_2863));
   AOI22_X1 i_8_0_2823 (.A1(n_8_0_3195), .A2(n_8_0_2865), .B1(n_8_0_2867), 
      .B2(n_8_0_6781), .ZN(n_8_0_2864));
   AOI21_X1 i_8_0_2824 (.A(n_8_0_1242), .B1(n_8_0_6784), .B2(n_8_0_2866), 
      .ZN(n_8_0_2865));
   INV_X1 i_8_0_2825 (.A(n_8_0_2867), .ZN(n_8_0_2866));
   NAND2_X1 i_8_0_2826 (.A1(n_8_0_5622), .A2(n_8_0_4325), .ZN(n_8_0_2867));
   OR2_X1 i_8_0_2827 (.A1(\out_as[1] [3]), .A2(n_8_0_600), .ZN(n_8_0_1242));
   OAI211_X1 i_8_0_2828 (.A(n_8_0_3207), .B(n_8_0_2870), .C1(n_8_0_3015), 
      .C2(\out_bs[0] [2]), .ZN(n_8_0_2868));
   AOI211_X1 i_8_0_2829 (.A(\out_bs[0] [2]), .B(n_8_0_3015), .C1(n_8_0_2870), 
      .C2(n_8_0_3207), .ZN(n_8_0_2869));
   NAND2_X1 i_8_0_2830 (.A1(n_8_0_3208), .A2(n_8_0_2870), .ZN(n_8_0_1243));
   INV_X1 i_8_0_2831 (.A(n_8_0_2870), .ZN(n_8_0_1244));
   NOR2_X1 i_8_0_2832 (.A1(\out_as[0] [3]), .A2(n_8_0_604), .ZN(n_8_0_2870));
   OAI22_X1 i_8_0_2833 (.A1(n_8_0_2873), .A2(n_8_0_2872), .B1(n_8_0_5455), 
      .B2(n_8_0_4728), .ZN(n_8_0_2871));
   AOI21_X1 i_8_0_2834 (.A(n_8_0_6755), .B1(n_8_0_5626), .B2(n_8_0_4563), 
      .ZN(n_8_0_2872));
   NOR2_X1 i_8_0_2835 (.A1(n_8_0_3203), .A2(n_8_0_1247), .ZN(n_8_0_2873));
   OR2_X1 i_8_0_2836 (.A1(n_8_0_1271), .A2(n_8_0_580), .ZN(n_8_0_1245));
   OR2_X1 i_8_0_2837 (.A1(n_8_0_1291), .A2(n_8_0_580), .ZN(n_8_0_1246));
   OR2_X1 i_8_0_2838 (.A1(\out_as[6] [3]), .A2(n_8_0_580), .ZN(n_8_0_1247));
   INV_X1 i_8_0_2839 (.A(n_8_0_2875), .ZN(n_8_0_2874));
   OAI21_X1 i_8_0_2840 (.A(n_8_0_2876), .B1(n_8_0_2877), .B2(n_8_0_2879), 
      .ZN(n_8_0_2875));
   NAND3_X1 i_8_0_2841 (.A1(n_8_0_6838), .A2(n_8_0_3181), .A3(n_8_0_2878), 
      .ZN(n_8_0_2876));
   AOI21_X1 i_8_0_2842 (.A(n_8_0_6838), .B1(n_8_0_3181), .B2(n_8_0_2878), 
      .ZN(n_8_0_2877));
   NAND3_X1 i_8_0_2843 (.A1(n_8_0_2878), .A2(n_8_0_7051), .A3(n_8_0_7052), 
      .ZN(n_8_0_1248));
   NAND2_X1 i_8_0_2844 (.A1(n_8_0_2878), .A2(n_8_0_7051), .ZN(n_8_0_1249));
   INV_X1 i_8_0_2845 (.A(n_8_0_2878), .ZN(n_8_0_1250));
   NOR2_X1 i_8_0_2846 (.A1(\out_as[3] [3]), .A2(n_8_0_592), .ZN(n_8_0_2878));
   NOR2_X1 i_8_0_2847 (.A1(n_8_0_3001), .A2(\out_bs[3] [2]), .ZN(n_8_0_2879));
   AOI21_X1 i_8_0_2848 (.A(n_8_0_6853), .B1(n_8_0_2881), .B2(n_8_0_2880), 
      .ZN(n_115));
   NOR3_X1 i_8_0_2849 (.A1(n_8_0_2909), .A2(n_8_0_2906), .A3(n_8_0_2883), 
      .ZN(n_8_0_2880));
   NOR4_X1 i_8_0_2850 (.A1(n_8_0_2896), .A2(n_8_0_2890), .A3(n_8_0_2882), 
      .A4(n_8_0_2901), .ZN(n_8_0_2881));
   OAI211_X1 i_8_0_2851 (.A(n_8_0_2913), .B(n_8_0_4132), .C1(n_8_0_5653), 
      .C2(n_8_0_6811), .ZN(n_8_0_2882));
   OAI21_X1 i_8_0_2852 (.A(n_8_0_2886), .B1(n_8_0_2884), .B2(n_8_0_3206), 
      .ZN(n_8_0_2883));
   OAI21_X1 i_8_0_2853 (.A(n_8_0_2885), .B1(n_8_0_3003), .B2(n_8_0_6522), 
      .ZN(n_8_0_2884));
   INV_X1 i_8_0_2854 (.A(n_8_0_2885), .ZN(n_8_0_1251));
   NOR2_X1 i_8_0_2855 (.A1(\out_as[0] [3]), .A2(n_8_0_572), .ZN(n_8_0_2885));
   AOI21_X1 i_8_0_2856 (.A(n_8_0_2887), .B1(n_8_0_2889), .B2(n_8_0_6794), 
      .ZN(n_8_0_2886));
   NOR2_X1 i_8_0_2857 (.A1(n_8_0_2888), .A2(n_8_0_556), .ZN(n_8_0_2887));
   OAI21_X1 i_8_0_2858 (.A(n_8_0_2987), .B1(n_8_0_3221), .B2(n_8_0_6191), 
      .ZN(n_8_0_2888));
   NAND2_X1 i_8_0_2859 (.A1(n_8_0_6192), .A2(n_8_0_3223), .ZN(n_8_0_2889));
   OR2_X1 i_8_0_2860 (.A1(\out_as[4] [3]), .A2(n_8_0_556), .ZN(n_8_0_1252));
   OAI21_X1 i_8_0_2861 (.A(n_8_0_2891), .B1(n_8_0_2892), .B2(n_8_0_2895), 
      .ZN(n_8_0_2890));
   NAND3_X1 i_8_0_2862 (.A1(n_8_0_6838), .A2(n_8_0_3181), .A3(n_8_0_2894), 
      .ZN(n_8_0_2891));
   AOI21_X1 i_8_0_2863 (.A(n_8_0_6838), .B1(n_8_0_3181), .B2(n_8_0_2894), 
      .ZN(n_8_0_2892));
   NAND3_X1 i_8_0_2864 (.A1(n_8_0_2894), .A2(n_8_0_7051), .A3(n_8_0_7052), 
      .ZN(n_8_0_1253));
   INV_X1 i_8_0_2865 (.A(n_8_0_2893), .ZN(n_8_0_1254));
   NOR2_X1 i_8_0_2866 (.A1(n_8_0_1353), .A2(\out_as[3] [3]), .ZN(n_8_0_2893));
   NAND2_X1 i_8_0_2867 (.A1(n_8_0_2894), .A2(n_8_0_7051), .ZN(n_8_0_1255));
   INV_X1 i_8_0_2868 (.A(n_8_0_2894), .ZN(n_8_0_1256));
   NOR2_X1 i_8_0_2869 (.A1(\out_as[3] [3]), .A2(n_8_0_560), .ZN(n_8_0_2894));
   NOR2_X1 i_8_0_2870 (.A1(n_8_0_6565), .A2(n_8_0_3001), .ZN(n_8_0_2895));
   AOI21_X1 i_8_0_2871 (.A(n_8_0_2897), .B1(n_8_0_2898), .B2(n_8_0_6824), 
      .ZN(n_8_0_2896));
   NOR3_X1 i_8_0_2872 (.A1(n_8_0_2899), .A2(n_8_0_3270), .A3(n_8_0_6210), 
      .ZN(n_8_0_2897));
   OAI21_X1 i_8_0_2873 (.A(n_8_0_2899), .B1(n_8_0_3270), .B2(n_8_0_6210), 
      .ZN(n_8_0_2898));
   NOR2_X1 i_8_0_2874 (.A1(n_8_0_3185), .A2(n_8_0_1258), .ZN(n_8_0_2899));
   OR2_X1 i_8_0_2875 (.A1(n_8_0_1289), .A2(n_8_0_552), .ZN(n_8_0_1257));
   OR2_X1 i_8_0_2876 (.A1(\out_as[5] [3]), .A2(n_8_0_552), .ZN(n_8_0_1258));
   INV_X1 i_8_0_2877 (.A(n_8_0_2901), .ZN(n_8_0_2900));
   OAI21_X1 i_8_0_2878 (.A(n_8_0_2902), .B1(n_8_0_2904), .B2(n_8_0_6755), 
      .ZN(n_8_0_2901));
   OAI211_X1 i_8_0_2879 (.A(n_8_0_3647), .B(n_8_0_2903), .C1(n_8_0_6757), 
      .C2(n_8_0_2905), .ZN(n_8_0_2902));
   NAND2_X1 i_8_0_2880 (.A1(n_8_0_2903), .A2(n_8_0_7017), .ZN(n_8_0_1259));
   INV_X1 i_8_0_2881 (.A(n_8_0_1260), .ZN(n_8_0_2903));
   OR2_X1 i_8_0_2882 (.A1(n_8_0_1291), .A2(n_8_0_548), .ZN(n_8_0_1260));
   OR2_X1 i_8_0_2883 (.A1(\out_as[6] [3]), .A2(n_8_0_548), .ZN(n_8_0_1261));
   INV_X1 i_8_0_2884 (.A(n_8_0_2905), .ZN(n_8_0_2904));
   NAND2_X1 i_8_0_2885 (.A1(n_8_0_6198), .A2(n_8_0_3237), .ZN(n_8_0_2905));
   AOI22_X1 i_8_0_2886 (.A1(n_8_0_2908), .A2(n_8_0_2907), .B1(n_8_0_5652), 
      .B2(n_8_0_3692), .ZN(n_8_0_2906));
   OAI21_X1 i_8_0_2887 (.A(n_8_0_6729), .B1(n_8_0_6201), .B2(n_8_0_3243), 
      .ZN(n_8_0_2907));
   OR2_X1 i_8_0_2888 (.A1(n_8_0_3211), .A2(n_8_0_1262), .ZN(n_8_0_2908));
   OR2_X1 i_8_0_2889 (.A1(\out_as[7] [3]), .A2(n_8_0_544), .ZN(n_8_0_1262));
   AOI22_X1 i_8_0_2890 (.A1(n_8_0_2912), .A2(n_8_0_2910), .B1(n_8_0_6537), 
      .B2(n_8_0_3019), .ZN(n_8_0_2909));
   NAND3_X1 i_8_0_2891 (.A1(n_8_0_3641), .A2(n_8_0_2911), .A3(n_8_0_7064), 
      .ZN(n_8_0_2910));
   NAND2_X1 i_8_0_2892 (.A1(n_8_0_2911), .A2(n_8_0_7064), .ZN(n_8_0_1263));
   INV_X1 i_8_0_2893 (.A(n_8_0_2911), .ZN(n_8_0_1264));
   NOR2_X1 i_8_0_2894 (.A1(\out_as[2] [3]), .A2(n_8_0_564), .ZN(n_8_0_2911));
   OAI21_X1 i_8_0_2895 (.A(n_8_0_6773), .B1(n_8_0_5642), .B2(n_8_0_4366), 
      .ZN(n_8_0_2912));
   OAI21_X1 i_8_0_2896 (.A(n_8_0_2914), .B1(n_8_0_6781), .B2(n_8_0_2915), 
      .ZN(n_8_0_2913));
   OAI21_X1 i_8_0_2897 (.A(n_8_0_2916), .B1(n_8_0_1267), .B2(n_8_0_3194), 
      .ZN(n_8_0_2914));
   NOR3_X1 i_8_0_2898 (.A1(n_8_0_2916), .A2(n_8_0_1267), .A3(n_8_0_3194), 
      .ZN(n_8_0_2915));
   NOR2_X1 i_8_0_2899 (.A1(n_8_0_5647), .A2(n_8_0_4324), .ZN(n_8_0_2916));
   NAND3_X1 i_8_0_2900 (.A1(n_8_0_2917), .A2(n_8_0_7076), .A3(n_8_0_7077), 
      .ZN(n_8_0_1265));
   NAND2_X1 i_8_0_2901 (.A1(n_8_0_2917), .A2(n_8_0_7076), .ZN(n_8_0_1266));
   INV_X1 i_8_0_2902 (.A(n_8_0_2917), .ZN(n_8_0_1267));
   NOR2_X1 i_8_0_2903 (.A1(\out_as[1] [3]), .A2(n_8_0_568), .ZN(n_8_0_2917));
   OAI22_X1 i_8_0_2908 (.A1(n_8_0_2923), .A2(n_8_0_2922), .B1(n_8_0_5690), 
      .B2(n_8_0_4384), .ZN(n_8_0_2921));
   NOR2_X1 i_8_0_2909 (.A1(n_8_0_3199), .A2(n_8_0_1269), .ZN(n_8_0_2922));
   OR2_X1 i_8_0_2910 (.A1(n_8_0_1297), .A2(n_8_0_520), .ZN(n_8_0_1268));
   OR2_X1 i_8_0_2911 (.A1(\out_as[4] [3]), .A2(n_8_0_520), .ZN(n_8_0_1269));
   AOI21_X1 i_8_0_2912 (.A(n_8_0_6795), .B1(n_8_0_6245), .B2(n_8_0_3223), 
      .ZN(n_8_0_2923));
   OAI33_X1 i_8_0_2913 (.A1(n_8_0_6759), .A2(n_8_0_6757), .A3(n_8_0_2926), 
      .B1(n_8_0_2925), .B2(n_8_0_5677), .B3(n_8_0_4562), .ZN(n_8_0_2924));
   NOR3_X1 i_8_0_2914 (.A1(\out_as[6] [6]), .A2(n_8_0_6763), .A3(n_8_0_1270), 
      .ZN(n_8_0_2925));
   NOR2_X1 i_8_0_2915 (.A1(n_8_0_3203), .A2(n_8_0_1273), .ZN(n_8_0_2926));
   NAND2_X1 i_8_0_2916 (.A1(n_8_0_3204), .A2(n_8_0_2927), .ZN(n_8_0_1270));
   NAND2_X1 i_8_0_2917 (.A1(n_8_0_3204), .A2(n_8_0_7015), .ZN(n_8_0_1271));
   NAND2_X1 i_8_0_2918 (.A1(n_8_0_2927), .A2(n_8_0_7016), .ZN(n_8_0_1272));
   INV_X1 i_8_0_2919 (.A(n_8_0_2927), .ZN(n_8_0_1273));
   NOR2_X1 i_8_0_2920 (.A1(\out_as[6] [3]), .A2(n_8_0_510), .ZN(n_8_0_2927));
   NAND2_X1 i_8_0_2922 (.A1(n_8_0_6824), .A2(n_8_0_2931), .ZN(n_8_0_2929));
   OAI21_X1 i_8_0_2923 (.A(n_8_0_3271), .B1(n_8_0_6831), .B2(n_8_0_2931), 
      .ZN(n_8_0_2930));
   NAND2_X1 i_8_0_2924 (.A1(n_8_0_3186), .A2(n_8_0_2932), .ZN(n_8_0_2931));
   NAND3_X1 i_8_0_2925 (.A1(n_8_0_2932), .A2(n_8_0_7028), .A3(n_8_0_7029), 
      .ZN(n_8_0_1274));
   NAND2_X1 i_8_0_2926 (.A1(n_8_0_2932), .A2(n_8_0_7028), .ZN(n_8_0_1275));
   INV_X1 i_8_0_2927 (.A(n_8_0_2932), .ZN(n_8_0_1276));
   NOR2_X1 i_8_0_2928 (.A1(\out_as[5] [3]), .A2(n_8_0_515), .ZN(n_8_0_2932));
   OAI211_X1 i_8_0_2929 (.A(n_8_0_3207), .B(n_8_0_2934), .C1(n_8_0_3003), 
      .C2(n_8_0_6668), .ZN(n_8_0_2933));
   OR2_X1 i_8_0_2930 (.A1(n_8_0_1295), .A2(n_8_0_540), .ZN(n_8_0_1277));
   INV_X1 i_8_0_2931 (.A(n_8_0_2934), .ZN(n_8_0_1278));
   NOR2_X1 i_8_0_2932 (.A1(\out_as[0] [3]), .A2(n_8_0_540), .ZN(n_8_0_2934));
   OAI21_X1 i_8_0_2934 (.A(n_8_0_4325), .B1(n_8_0_3194), .B2(n_8_0_1281), 
      .ZN(n_8_0_2936));
   AOI211_X1 i_8_0_2935 (.A(n_8_0_3194), .B(n_8_0_1281), .C1(n_8_0_5669), 
      .C2(n_8_0_4325), .ZN(n_8_0_2937));
   NAND3_X1 i_8_0_2936 (.A1(n_8_0_2938), .A2(n_8_0_7076), .A3(n_8_0_7077), 
      .ZN(n_8_0_1279));
   NAND2_X1 i_8_0_2937 (.A1(n_8_0_2938), .A2(n_8_0_7076), .ZN(n_8_0_1280));
   INV_X1 i_8_0_2938 (.A(n_8_0_2938), .ZN(n_8_0_1281));
   NOR2_X1 i_8_0_2939 (.A1(\out_as[1] [3]), .A2(n_8_0_535), .ZN(n_8_0_2938));
   OAI21_X1 i_8_0_2941 (.A(n_8_0_2942), .B1(n_8_0_4366), .B2(n_8_0_5664), 
      .ZN(n_8_0_2940));
   NOR3_X1 i_8_0_2942 (.A1(n_8_0_2942), .A2(n_8_0_4366), .A3(n_8_0_5664), 
      .ZN(n_8_0_2941));
   NOR2_X1 i_8_0_2943 (.A1(n_8_0_3190), .A2(n_8_0_1284), .ZN(n_8_0_2942));
   OR2_X1 i_8_0_2944 (.A1(n_8_0_1355), .A2(n_8_0_1284), .ZN(n_8_0_1282));
   OR2_X1 i_8_0_2945 (.A1(n_8_0_1293), .A2(n_8_0_530), .ZN(n_8_0_1283));
   OR2_X1 i_8_0_2946 (.A1(\out_as[2] [3]), .A2(n_8_0_530), .ZN(n_8_0_1284));
   OAI21_X1 i_8_0_2949 (.A(n_8_0_6729), .B1(n_8_0_6237), .B2(n_8_0_3243), 
      .ZN(n_8_0_2945));
   OR2_X1 i_8_0_2950 (.A1(n_8_0_1296), .A2(n_8_0_505), .ZN(n_8_0_1285));
   OR2_X1 i_8_0_2951 (.A1(\out_as[7] [3]), .A2(n_8_0_505), .ZN(n_8_0_1286));
   AOI21_X1 i_8_0_2953 (.A(n_8_0_2948), .B1(n_8_0_6838), .B2(n_8_0_2949), 
      .ZN(n_8_0_2947));
   NOR3_X1 i_8_0_2954 (.A1(n_8_0_2950), .A2(n_8_0_1288), .A3(n_8_0_3180), 
      .ZN(n_8_0_2948));
   OAI21_X1 i_8_0_2955 (.A(n_8_0_2950), .B1(n_8_0_2961), .B2(n_8_0_525), 
      .ZN(n_8_0_2949));
   OR2_X1 i_8_0_2956 (.A1(n_8_0_1290), .A2(n_8_0_525), .ZN(n_8_0_1287));
   OR2_X1 i_8_0_2957 (.A1(\out_as[3] [3]), .A2(n_8_0_525), .ZN(n_8_0_1288));
   NOR2_X1 i_8_0_2958 (.A1(n_8_0_5687), .A2(n_8_0_3685), .ZN(n_8_0_2950));
   NOR2_X1 i_8_0_2959 (.A1(n_8_0_2951), .A2(n_8_0_6853), .ZN(n_116));
   NOR2_X1 i_8_0_2960 (.A1(n_8_0_2953), .A2(n_8_0_2952), .ZN(n_8_0_2951));
   NAND4_X1 i_8_0_2961 (.A1(n_8_0_2984), .A2(n_8_0_2979), .A3(n_8_0_2972), 
      .A4(n_8_0_2964), .ZN(n_8_0_2952));
   NAND4_X1 i_8_0_2962 (.A1(n_8_0_2955), .A2(n_8_0_2954), .A3(n_8_0_2967), 
      .A4(n_8_0_2959), .ZN(n_8_0_2953));
   OAI21_X1 i_8_0_2963 (.A(n_8_0_2971), .B1(n_8_0_6810), .B2(n_8_0_2976), 
      .ZN(n_8_0_2954));
   OAI22_X1 i_8_0_2964 (.A1(n_8_0_2957), .A2(n_8_0_2956), .B1(n_8_0_6299), 
      .B2(n_8_0_3226), .ZN(n_8_0_2955));
   AOI21_X1 i_8_0_2965 (.A(n_8_0_6824), .B1(n_8_0_6298), .B2(n_8_0_3271), 
      .ZN(n_8_0_2956));
   NOR2_X1 i_8_0_2966 (.A1(n_8_0_3664), .A2(n_8_0_1289), .ZN(n_8_0_2957));
   INV_X1 i_8_0_2967 (.A(n_8_0_2958), .ZN(n_8_0_1289));
   NOR2_X1 i_8_0_2968 (.A1(\out_as[5] [4]), .A2(\out_as[5] [3]), .ZN(n_8_0_2958));
   OAI21_X1 i_8_0_2969 (.A(n_8_0_2960), .B1(n_8_0_2962), .B2(n_8_0_6838), 
      .ZN(n_8_0_2959));
   OAI211_X1 i_8_0_2970 (.A(n_8_0_5696), .B(n_8_0_3686), .C1(n_8_0_2961), 
      .C2(n_8_0_6837), .ZN(n_8_0_2960));
   NAND2_X1 i_8_0_2971 (.A1(n_8_0_3677), .A2(n_8_0_2963), .ZN(n_8_0_2961));
   NOR2_X1 i_8_0_2972 (.A1(n_8_0_3676), .A2(n_8_0_1290), .ZN(n_8_0_2962));
   INV_X1 i_8_0_2973 (.A(n_8_0_2963), .ZN(n_8_0_1290));
   NOR2_X1 i_8_0_2974 (.A1(\out_as[3] [4]), .A2(\out_as[3] [3]), .ZN(n_8_0_2963));
   OAI22_X1 i_8_0_2975 (.A1(n_8_0_5722), .A2(n_8_0_4560), .B1(n_8_0_4346), 
      .B2(n_8_0_2965), .ZN(n_8_0_2964));
   OAI21_X1 i_8_0_2976 (.A(n_8_0_2966), .B1(n_8_0_3203), .B2(\out_as[6] [3]), 
      .ZN(n_8_0_2965));
   NAND2_X1 i_8_0_2977 (.A1(n_8_0_7016), .A2(n_8_0_7015), .ZN(n_8_0_1291));
   NAND2_X1 i_8_0_2978 (.A1(n_8_0_6754), .A2(n_8_0_5722), .ZN(n_8_0_2966));
   OAI21_X1 i_8_0_2979 (.A(n_8_0_2968), .B1(n_8_0_4198), .B2(n_8_0_5711), 
      .ZN(n_8_0_2967));
   OAI21_X1 i_8_0_2980 (.A(n_8_0_2969), .B1(n_8_0_3194), .B2(\out_as[1] [3]), 
      .ZN(n_8_0_2968));
   OAI21_X1 i_8_0_2981 (.A(n_8_0_6781), .B1(n_8_0_5711), .B2(n_8_0_4324), 
      .ZN(n_8_0_2969));
   INV_X1 i_8_0_2982 (.A(n_8_0_2970), .ZN(n_8_0_1292));
   NOR2_X1 i_8_0_2983 (.A1(\out_as[1] [4]), .A2(\out_as[1] [3]), .ZN(n_8_0_2970));
   OAI211_X1 i_8_0_2984 (.A(n_8_0_6665), .B(n_8_0_3016), .C1(n_8_0_1295), 
      .C2(n_8_0_3643), .ZN(n_8_0_2971));
   OAI21_X1 i_8_0_2985 (.A(n_8_0_2974), .B1(n_8_0_2975), .B2(n_8_0_2973), 
      .ZN(n_8_0_2972));
   NAND2_X1 i_8_0_2986 (.A1(n_8_0_5707), .A2(n_8_0_4367), .ZN(n_8_0_2973));
   OAI21_X1 i_8_0_2987 (.A(n_8_0_6772), .B1(n_8_0_3190), .B2(\out_as[2] [3]), 
      .ZN(n_8_0_2974));
   NOR3_X1 i_8_0_2988 (.A1(n_8_0_6774), .A2(n_8_0_3640), .A3(n_8_0_1293), 
      .ZN(n_8_0_2975));
   NAND2_X1 i_8_0_2989 (.A1(n_8_0_7064), .A2(n_8_0_7063), .ZN(n_8_0_1293));
   AOI211_X1 i_8_0_2990 (.A(n_8_0_3643), .B(n_8_0_1295), .C1(n_8_0_3016), 
      .C2(n_8_0_6665), .ZN(n_8_0_2976));
   INV_X1 i_8_0_2991 (.A(n_8_0_2977), .ZN(n_8_0_1294));
   NOR2_X1 i_8_0_2992 (.A1(n_8_0_1359), .A2(\out_as[0] [3]), .ZN(n_8_0_2977));
   INV_X1 i_8_0_2993 (.A(n_8_0_2978), .ZN(n_8_0_1295));
   NOR2_X1 i_8_0_2994 (.A1(\out_as[0] [4]), .A2(\out_as[0] [3]), .ZN(n_8_0_2978));
   INV_X1 i_8_0_2999 (.A(n_8_0_2983), .ZN(n_8_0_1296));
   NOR2_X1 i_8_0_3000 (.A1(\out_as[7] [4]), .A2(\out_as[7] [3]), .ZN(n_8_0_2983));
   OAI21_X1 i_8_0_3001 (.A(n_8_0_2985), .B1(n_8_0_6794), .B2(n_8_0_2987), 
      .ZN(n_8_0_2984));
   OAI211_X1 i_8_0_3002 (.A(n_8_0_6629), .B(n_8_0_2997), .C1(n_8_0_6801), 
      .C2(n_8_0_2986), .ZN(n_8_0_2985));
   NAND2_X1 i_8_0_3003 (.A1(n_8_0_3670), .A2(n_8_0_2988), .ZN(n_8_0_2986));
   NOR2_X1 i_8_0_3004 (.A1(n_8_0_3669), .A2(n_8_0_1297), .ZN(n_8_0_2987));
   INV_X1 i_8_0_3005 (.A(n_8_0_2988), .ZN(n_8_0_1297));
   NOR2_X1 i_8_0_3006 (.A1(\out_as[4] [4]), .A2(\out_as[4] [3]), .ZN(n_8_0_2988));
   OAI21_X1 i_8_0_3012 (.A(n_8_0_3186), .B1(n_8_0_3226), .B2(\out_bs[5] [3]), 
      .ZN(n_8_0_2993));
   OR2_X1 i_8_0_3013 (.A1(\out_as[5] [4]), .A2(n_8_0_686), .ZN(n_8_0_1298));
   INV_X1 i_8_0_3015 (.A(n_8_0_2996), .ZN(n_8_0_2995));
   AOI211_X1 i_8_0_3016 (.A(n_8_0_3199), .B(n_8_0_689), .C1(n_8_0_6795), 
      .C2(n_8_0_2997), .ZN(n_8_0_2996));
   OR2_X1 i_8_0_3017 (.A1(\out_as[4] [4]), .A2(n_8_0_689), .ZN(n_8_0_1299));
   NOR2_X1 i_8_0_3018 (.A1(n_8_0_5744), .A2(n_8_0_4486), .ZN(n_8_0_2997));
   NOR3_X1 i_8_0_3020 (.A1(n_8_0_3000), .A2(n_8_0_1301), .A3(n_8_0_3676), 
      .ZN(n_8_0_2999));
   OR2_X1 i_8_0_3021 (.A1(n_8_0_1353), .A2(n_8_0_692), .ZN(n_8_0_1300));
   OR2_X1 i_8_0_3022 (.A1(\out_as[3] [4]), .A2(n_8_0_692), .ZN(n_8_0_1301));
   NOR2_X1 i_8_0_3023 (.A1(n_8_0_6838), .A2(n_8_0_3001), .ZN(n_8_0_3000));
   NAND2_X1 i_8_0_3024 (.A1(n_8_0_6008), .A2(n_8_0_3686), .ZN(n_8_0_3001));
   OR2_X1 i_8_0_3026 (.A1(n_8_0_1359), .A2(n_8_0_701), .ZN(n_8_0_1302));
   OR2_X1 i_8_0_3027 (.A1(\out_as[0] [4]), .A2(n_8_0_701), .ZN(n_8_0_1303));
   AOI211_X1 i_8_0_3030 (.A(n_8_0_683), .B(n_8_0_3203), .C1(n_8_0_4561), 
      .C2(n_8_0_5894), .ZN(n_8_0_3005));
   AOI21_X1 i_8_0_3031 (.A(n_8_0_6755), .B1(n_8_0_5894), .B2(n_8_0_4563), 
      .ZN(n_8_0_3006));
   OR2_X1 i_8_0_3032 (.A1(\out_as[6] [4]), .A2(n_8_0_683), .ZN(n_8_0_1304));
   OAI21_X1 i_8_0_3036 (.A(n_8_0_6729), .B1(n_8_0_3243), .B2(\out_bs[7] [3]), 
      .ZN(n_8_0_3010));
   OR2_X1 i_8_0_3037 (.A1(\out_as[7] [4]), .A2(n_8_0_680), .ZN(n_8_0_1305));
   NOR2_X1 i_8_0_3039 (.A1(n_8_0_3194), .A2(n_8_0_698), .ZN(n_8_0_3012));
   OR2_X1 i_8_0_3040 (.A1(\out_as[1] [4]), .A2(n_8_0_698), .ZN(n_8_0_1306));
   AOI21_X1 i_8_0_3041 (.A(n_8_0_6782), .B1(n_8_0_5984), .B2(n_8_0_4325), 
      .ZN(n_8_0_3013));
   NAND2_X1 i_8_0_3043 (.A1(n_8_0_5944), .A2(n_8_0_4604), .ZN(n_8_0_3015));
   NOR2_X1 i_8_0_3044 (.A1(n_8_0_5943), .A2(n_8_0_4603), .ZN(n_8_0_3016));
   OAI21_X1 i_8_0_3045 (.A(n_8_0_3018), .B1(n_8_0_4834), .B2(n_8_0_5427), 
      .ZN(n_8_0_3017));
   OAI22_X1 i_8_0_3046 (.A1(n_8_0_6772), .A2(n_8_0_3020), .B1(n_8_0_3190), 
      .B2(n_8_0_695), .ZN(n_8_0_3018));
   OR2_X1 i_8_0_3047 (.A1(\out_as[2] [4]), .A2(n_8_0_695), .ZN(n_8_0_1307));
   NOR2_X1 i_8_0_3048 (.A1(n_8_0_5427), .A2(n_8_0_4834), .ZN(n_8_0_3019));
   NOR2_X1 i_8_0_3049 (.A1(n_8_0_5814), .A2(n_8_0_4366), .ZN(n_8_0_3020));
   AOI21_X1 i_8_0_3050 (.A(n_8_0_6853), .B1(n_8_0_3021), .B2(n_8_0_3035), 
      .ZN(n_117));
   AND4_X1 i_8_0_3051 (.A1(n_8_0_3038), .A2(n_8_0_3029), .A3(n_8_0_3022), 
      .A4(n_8_0_3045), .ZN(n_8_0_3021));
   NOR3_X1 i_8_0_3052 (.A1(n_8_0_3023), .A2(n_8_0_4133), .A3(n_8_0_3024), 
      .ZN(n_8_0_3022));
   OAI211_X1 i_8_0_3053 (.A(n_8_0_3031), .B(n_8_0_3026), .C1(n_8_0_677), 
      .C2(n_8_0_3041), .ZN(n_8_0_3023));
   INV_X1 i_8_0_3054 (.A(n_8_0_3025), .ZN(n_8_0_3024));
   AOI211_X1 i_8_0_3055 (.A(n_8_0_3044), .B(n_8_0_3043), .C1(n_8_0_6810), 
      .C2(n_8_0_5771), .ZN(n_8_0_3025));
   AOI21_X1 i_8_0_3056 (.A(n_8_0_3028), .B1(n_8_0_3027), .B2(n_8_0_3677), 
      .ZN(n_8_0_3026));
   AOI21_X1 i_8_0_3057 (.A(n_8_0_1308), .B1(n_8_0_3452), .B2(n_8_0_5788), 
      .ZN(n_8_0_3027));
   OR2_X1 i_8_0_3058 (.A1(\out_as[3] [4]), .A2(n_8_0_668), .ZN(n_8_0_1308));
   AOI21_X1 i_8_0_3059 (.A(n_8_0_6837), .B1(n_8_0_5788), .B2(n_8_0_3686), 
      .ZN(n_8_0_3028));
   OAI22_X1 i_8_0_3060 (.A1(n_8_0_3030), .A2(n_8_0_4059), .B1(n_8_0_6351), 
      .B2(n_8_0_3221), .ZN(n_8_0_3029));
   OAI22_X1 i_8_0_3061 (.A1(n_8_0_6795), .A2(n_8_0_5783), .B1(n_8_0_3199), 
      .B2(n_8_0_665), .ZN(n_8_0_3030));
   OR2_X1 i_8_0_3062 (.A1(\out_as[4] [4]), .A2(n_8_0_665), .ZN(n_8_0_1309));
   OAI21_X1 i_8_0_3063 (.A(n_8_0_3033), .B1(n_8_0_3032), .B2(n_8_0_3034), 
      .ZN(n_8_0_3031));
   NOR3_X1 i_8_0_3064 (.A1(n_8_0_6831), .A2(n_8_0_3664), .A3(n_8_0_1310), 
      .ZN(n_8_0_3032));
   OAI21_X1 i_8_0_3065 (.A(n_8_0_6824), .B1(n_8_0_3185), .B2(n_8_0_662), 
      .ZN(n_8_0_3033));
   NAND2_X1 i_8_0_3066 (.A1(n_8_0_5775), .A2(n_8_0_4110), .ZN(n_8_0_3034));
   OR2_X1 i_8_0_3067 (.A1(\out_as[5] [4]), .A2(n_8_0_662), .ZN(n_8_0_1310));
   OAI21_X1 i_8_0_3068 (.A(n_8_0_3036), .B1(n_8_0_3691), .B2(n_8_0_5763), 
      .ZN(n_8_0_3035));
   OAI21_X1 i_8_0_3069 (.A(n_8_0_3037), .B1(n_8_0_3211), .B2(n_8_0_656), 
      .ZN(n_8_0_3036));
   OR2_X1 i_8_0_3070 (.A1(\out_as[7] [4]), .A2(n_8_0_656), .ZN(n_8_0_1311));
   OAI21_X1 i_8_0_3071 (.A(n_8_0_6729), .B1(n_8_0_6362), .B2(n_8_0_3243), 
      .ZN(n_8_0_3037));
   NOR3_X1 i_8_0_3072 (.A1(n_8_0_4365), .A2(n_8_0_3040), .A3(n_8_0_3039), 
      .ZN(n_8_0_3038));
   NOR2_X1 i_8_0_3073 (.A1(n_8_0_6772), .A2(n_8_0_5779), .ZN(n_8_0_3039));
   AOI211_X1 i_8_0_3074 (.A(n_8_0_671), .B(n_8_0_3190), .C1(n_8_0_4127), 
      .C2(n_8_0_5779), .ZN(n_8_0_3040));
   OR2_X1 i_8_0_3075 (.A1(\out_as[2] [4]), .A2(n_8_0_671), .ZN(n_8_0_1312));
   OAI21_X1 i_8_0_3076 (.A(n_8_0_3207), .B1(n_8_0_3696), .B2(n_8_0_5771), 
      .ZN(n_8_0_3041));
   OR2_X1 i_8_0_3077 (.A1(\out_as[0] [4]), .A2(n_8_0_677), .ZN(n_8_0_1313));
   NOR2_X1 i_8_0_3078 (.A1(n_8_0_3044), .A2(n_8_0_3043), .ZN(n_8_0_3042));
   AOI211_X1 i_8_0_3079 (.A(n_8_0_674), .B(n_8_0_3194), .C1(n_8_0_4199), 
      .C2(n_8_0_5758), .ZN(n_8_0_3043));
   OR2_X1 i_8_0_3080 (.A1(\out_as[1] [4]), .A2(n_8_0_674), .ZN(n_8_0_1314));
   AOI21_X1 i_8_0_3081 (.A(n_8_0_6782), .B1(n_8_0_5758), .B2(n_8_0_4325), 
      .ZN(n_8_0_3044));
   OAI221_X1 i_8_0_3082 (.A(n_8_0_3201), .B1(n_8_0_3202), .B2(n_8_0_5767), 
      .C1(n_8_0_3046), .C2(n_8_0_6855), .ZN(n_8_0_3045));
   AOI21_X1 i_8_0_3083 (.A(n_8_0_6755), .B1(n_8_0_5768), .B2(n_8_0_4563), 
      .ZN(n_8_0_3046));
   AOI21_X1 i_8_0_3084 (.A(n_8_0_6853), .B1(n_8_0_3072), .B2(n_8_0_3047), 
      .ZN(n_118));
   NOR4_X1 i_8_0_3085 (.A1(n_8_0_3061), .A2(n_8_0_3058), .A3(n_8_0_3054), 
      .A4(n_8_0_3048), .ZN(n_8_0_3047));
   OAI211_X1 i_8_0_3086 (.A(n_8_0_3050), .B(n_8_0_3049), .C1(n_8_0_653), 
      .C2(n_8_0_3053), .ZN(n_8_0_3048));
   OAI21_X1 i_8_0_3087 (.A(n_8_0_6810), .B1(n_8_0_5805), .B2(n_8_0_4603), 
      .ZN(n_8_0_3049));
   OAI21_X1 i_8_0_3088 (.A(n_8_0_3051), .B1(n_8_0_3052), .B2(n_8_0_6233), 
      .ZN(n_8_0_3050));
   OAI211_X1 i_8_0_3089 (.A(n_8_0_3244), .B(n_8_0_6403), .C1(n_8_0_3211), 
      .C2(n_8_0_632), .ZN(n_8_0_3051));
   AOI211_X1 i_8_0_3090 (.A(n_8_0_3658), .B(n_8_0_1315), .C1(n_8_0_3244), 
      .C2(n_8_0_6403), .ZN(n_8_0_3052));
   OR2_X1 i_8_0_3091 (.A1(\out_as[7] [4]), .A2(n_8_0_632), .ZN(n_8_0_1315));
   OAI21_X1 i_8_0_3092 (.A(n_8_0_3207), .B1(n_8_0_3696), .B2(n_8_0_5805), 
      .ZN(n_8_0_3053));
   OR2_X1 i_8_0_3093 (.A1(\out_as[0] [4]), .A2(n_8_0_653), .ZN(n_8_0_1316));
   NAND2_X1 i_8_0_3094 (.A1(n_8_0_4231), .A2(n_8_0_3055), .ZN(n_8_0_3054));
   NAND2_X1 i_8_0_3095 (.A1(n_8_0_3057), .A2(n_8_0_3056), .ZN(n_8_0_3055));
   NAND2_X1 i_8_0_3096 (.A1(n_8_0_4199), .A2(n_8_0_5819), .ZN(n_8_0_3056));
   OAI22_X1 i_8_0_3097 (.A1(n_8_0_6782), .A2(n_8_0_5819), .B1(n_8_0_3194), 
      .B2(n_8_0_650), .ZN(n_8_0_3057));
   OR2_X1 i_8_0_3098 (.A1(\out_as[1] [4]), .A2(n_8_0_650), .ZN(n_8_0_1317));
   OAI211_X1 i_8_0_3099 (.A(n_8_0_3059), .B(n_8_0_4347), .C1(n_8_0_5823), 
      .C2(n_8_0_6755), .ZN(n_8_0_3058));
   INV_X1 i_8_0_3100 (.A(n_8_0_3060), .ZN(n_8_0_3059));
   AOI211_X1 i_8_0_3101 (.A(n_8_0_635), .B(n_8_0_3203), .C1(n_8_0_4561), 
      .C2(n_8_0_5823), .ZN(n_8_0_3060));
   OR2_X1 i_8_0_3102 (.A1(\out_as[6] [4]), .A2(n_8_0_635), .ZN(n_8_0_1318));
   NAND3_X1 i_8_0_3103 (.A1(n_8_0_3066), .A2(n_8_0_3062), .A3(n_8_0_3069), 
      .ZN(n_8_0_3061));
   OAI21_X1 i_8_0_3104 (.A(n_8_0_3063), .B1(n_8_0_3065), .B2(n_8_0_6794), 
      .ZN(n_8_0_3062));
   OAI22_X1 i_8_0_3105 (.A1(n_8_0_6795), .A2(n_8_0_3064), .B1(n_8_0_3199), 
      .B2(n_8_0_641), .ZN(n_8_0_3063));
   OR2_X1 i_8_0_3106 (.A1(\out_as[4] [4]), .A2(n_8_0_641), .ZN(n_8_0_1319));
   INV_X1 i_8_0_3107 (.A(n_8_0_3065), .ZN(n_8_0_3064));
   OR2_X1 i_8_0_3108 (.A1(n_8_0_6381), .A2(n_8_0_3222), .ZN(n_8_0_3065));
   OAI21_X1 i_8_0_3109 (.A(n_8_0_3067), .B1(n_8_0_4126), .B2(n_8_0_5813), 
      .ZN(n_8_0_3066));
   OAI21_X1 i_8_0_3110 (.A(n_8_0_3068), .B1(n_8_0_3190), .B2(n_8_0_647), 
      .ZN(n_8_0_3067));
   OR2_X1 i_8_0_3111 (.A1(\out_as[2] [4]), .A2(n_8_0_647), .ZN(n_8_0_1320));
   OAI21_X1 i_8_0_3112 (.A(n_8_0_6773), .B1(n_8_0_5813), .B2(n_8_0_4366), 
      .ZN(n_8_0_3068));
   OAI21_X1 i_8_0_3113 (.A(n_8_0_3071), .B1(n_8_0_3070), .B2(n_8_0_5793), 
      .ZN(n_8_0_3069));
   OAI21_X1 i_8_0_3114 (.A(n_8_0_3686), .B1(n_8_0_3179), .B2(n_8_0_644), 
      .ZN(n_8_0_3070));
   OAI21_X1 i_8_0_3115 (.A(n_8_0_6837), .B1(n_8_0_3180), .B2(n_8_0_644), 
      .ZN(n_8_0_3071));
   OR2_X1 i_8_0_3116 (.A1(\out_as[3] [4]), .A2(n_8_0_644), .ZN(n_8_0_1321));
   OAI211_X1 i_8_0_3117 (.A(n_8_0_3184), .B(n_8_0_3073), .C1(n_8_0_3183), 
      .C2(n_8_0_6409), .ZN(n_8_0_3072));
   OAI211_X1 i_8_0_3118 (.A(n_8_0_638), .B(n_8_0_3227), .C1(n_8_0_6408), 
      .C2(n_8_0_6824), .ZN(n_8_0_3073));
   NOR3_X1 i_8_0_3122 (.A1(n_8_0_3082), .A2(n_8_0_3078), .A3(n_8_0_3077), 
      .ZN(n_8_0_3076));
   AOI21_X1 i_8_0_3123 (.A(n_8_0_6811), .B1(n_8_0_5854), .B2(n_8_0_4604), 
      .ZN(n_8_0_3077));
   AOI211_X1 i_8_0_3124 (.A(n_8_0_629), .B(n_8_0_3206), .C1(n_8_0_3697), 
      .C2(n_8_0_5854), .ZN(n_8_0_3078));
   OR2_X1 i_8_0_3128 (.A1(\out_as[7] [4]), .A2(n_8_0_608), .ZN(n_8_0_1322));
   OR2_X1 i_8_0_3129 (.A1(\out_as[0] [4]), .A2(n_8_0_629), .ZN(n_8_0_1323));
   OAI211_X1 i_8_0_3130 (.A(n_8_0_4231), .B(n_8_0_3083), .C1(n_8_0_6782), 
      .C2(n_8_0_5849), .ZN(n_8_0_3082));
   INV_X1 i_8_0_3131 (.A(n_8_0_3084), .ZN(n_8_0_3083));
   AOI211_X1 i_8_0_3132 (.A(n_8_0_626), .B(n_8_0_3194), .C1(n_8_0_4199), 
      .C2(n_8_0_5849), .ZN(n_8_0_3084));
   OR2_X1 i_8_0_3133 (.A1(\out_as[1] [4]), .A2(n_8_0_626), .ZN(n_8_0_1324));
   AOI21_X1 i_8_0_3135 (.A(n_8_0_4366), .B1(n_8_0_3189), .B2(n_8_0_6856), 
      .ZN(n_8_0_3086));
   NAND2_X1 i_8_0_3136 (.A1(n_8_0_3191), .A2(n_8_0_6856), .ZN(n_8_0_1325));
   NAND2_X1 i_8_0_3137 (.A1(n_8_0_7064), .A2(n_8_0_6856), .ZN(n_8_0_1326));
   OAI211_X1 i_8_0_3138 (.A(n_8_0_3184), .B(n_8_0_3088), .C1(n_8_0_3183), 
      .C2(n_8_0_6460), .ZN(n_8_0_3087));
   OAI21_X1 i_8_0_3139 (.A(n_8_0_614), .B1(n_8_0_6824), .B2(n_8_0_3089), 
      .ZN(n_8_0_3088));
   NOR2_X1 i_8_0_3140 (.A1(n_8_0_6460), .A2(n_8_0_3270), .ZN(n_8_0_3089));
   AOI21_X1 i_8_0_3142 (.A(n_8_0_6755), .B1(n_8_0_5828), .B2(n_8_0_4563), 
      .ZN(n_8_0_3091));
   AOI21_X1 i_8_0_3143 (.A(n_8_0_1328), .B1(n_8_0_4561), .B2(n_8_0_5828), 
      .ZN(n_8_0_3092));
   OR2_X1 i_8_0_3144 (.A1(n_8_0_1358), .A2(n_8_0_611), .ZN(n_8_0_1327));
   OR2_X1 i_8_0_3145 (.A1(\out_as[6] [4]), .A2(n_8_0_611), .ZN(n_8_0_1328));
   AOI211_X1 i_8_0_3146 (.A(n_8_0_4059), .B(n_8_0_3094), .C1(n_8_0_6794), 
      .C2(n_8_0_5835), .ZN(n_8_0_3093));
   AOI211_X1 i_8_0_3147 (.A(n_8_0_617), .B(n_8_0_3199), .C1(n_8_0_4385), 
      .C2(n_8_0_5836), .ZN(n_8_0_3094));
   OR2_X1 i_8_0_3148 (.A1(\out_as[4] [4]), .A2(n_8_0_617), .ZN(n_8_0_1329));
   AOI211_X1 i_8_0_3150 (.A(n_8_0_620), .B(n_8_0_3180), .C1(n_8_0_3452), 
      .C2(n_8_0_5859), .ZN(n_8_0_3096));
   OR2_X1 i_8_0_3151 (.A1(\out_as[3] [4]), .A2(n_8_0_620), .ZN(n_8_0_1330));
   AOI21_X1 i_8_0_3152 (.A(n_8_0_6837), .B1(n_8_0_5859), .B2(n_8_0_3686), 
      .ZN(n_8_0_3097));
   OAI21_X1 i_8_0_3157 (.A(n_8_0_3207), .B1(n_8_0_3696), .B2(n_8_0_5942), 
      .ZN(n_8_0_3101));
   OR2_X1 i_8_0_3158 (.A1(\out_as[0] [4]), .A2(n_8_0_605), .ZN(n_8_0_1331));
   AOI211_X1 i_8_0_3160 (.A(n_8_0_581), .B(n_8_0_3203), .C1(n_8_0_4561), 
      .C2(n_8_0_5970), .ZN(n_8_0_3103));
   AOI21_X1 i_8_0_3161 (.A(n_8_0_6755), .B1(n_8_0_5970), .B2(n_8_0_4563), 
      .ZN(n_8_0_3104));
   OR2_X1 i_8_0_3162 (.A1(\out_as[6] [4]), .A2(n_8_0_581), .ZN(n_8_0_1332));
   NOR2_X1 i_8_0_3163 (.A1(n_8_0_3107), .A2(n_8_0_3106), .ZN(n_8_0_3105));
   AOI211_X1 i_8_0_3164 (.A(n_8_0_589), .B(n_8_0_3199), .C1(n_8_0_4385), 
      .C2(n_8_0_5871), .ZN(n_8_0_3106));
   AOI21_X1 i_8_0_3165 (.A(n_8_0_6795), .B1(n_8_0_6641), .B2(n_8_0_3223), 
      .ZN(n_8_0_3107));
   OR2_X1 i_8_0_3166 (.A1(\out_as[4] [4]), .A2(n_8_0_589), .ZN(n_8_0_1333));
   OAI21_X1 i_8_0_3167 (.A(n_8_0_3109), .B1(n_8_0_6781), .B2(n_8_0_3110), 
      .ZN(n_8_0_3108));
   OAI211_X1 i_8_0_3168 (.A(n_8_0_4325), .B(n_8_0_5980), .C1(n_8_0_1334), 
      .C2(n_8_0_3653), .ZN(n_8_0_3109));
   AOI211_X1 i_8_0_3169 (.A(n_8_0_3653), .B(n_8_0_1334), .C1(n_8_0_5980), 
      .C2(n_8_0_4325), .ZN(n_8_0_3110));
   OR2_X1 i_8_0_3170 (.A1(\out_as[1] [4]), .A2(n_8_0_601), .ZN(n_8_0_1334));
   AOI22_X1 i_8_0_3171 (.A1(n_8_0_3113), .A2(n_8_0_3112), .B1(n_8_0_3189), 
      .B2(n_8_0_6857), .ZN(n_8_0_3111));
   OAI21_X1 i_8_0_3172 (.A(n_8_0_6772), .B1(n_8_0_3190), .B2(n_8_0_597), 
      .ZN(n_8_0_3112));
   NAND2_X1 i_8_0_3173 (.A1(n_8_0_7064), .A2(n_8_0_6857), .ZN(n_8_0_1335));
   NAND2_X1 i_8_0_3174 (.A1(n_8_0_5991), .A2(n_8_0_4367), .ZN(n_8_0_3113));
   NAND2_X1 i_8_0_3178 (.A1(n_8_0_7004), .A2(n_8_0_6859), .ZN(n_8_0_1336));
   OAI22_X1 i_8_0_3180 (.A1(n_8_0_3119), .A2(n_8_0_3684), .B1(n_8_0_5864), 
      .B2(n_8_0_3675), .ZN(n_8_0_3118));
   OAI22_X1 i_8_0_3181 (.A1(n_8_0_6837), .A2(n_8_0_5865), .B1(n_8_0_3180), 
      .B2(n_8_0_593), .ZN(n_8_0_3119));
   OR2_X1 i_8_0_3182 (.A1(\out_as[3] [4]), .A2(n_8_0_593), .ZN(n_8_0_1337));
   INV_X1 i_8_0_3183 (.A(n_8_0_3121), .ZN(n_8_0_3120));
   OAI211_X1 i_8_0_3184 (.A(n_8_0_3184), .B(n_8_0_3122), .C1(n_8_0_3183), 
      .C2(n_8_0_6679), .ZN(n_8_0_3121));
   OAI211_X1 i_8_0_3185 (.A(n_8_0_585), .B(n_8_0_3227), .C1(n_8_0_6678), 
      .C2(n_8_0_6824), .ZN(n_8_0_3122));
   NOR3_X1 i_8_0_3189 (.A1(n_8_0_3134), .A2(n_8_0_3127), .A3(n_8_0_3126), 
      .ZN(n_8_0_3125));
   AOI211_X1 i_8_0_3190 (.A(n_8_0_573), .B(n_8_0_3206), .C1(n_8_0_3697), 
      .C2(n_8_0_5908), .ZN(n_8_0_3126));
   AOI21_X1 i_8_0_3191 (.A(n_8_0_6811), .B1(n_8_0_5908), .B2(n_8_0_4604), 
      .ZN(n_8_0_3127));
   AOI211_X1 i_8_0_3193 (.A(n_8_0_4059), .B(n_8_0_3130), .C1(n_8_0_6794), 
      .C2(n_8_0_5897), .ZN(n_8_0_3129));
   AOI211_X1 i_8_0_3194 (.A(n_8_0_3199), .B(n_8_0_557), .C1(n_8_0_5460), 
      .C2(n_8_0_4976), .ZN(n_8_0_3130));
   OR2_X1 i_8_0_3195 (.A1(\out_as[4] [4]), .A2(n_8_0_557), .ZN(n_8_0_1338));
   NOR2_X1 i_8_0_3196 (.A1(n_8_0_3133), .A2(n_8_0_3132), .ZN(n_8_0_3131));
   AOI21_X1 i_8_0_3197 (.A(n_8_0_6755), .B1(n_8_0_5892), .B2(n_8_0_4563), 
      .ZN(n_8_0_3132));
   AOI211_X1 i_8_0_3198 (.A(n_8_0_549), .B(n_8_0_3203), .C1(n_8_0_4561), 
      .C2(n_8_0_5892), .ZN(n_8_0_3133));
   OR2_X1 i_8_0_3199 (.A1(\out_as[6] [4]), .A2(n_8_0_549), .ZN(n_8_0_1339));
   OAI211_X1 i_8_0_3200 (.A(n_8_0_4231), .B(n_8_0_3135), .C1(n_8_0_6782), 
      .C2(n_8_0_5901), .ZN(n_8_0_3134));
   INV_X1 i_8_0_3201 (.A(n_8_0_3136), .ZN(n_8_0_3135));
   AOI211_X1 i_8_0_3202 (.A(n_8_0_569), .B(n_8_0_3194), .C1(n_8_0_4199), 
      .C2(n_8_0_5901), .ZN(n_8_0_3136));
   OR2_X1 i_8_0_3203 (.A1(\out_as[1] [4]), .A2(n_8_0_569), .ZN(n_8_0_1340));
   AOI211_X1 i_8_0_3204 (.A(n_8_0_4365), .B(n_8_0_3138), .C1(n_8_0_6773), 
      .C2(n_8_0_5905), .ZN(n_8_0_3137));
   AOI211_X1 i_8_0_3205 (.A(n_8_0_3190), .B(n_8_0_565), .C1(n_8_0_5428), 
      .C2(n_8_0_4963), .ZN(n_8_0_3138));
   OR2_X1 i_8_0_3206 (.A1(\out_as[2] [4]), .A2(n_8_0_565), .ZN(n_8_0_1341));
   OR2_X1 i_8_0_3207 (.A1(\out_as[0] [4]), .A2(n_8_0_573), .ZN(n_8_0_1342));
   OR2_X1 i_8_0_3211 (.A1(\out_as[7] [4]), .A2(n_8_0_545), .ZN(n_8_0_1343));
   OAI221_X1 i_8_0_3213 (.A(n_8_0_3686), .B1(n_8_0_5918), .B2(n_8_0_6008), 
      .C1(n_8_0_3179), .C2(n_8_0_561), .ZN(n_8_0_3143));
   OAI21_X1 i_8_0_3214 (.A(n_8_0_6837), .B1(n_8_0_3180), .B2(n_8_0_561), 
      .ZN(n_8_0_3144));
   OR2_X1 i_8_0_3215 (.A1(\out_as[3] [4]), .A2(n_8_0_561), .ZN(n_8_0_1344));
   OAI211_X1 i_8_0_3217 (.A(n_8_0_553), .B(n_8_0_3227), .C1(n_8_0_6515), 
      .C2(n_8_0_6824), .ZN(n_8_0_3146));
   AOI21_X1 i_8_0_3218 (.A(n_8_0_6853), .B1(n_8_0_3171), .B2(n_8_0_3147), 
      .ZN(n_119));
   NOR2_X1 i_8_0_3219 (.A1(n_8_0_3155), .A2(n_8_0_3148), .ZN(n_8_0_3147));
   NAND3_X1 i_8_0_3220 (.A1(n_8_0_3149), .A2(n_8_0_3165), .A3(n_8_0_3163), 
      .ZN(n_8_0_3148));
   NOR4_X1 i_8_0_3221 (.A1(n_8_0_3153), .A2(n_8_0_3168), .A3(n_8_0_3159), 
      .A4(n_8_0_3150), .ZN(n_8_0_3149));
   OAI21_X1 i_8_0_3222 (.A(n_8_0_3152), .B1(n_8_0_3151), .B2(n_8_0_541), 
      .ZN(n_8_0_3150));
   OAI21_X1 i_8_0_3223 (.A(n_8_0_3207), .B1(n_8_0_3696), .B2(n_8_0_5940), 
      .ZN(n_8_0_3151));
   OAI21_X1 i_8_0_3224 (.A(n_8_0_6810), .B1(n_8_0_5940), .B2(n_8_0_4603), 
      .ZN(n_8_0_3152));
   OAI221_X1 i_8_0_3225 (.A(n_8_0_3803), .B1(n_8_0_5957), .B2(n_8_0_6824), 
      .C1(n_8_0_3154), .C2(n_8_0_516), .ZN(n_8_0_3153));
   OAI21_X1 i_8_0_3226 (.A(n_8_0_3186), .B1(n_8_0_3226), .B2(n_8_0_6676), 
      .ZN(n_8_0_3154));
   OR2_X1 i_8_0_3227 (.A1(\out_as[5] [4]), .A2(n_8_0_516), .ZN(n_8_0_1345));
   OAI21_X1 i_8_0_3228 (.A(n_8_0_3156), .B1(n_8_0_3157), .B2(n_8_0_6795), 
      .ZN(n_8_0_3155));
   OAI22_X1 i_8_0_3229 (.A1(n_8_0_6794), .A2(n_8_0_3158), .B1(n_8_0_3222), 
      .B2(n_8_0_6640), .ZN(n_8_0_3156));
   INV_X1 i_8_0_3230 (.A(n_8_0_3158), .ZN(n_8_0_3157));
   NOR2_X1 i_8_0_3231 (.A1(n_8_0_3199), .A2(n_8_0_521), .ZN(n_8_0_3158));
   OR2_X1 i_8_0_3232 (.A1(\out_as[4] [4]), .A2(n_8_0_521), .ZN(n_8_0_1346));
   OR2_X1 i_8_0_3233 (.A1(n_8_0_3161), .A2(n_8_0_3160), .ZN(n_8_0_3159));
   AOI211_X1 i_8_0_3234 (.A(n_8_0_526), .B(n_8_0_3180), .C1(n_8_0_3452), 
      .C2(n_8_0_5932), .ZN(n_8_0_3160));
   OR2_X1 i_8_0_3235 (.A1(\out_as[3] [4]), .A2(n_8_0_526), .ZN(n_8_0_1347));
   AOI21_X1 i_8_0_3236 (.A(n_8_0_6837), .B1(n_8_0_5932), .B2(n_8_0_3686), 
      .ZN(n_8_0_3161));
   INV_X1 i_8_0_3237 (.A(n_8_0_3163), .ZN(n_8_0_3162));
   AOI211_X1 i_8_0_3238 (.A(n_8_0_4346), .B(n_8_0_3164), .C1(n_8_0_6754), 
      .C2(n_8_0_5935), .ZN(n_8_0_3163));
   AOI211_X1 i_8_0_3239 (.A(n_8_0_511), .B(n_8_0_3203), .C1(n_8_0_4561), 
      .C2(n_8_0_5936), .ZN(n_8_0_3164));
   OR2_X1 i_8_0_3240 (.A1(\out_as[6] [4]), .A2(n_8_0_511), .ZN(n_8_0_1348));
   NAND2_X1 i_8_0_3241 (.A1(n_8_0_3167), .A2(n_8_0_3166), .ZN(n_8_0_3165));
   OAI21_X1 i_8_0_3242 (.A(n_8_0_6772), .B1(n_8_0_3190), .B2(n_8_0_531), 
      .ZN(n_8_0_3166));
   OAI211_X1 i_8_0_3243 (.A(n_8_0_5947), .B(n_8_0_4367), .C1(n_8_0_3638), 
      .C2(n_8_0_1349), .ZN(n_8_0_3167));
   OR2_X1 i_8_0_3244 (.A1(\out_as[2] [4]), .A2(n_8_0_531), .ZN(n_8_0_1349));
   OR2_X1 i_8_0_3245 (.A1(\out_as[0] [4]), .A2(n_8_0_541), .ZN(n_8_0_1350));
   AOI21_X1 i_8_0_3246 (.A(n_8_0_3169), .B1(n_8_0_4199), .B2(n_8_0_5961), 
      .ZN(n_8_0_3168));
   INV_X1 i_8_0_3247 (.A(n_8_0_3170), .ZN(n_8_0_3169));
   OAI221_X1 i_8_0_3248 (.A(n_8_0_4231), .B1(n_8_0_3194), .B2(n_8_0_536), 
      .C1(n_8_0_6782), .C2(n_8_0_5961), .ZN(n_8_0_3170));
   OR2_X1 i_8_0_3249 (.A1(\out_as[1] [4]), .A2(n_8_0_536), .ZN(n_8_0_1351));
   OAI21_X1 i_8_0_3250 (.A(n_8_0_3172), .B1(n_8_0_3691), .B2(n_8_0_5952), 
      .ZN(n_8_0_3171));
   OAI21_X1 i_8_0_3251 (.A(n_8_0_3173), .B1(n_8_0_3211), .B2(n_8_0_506), 
      .ZN(n_8_0_3172));
   OAI21_X1 i_8_0_3252 (.A(n_8_0_6729), .B1(n_8_0_5952), .B2(n_8_0_4423), 
      .ZN(n_8_0_3173));
   OR2_X1 i_8_0_3253 (.A1(\out_as[7] [4]), .A2(n_8_0_506), .ZN(n_8_0_1352));
   NAND3_X1 i_8_0_3259 (.A1(n_8_0_3179), .A2(n_8_0_3686), .A3(n_8_0_6006), 
      .ZN(n_8_0_3178));
   NAND2_X1 i_8_0_3260 (.A1(n_8_0_6841), .A2(n_8_0_3181), .ZN(n_8_0_3179));
   NAND2_X1 i_8_0_3261 (.A1(n_8_0_3677), .A2(n_8_0_7051), .ZN(n_8_0_3180));
   NOR2_X1 i_8_0_3262 (.A1(n_8_0_3676), .A2(\out_as[3] [4]), .ZN(n_8_0_3181));
   NAND2_X1 i_8_0_3263 (.A1(n_8_0_7052), .A2(n_8_0_7051), .ZN(n_8_0_1353));
   OAI21_X1 i_8_0_3264 (.A(n_8_0_3184), .B1(n_8_0_3183), .B2(n_8_0_6674), 
      .ZN(n_8_0_3182));
   OAI21_X1 i_8_0_3265 (.A(n_8_0_3271), .B1(n_8_0_3185), .B2(n_8_0_6824), 
      .ZN(n_8_0_3183));
   NAND2_X1 i_8_0_3266 (.A1(n_8_0_6824), .A2(n_8_0_3185), .ZN(n_8_0_3184));
   NAND2_X1 i_8_0_3267 (.A1(n_8_0_3665), .A2(n_8_0_7028), .ZN(n_8_0_3185));
   NOR2_X1 i_8_0_3268 (.A1(n_8_0_3664), .A2(\out_as[5] [4]), .ZN(n_8_0_3186));
   NAND2_X1 i_8_0_3269 (.A1(n_8_0_7029), .A2(n_8_0_7028), .ZN(n_8_0_1354));
   NOR3_X1 i_8_0_3271 (.A1(n_8_0_5989), .A2(n_8_0_3189), .A3(n_8_0_4366), 
      .ZN(n_8_0_3188));
   NOR2_X1 i_8_0_3272 (.A1(n_8_0_6772), .A2(n_8_0_3190), .ZN(n_8_0_3189));
   NAND2_X1 i_8_0_3273 (.A1(n_8_0_3641), .A2(n_8_0_7064), .ZN(n_8_0_3190));
   INV_X1 i_8_0_3274 (.A(n_8_0_3191), .ZN(n_8_0_1355));
   NOR2_X1 i_8_0_3275 (.A1(\out_as[2] [5]), .A2(\out_as[2] [4]), .ZN(n_8_0_3191));
   OAI22_X1 i_8_0_3276 (.A1(n_8_0_6781), .A2(n_8_0_3195), .B1(n_8_0_3193), 
      .B2(n_8_0_5979), .ZN(n_8_0_3192));
   OAI21_X1 i_8_0_3277 (.A(n_8_0_4325), .B1(n_8_0_6786), .B2(n_8_0_3194), 
      .ZN(n_8_0_3193));
   NAND2_X1 i_8_0_3278 (.A1(n_8_0_3654), .A2(n_8_0_7076), .ZN(n_8_0_3194));
   NOR2_X1 i_8_0_3279 (.A1(n_8_0_3653), .A2(\out_as[1] [4]), .ZN(n_8_0_3195));
   NAND2_X1 i_8_0_3280 (.A1(n_8_0_7077), .A2(n_8_0_7076), .ZN(n_8_0_1356));
   OAI211_X1 i_8_0_3282 (.A(n_8_0_5996), .B(n_8_0_4487), .C1(n_8_0_6795), 
      .C2(n_8_0_3199), .ZN(n_8_0_3197));
   NAND2_X1 i_8_0_3283 (.A1(n_8_0_6795), .A2(n_8_0_3199), .ZN(n_8_0_3198));
   NAND2_X1 i_8_0_3284 (.A1(n_8_0_3670), .A2(n_8_0_7039), .ZN(n_8_0_3199));
   OR2_X1 i_8_0_3285 (.A1(\out_as[4] [5]), .A2(\out_as[4] [4]), .ZN(n_8_0_1357));
   NAND2_X1 i_8_0_3287 (.A1(n_8_0_6755), .A2(n_8_0_3203), .ZN(n_8_0_3201));
   OAI21_X1 i_8_0_3288 (.A(n_8_0_4563), .B1(n_8_0_6763), .B2(n_8_0_3203), 
      .ZN(n_8_0_3202));
   NAND2_X1 i_8_0_3289 (.A1(n_8_0_3647), .A2(n_8_0_7016), .ZN(n_8_0_3203));
   INV_X1 i_8_0_3290 (.A(n_8_0_3204), .ZN(n_8_0_1358));
   NOR2_X1 i_8_0_3291 (.A1(\out_as[6] [5]), .A2(\out_as[6] [4]), .ZN(n_8_0_3204));
   NAND2_X1 i_8_0_3293 (.A1(n_8_0_3208), .A2(n_8_0_7089), .ZN(n_8_0_3206));
   NOR2_X1 i_8_0_3294 (.A1(n_8_0_3643), .A2(\out_as[0] [4]), .ZN(n_8_0_3207));
   INV_X1 i_8_0_3295 (.A(n_8_0_3208), .ZN(n_8_0_1359));
   NOR2_X1 i_8_0_3296 (.A1(\out_as[0] [5]), .A2(\out_as[0] [4]), .ZN(n_8_0_3208));
   OR2_X1 i_8_0_3301 (.A1(\out_as[7] [5]), .A2(\out_as[7] [4]), .ZN(n_8_0_1360));
   OAI21_X1 i_8_0_3306 (.A(n_8_0_3217), .B1(n_8_0_1361), .B2(n_8_0_4197), 
      .ZN(n_8_0_3216));
   OAI21_X1 i_8_0_3307 (.A(n_8_0_3218), .B1(n_8_0_4232), .B2(\out_bs[1] [4]), 
      .ZN(n_8_0_3217));
   OAI21_X1 i_8_0_3308 (.A(n_8_0_6782), .B1(n_8_0_3653), .B2(n_8_0_828), 
      .ZN(n_8_0_3218));
   OR2_X1 i_8_0_3309 (.A1(\out_as[1] [5]), .A2(n_8_0_828), .ZN(n_8_0_1361));
   OAI21_X1 i_8_0_3311 (.A(n_8_0_6622), .B1(n_8_0_3669), .B2(n_8_0_822), 
      .ZN(n_8_0_3220));
   OR2_X1 i_8_0_3312 (.A1(\out_as[4] [5]), .A2(n_8_0_822), .ZN(n_8_0_1362));
   NAND2_X1 i_8_0_3313 (.A1(n_8_0_6801), .A2(n_8_0_3223), .ZN(n_8_0_3221));
   NAND2_X1 i_8_0_3314 (.A1(n_8_0_5224), .A2(n_8_0_7035), .ZN(n_8_0_3222));
   NOR2_X1 i_8_0_3315 (.A1(n_8_0_5223), .A2(\out_bs[4] [6]), .ZN(n_8_0_3223));
   AND2_X1 i_8_0_3316 (.A1(n_8_0_3226), .A2(n_8_0_3225), .ZN(n_8_0_3224));
   OAI21_X1 i_8_0_3317 (.A(n_8_0_3227), .B1(n_8_0_3664), .B2(n_8_0_820), 
      .ZN(n_8_0_3225));
   NAND2_X1 i_8_0_3318 (.A1(n_8_0_6828), .A2(n_8_0_3271), .ZN(n_8_0_3226));
   NAND2_X1 i_8_0_3319 (.A1(n_8_0_6825), .A2(n_8_0_3270), .ZN(n_8_0_3227));
   OAI21_X1 i_8_0_3321 (.A(n_8_0_3686), .B1(n_8_0_3673), .B2(n_8_0_824), 
      .ZN(n_8_0_3229));
   OAI21_X1 i_8_0_3322 (.A(n_8_0_6837), .B1(n_8_0_3676), .B2(n_8_0_824), 
      .ZN(n_8_0_3230));
   OR2_X1 i_8_0_3323 (.A1(\out_as[3] [5]), .A2(n_8_0_824), .ZN(n_8_0_1363));
   OAI21_X1 i_8_0_3325 (.A(n_8_0_6772), .B1(n_8_0_3640), .B2(n_8_0_826), 
      .ZN(n_8_0_3232));
   NAND2_X1 i_8_0_3326 (.A1(n_8_0_7058), .A2(n_8_0_4364), .ZN(n_8_0_3233));
   NOR2_X1 i_8_0_3327 (.A1(n_8_0_4125), .A2(n_8_0_1364), .ZN(n_8_0_3234));
   OR2_X1 i_8_0_3328 (.A1(\out_as[2] [5]), .A2(n_8_0_826), .ZN(n_8_0_1364));
   OAI21_X1 i_8_0_3330 (.A(n_8_0_3647), .B1(n_8_0_4560), .B2(\out_bs[6] [4]), 
      .ZN(n_8_0_3236));
   NOR2_X1 i_8_0_3331 (.A1(n_8_0_4562), .A2(\out_bs[6] [4]), .ZN(n_8_0_3237));
   OR2_X1 i_8_0_3332 (.A1(\out_as[6] [5]), .A2(n_8_0_818), .ZN(n_8_0_1365));
   NOR2_X1 i_8_0_3335 (.A1(n_8_0_4603), .A2(\out_bs[0] [4]), .ZN(n_8_0_3240));
   OR2_X1 i_8_0_3338 (.A1(\out_as[7] [5]), .A2(n_8_0_816), .ZN(n_8_0_1366));
   AOI21_X1 i_8_0_3341 (.A(n_8_0_6853), .B1(n_8_0_3246), .B2(n_8_0_3245), 
      .ZN(n_120));
   NOR4_X1 i_8_0_3342 (.A1(n_8_0_3266), .A2(n_8_0_3263), .A3(n_8_0_3250), 
      .A4(n_8_0_3247), .ZN(n_8_0_3245));
   AND3_X1 i_8_0_3343 (.A1(n_8_0_3273), .A2(n_8_0_3256), .A3(n_8_0_3253), 
      .ZN(n_8_0_3246));
   OAI21_X1 i_8_0_3344 (.A(n_8_0_3248), .B1(n_8_0_6054), .B2(n_8_0_6811), 
      .ZN(n_8_0_3247));
   NOR3_X1 i_8_0_3345 (.A1(n_8_0_3259), .A2(n_8_0_3249), .A3(n_8_0_4133), 
      .ZN(n_8_0_3248));
   AOI211_X1 i_8_0_3346 (.A(n_8_0_814), .B(n_8_0_3643), .C1(n_8_0_3697), 
      .C2(n_8_0_6054), .ZN(n_8_0_3249));
   OAI211_X1 i_8_0_3347 (.A(n_8_0_3251), .B(n_8_0_3448), .C1(n_8_0_3451), 
      .C2(n_8_0_808), .ZN(n_8_0_3250));
   NAND2_X1 i_8_0_3348 (.A1(n_8_0_6357), .A2(n_8_0_3252), .ZN(n_8_0_3251));
   OAI21_X1 i_8_0_3349 (.A(n_8_0_4309), .B1(n_8_0_3402), .B2(n_8_0_808), 
      .ZN(n_8_0_3252));
   AOI211_X1 i_8_0_3350 (.A(n_8_0_4059), .B(n_8_0_3254), .C1(n_8_0_6623), 
      .C2(n_8_0_6031), .ZN(n_8_0_3253));
   NOR2_X1 i_8_0_3351 (.A1(n_8_0_806), .A2(n_8_0_3255), .ZN(n_8_0_3254));
   AOI21_X1 i_8_0_3352 (.A(n_8_0_3559), .B1(n_8_0_3406), .B2(n_8_0_6031), 
      .ZN(n_8_0_3255));
   NAND2_X1 i_8_0_3353 (.A1(n_8_0_3258), .A2(n_8_0_3257), .ZN(n_8_0_3256));
   OAI221_X1 i_8_0_3354 (.A(n_8_0_4424), .B1(n_8_0_6041), .B2(n_8_0_6998), 
      .C1(n_8_0_3657), .C2(n_8_0_800), .ZN(n_8_0_3257));
   OAI21_X1 i_8_0_3355 (.A(n_8_0_6730), .B1(n_8_0_3658), .B2(n_8_0_800), 
      .ZN(n_8_0_3258));
   OR2_X1 i_8_0_3356 (.A1(\out_as[7] [5]), .A2(n_8_0_800), .ZN(n_8_0_1367));
   OR2_X1 i_8_0_3357 (.A1(\out_as[0] [5]), .A2(n_8_0_814), .ZN(n_8_0_1368));
   INV_X1 i_8_0_3358 (.A(n_8_0_3260), .ZN(n_8_0_3259));
   NOR2_X1 i_8_0_3359 (.A1(n_8_0_3262), .A2(n_8_0_3261), .ZN(n_8_0_3260));
   AOI211_X1 i_8_0_3360 (.A(n_8_0_812), .B(n_8_0_3653), .C1(n_8_0_4199), 
      .C2(n_8_0_6049), .ZN(n_8_0_3261));
   OR2_X1 i_8_0_3361 (.A1(\out_as[1] [5]), .A2(n_8_0_812), .ZN(n_8_0_1369));
   AOI21_X1 i_8_0_3362 (.A(n_8_0_6782), .B1(n_8_0_6049), .B2(n_8_0_4325), 
      .ZN(n_8_0_3262));
   AND2_X1 i_8_0_3363 (.A1(n_8_0_3265), .A2(n_8_0_3264), .ZN(n_8_0_3263));
   OAI211_X1 i_8_0_3364 (.A(n_8_0_6046), .B(n_8_0_4367), .C1(n_8_0_3638), 
      .C2(n_8_0_810), .ZN(n_8_0_3264));
   OAI21_X1 i_8_0_3365 (.A(n_8_0_6772), .B1(n_8_0_3640), .B2(n_8_0_810), 
      .ZN(n_8_0_3265));
   OR2_X1 i_8_0_3366 (.A1(\out_as[2] [5]), .A2(n_8_0_810), .ZN(n_8_0_1370));
   AOI21_X1 i_8_0_3367 (.A(n_8_0_3267), .B1(n_8_0_6824), .B2(n_8_0_804), 
      .ZN(n_8_0_3266));
   OAI21_X1 i_8_0_3368 (.A(n_8_0_3663), .B1(n_8_0_3269), .B2(n_8_0_3268), 
      .ZN(n_8_0_3267));
   NOR2_X1 i_8_0_3369 (.A1(n_8_0_3662), .A2(n_8_0_804), .ZN(n_8_0_3268));
   NAND2_X1 i_8_0_3370 (.A1(n_8_0_6057), .A2(n_8_0_4110), .ZN(n_8_0_3269));
   NAND2_X1 i_8_0_3371 (.A1(n_8_0_4110), .A2(n_8_0_7022), .ZN(n_8_0_3270));
   NOR2_X1 i_8_0_3372 (.A1(n_8_0_4109), .A2(\out_bs[5] [4]), .ZN(n_8_0_3271));
   INV_X1 i_8_0_3373 (.A(n_8_0_3273), .ZN(n_8_0_3272));
   AOI211_X1 i_8_0_3374 (.A(n_8_0_4346), .B(n_8_0_3274), .C1(n_8_0_3275), 
      .C2(n_8_0_6035), .ZN(n_8_0_3273));
   NOR2_X1 i_8_0_3375 (.A1(n_8_0_4558), .A2(n_8_0_1371), .ZN(n_8_0_3274));
   OAI21_X1 i_8_0_3376 (.A(n_8_0_6755), .B1(n_8_0_3646), .B2(n_8_0_802), 
      .ZN(n_8_0_3275));
   OR2_X1 i_8_0_3377 (.A1(\out_as[6] [5]), .A2(n_8_0_802), .ZN(n_8_0_1371));
   AOI21_X1 i_8_0_3384 (.A(n_8_0_3674), .B1(n_8_0_3403), .B2(n_8_0_5116), 
      .ZN(n_8_0_3281));
   AOI211_X1 i_8_0_3386 (.A(n_8_0_3288), .B(n_8_0_3285), .C1(n_8_0_3284), 
      .C2(n_8_0_6082), .ZN(n_8_0_3283));
   OAI21_X1 i_8_0_3387 (.A(n_8_0_6811), .B1(n_8_0_3643), .B2(n_8_0_798), 
      .ZN(n_8_0_3284));
   OAI21_X1 i_8_0_3389 (.A(n_8_0_6754), .B1(n_8_0_6087), .B2(n_8_0_4562), 
      .ZN(n_8_0_3286));
   OAI21_X1 i_8_0_3390 (.A(n_8_0_3647), .B1(n_8_0_4560), .B2(n_8_0_6087), 
      .ZN(n_8_0_3287));
   OR2_X1 i_8_0_3391 (.A1(\out_as[6] [5]), .A2(n_8_0_786), .ZN(n_8_0_1372));
   NAND4_X1 i_8_0_3392 (.A1(n_8_0_4132), .A2(n_8_0_3293), .A3(n_8_0_3290), 
      .A4(n_8_0_3289), .ZN(n_8_0_3288));
   OR3_X1 i_8_0_3393 (.A1(n_8_0_798), .A2(n_8_0_3697), .A3(n_8_0_3643), .ZN(
      n_8_0_3289));
   NOR2_X1 i_8_0_3394 (.A1(n_8_0_3292), .A2(n_8_0_3291), .ZN(n_8_0_3290));
   AOI211_X1 i_8_0_3395 (.A(n_8_0_796), .B(n_8_0_3653), .C1(n_8_0_4199), 
      .C2(n_8_0_6075), .ZN(n_8_0_3291));
   OR2_X1 i_8_0_3396 (.A1(\out_as[1] [5]), .A2(n_8_0_796), .ZN(n_8_0_1373));
   AOI21_X1 i_8_0_3397 (.A(n_8_0_6782), .B1(n_8_0_6075), .B2(n_8_0_4325), 
      .ZN(n_8_0_3292));
   OAI21_X1 i_8_0_3398 (.A(n_8_0_3295), .B1(n_8_0_3294), .B2(n_8_0_6069), 
      .ZN(n_8_0_3293));
   OAI21_X1 i_8_0_3399 (.A(n_8_0_4367), .B1(n_8_0_3638), .B2(n_8_0_794), 
      .ZN(n_8_0_3294));
   OAI21_X1 i_8_0_3400 (.A(n_8_0_6772), .B1(n_8_0_3640), .B2(n_8_0_794), 
      .ZN(n_8_0_3295));
   OR2_X1 i_8_0_3401 (.A1(\out_as[2] [5]), .A2(n_8_0_794), .ZN(n_8_0_1374));
   AOI21_X1 i_8_0_3403 (.A(n_8_0_3620), .B1(n_8_0_3619), .B2(n_8_0_6097), 
      .ZN(n_8_0_3297));
   OAI21_X1 i_8_0_3405 (.A(n_8_0_4058), .B1(n_8_0_3300), .B2(n_8_0_790), 
      .ZN(n_8_0_3299));
   AOI21_X1 i_8_0_3406 (.A(n_8_0_3559), .B1(n_8_0_3406), .B2(n_8_0_6092), 
      .ZN(n_8_0_3300));
   AOI21_X1 i_8_0_3407 (.A(n_8_0_6853), .B1(n_8_0_3319), .B2(n_8_0_3301), 
      .ZN(n_121));
   NOR2_X1 i_8_0_3408 (.A1(n_8_0_3305), .A2(n_8_0_3302), .ZN(n_8_0_3301));
   OAI21_X1 i_8_0_3411 (.A(n_8_0_6471), .B1(n_8_0_3477), .B2(n_8_0_768), 
      .ZN(n_8_0_3304));
   NAND3_X1 i_8_0_3412 (.A1(n_8_0_3313), .A2(n_8_0_3310), .A3(n_8_0_3306), 
      .ZN(n_8_0_3305));
   NAND3_X1 i_8_0_3413 (.A1(n_8_0_3663), .A2(n_8_0_3308), .A3(n_8_0_3307), 
      .ZN(n_8_0_3306));
   OAI221_X1 i_8_0_3414 (.A(n_8_0_4110), .B1(n_8_0_6135), .B2(n_8_0_7022), 
      .C1(n_8_0_3662), .C2(n_8_0_772), .ZN(n_8_0_3307));
   NAND2_X1 i_8_0_3415 (.A1(n_8_0_6824), .A2(n_8_0_772), .ZN(n_8_0_3308));
   NOR2_X1 i_8_0_3417 (.A1(n_8_0_3312), .A2(n_8_0_3311), .ZN(n_8_0_3310));
   AOI21_X1 i_8_0_3418 (.A(n_8_0_6755), .B1(n_8_0_6123), .B2(n_8_0_4563), 
      .ZN(n_8_0_3311));
   AOI211_X1 i_8_0_3419 (.A(n_8_0_770), .B(n_8_0_3646), .C1(n_8_0_4561), 
      .C2(n_8_0_6123), .ZN(n_8_0_3312));
   OR2_X1 i_8_0_3420 (.A1(\out_as[6] [5]), .A2(n_8_0_770), .ZN(n_8_0_1375));
   AOI211_X1 i_8_0_3421 (.A(n_8_0_4133), .B(n_8_0_3316), .C1(n_8_0_3315), 
      .C2(n_8_0_3314), .ZN(n_8_0_3313));
   NAND2_X1 i_8_0_3422 (.A1(n_8_0_6139), .A2(n_8_0_3697), .ZN(n_8_0_3314));
   OAI22_X1 i_8_0_3423 (.A1(n_8_0_6811), .A2(n_8_0_6139), .B1(n_8_0_3643), 
      .B2(n_8_0_782), .ZN(n_8_0_3315));
   OAI21_X1 i_8_0_3424 (.A(n_8_0_3317), .B1(n_8_0_3318), .B2(n_8_0_780), 
      .ZN(n_8_0_3316));
   OAI21_X1 i_8_0_3425 (.A(n_8_0_6781), .B1(n_8_0_6127), .B2(n_8_0_4324), 
      .ZN(n_8_0_3317));
   OAI21_X1 i_8_0_3426 (.A(n_8_0_3654), .B1(n_8_0_4198), .B2(n_8_0_6127), 
      .ZN(n_8_0_3318));
   OR2_X1 i_8_0_3427 (.A1(\out_as[1] [5]), .A2(n_8_0_780), .ZN(n_8_0_1376));
   OR2_X1 i_8_0_3428 (.A1(\out_as[0] [5]), .A2(n_8_0_782), .ZN(n_8_0_1377));
   NOR3_X1 i_8_0_3429 (.A1(n_8_0_3326), .A2(n_8_0_3322), .A3(n_8_0_3320), 
      .ZN(n_8_0_3319));
   OAI221_X1 i_8_0_3430 (.A(n_8_0_3683), .B1(n_8_0_3321), .B2(n_8_0_776), 
      .C1(n_8_0_4309), .C2(n_8_0_6109), .ZN(n_8_0_3320));
   AOI21_X1 i_8_0_3431 (.A(n_8_0_3674), .B1(n_8_0_3403), .B2(n_8_0_6108), 
      .ZN(n_8_0_3321));
   NAND3_X1 i_8_0_3432 (.A1(n_8_0_4364), .A2(n_8_0_3324), .A3(n_8_0_3323), 
      .ZN(n_8_0_3322));
   NAND2_X1 i_8_0_3433 (.A1(n_8_0_6773), .A2(n_8_0_6131), .ZN(n_8_0_3323));
   OAI21_X1 i_8_0_3434 (.A(n_8_0_3325), .B1(n_8_0_4126), .B2(n_8_0_6131), 
      .ZN(n_8_0_3324));
   NOR2_X1 i_8_0_3435 (.A1(n_8_0_3640), .A2(n_8_0_778), .ZN(n_8_0_3325));
   OAI221_X1 i_8_0_3436 (.A(n_8_0_4058), .B1(n_8_0_3327), .B2(n_8_0_774), 
      .C1(n_8_0_6622), .C2(n_8_0_6114), .ZN(n_8_0_3326));
   AOI21_X1 i_8_0_3437 (.A(n_8_0_3559), .B1(n_8_0_3406), .B2(n_8_0_6113), 
      .ZN(n_8_0_3327));
   NAND2_X1 i_8_0_3440 (.A1(n_8_0_3343), .A2(n_8_0_3333), .ZN(n_8_0_3329));
   NAND3_X1 i_8_0_3442 (.A1(n_8_0_3347), .A2(n_8_0_3340), .A3(n_8_0_3332), 
      .ZN(n_8_0_3331));
   NOR2_X1 i_8_0_3443 (.A1(n_8_0_3345), .A2(n_8_0_3339), .ZN(n_8_0_3332));
   AOI21_X1 i_8_0_3444 (.A(n_8_0_3334), .B1(n_8_0_4310), .B2(n_8_0_6160), 
      .ZN(n_8_0_3333));
   OAI21_X1 i_8_0_3445 (.A(n_8_0_3683), .B1(n_8_0_3335), .B2(n_8_0_760), 
      .ZN(n_8_0_3334));
   AOI21_X1 i_8_0_3446 (.A(n_8_0_3674), .B1(n_8_0_3403), .B2(n_8_0_6160), 
      .ZN(n_8_0_3335));
   OAI21_X1 i_8_0_3449 (.A(n_8_0_6471), .B1(n_8_0_3477), .B2(n_8_0_752), 
      .ZN(n_8_0_3338));
   AOI21_X1 i_8_0_3450 (.A(n_8_0_6811), .B1(n_8_0_6174), .B2(n_8_0_4604), 
      .ZN(n_8_0_3339));
   NAND3_X1 i_8_0_3451 (.A1(n_8_0_3651), .A2(n_8_0_3342), .A3(n_8_0_3341), 
      .ZN(n_8_0_3340));
   OAI211_X1 i_8_0_3452 (.A(n_8_0_6147), .B(n_8_0_4325), .C1(n_8_0_3586), 
      .C2(n_8_0_764), .ZN(n_8_0_3341));
   NAND2_X1 i_8_0_3453 (.A1(n_8_0_764), .A2(n_8_0_6782), .ZN(n_8_0_3342));
   AOI211_X1 i_8_0_3454 (.A(n_8_0_4365), .B(n_8_0_3344), .C1(n_8_0_6773), 
      .C2(n_8_0_6150), .ZN(n_8_0_3343));
   AOI211_X1 i_8_0_3455 (.A(n_8_0_762), .B(n_8_0_3640), .C1(n_8_0_4127), 
      .C2(n_8_0_6151), .ZN(n_8_0_3344));
   AOI211_X1 i_8_0_3456 (.A(n_8_0_766), .B(n_8_0_3643), .C1(n_8_0_3697), 
      .C2(n_8_0_6174), .ZN(n_8_0_3345));
   OR2_X1 i_8_0_3457 (.A1(\out_as[0] [5]), .A2(n_8_0_766), .ZN(n_8_0_1378));
   INV_X1 i_8_0_3458 (.A(n_8_0_3347), .ZN(n_8_0_3346));
   NOR2_X1 i_8_0_3459 (.A1(n_8_0_3349), .A2(n_8_0_3348), .ZN(n_8_0_3347));
   AOI211_X1 i_8_0_3460 (.A(n_8_0_754), .B(n_8_0_3646), .C1(n_8_0_4561), 
      .C2(n_8_0_6293), .ZN(n_8_0_3348));
   OR2_X1 i_8_0_3461 (.A1(\out_as[6] [5]), .A2(n_8_0_754), .ZN(n_8_0_1379));
   AOI21_X1 i_8_0_3462 (.A(n_8_0_6755), .B1(n_8_0_6293), .B2(n_8_0_4563), 
      .ZN(n_8_0_3349));
   OAI221_X1 i_8_0_3463 (.A(n_8_0_3803), .B1(n_8_0_3623), .B2(n_8_0_6166), 
      .C1(n_8_0_3351), .C2(n_8_0_756), .ZN(n_8_0_3350));
   AOI21_X1 i_8_0_3464 (.A(n_8_0_3620), .B1(n_8_0_3619), .B2(n_8_0_6165), 
      .ZN(n_8_0_3351));
   AOI21_X1 i_8_0_3466 (.A(n_8_0_3559), .B1(n_8_0_3406), .B2(n_8_0_6170), 
      .ZN(n_8_0_3353));
   NAND4_X1 i_8_0_3470 (.A1(n_8_0_4132), .A2(n_8_0_3363), .A3(n_8_0_3360), 
      .A4(n_8_0_3369), .ZN(n_8_0_3356));
   OAI21_X1 i_8_0_3472 (.A(n_8_0_3359), .B1(n_8_0_3643), .B2(n_8_0_750), 
      .ZN(n_8_0_3358));
   NAND2_X1 i_8_0_3473 (.A1(n_8_0_6810), .A2(n_8_0_6185), .ZN(n_8_0_3359));
   AOI21_X1 i_8_0_3474 (.A(n_8_0_3361), .B1(n_8_0_3362), .B2(n_8_0_3651), 
      .ZN(n_8_0_3360));
   NOR2_X1 i_8_0_3475 (.A1(n_8_0_4197), .A2(n_8_0_1380), .ZN(n_8_0_3361));
   OR2_X1 i_8_0_3476 (.A1(\out_as[1] [5]), .A2(n_8_0_748), .ZN(n_8_0_1380));
   AOI22_X1 i_8_0_3477 (.A1(n_8_0_6206), .A2(n_8_0_4231), .B1(n_8_0_748), 
      .B2(n_8_0_6782), .ZN(n_8_0_3362));
   AOI211_X1 i_8_0_3478 (.A(n_8_0_4365), .B(n_8_0_3364), .C1(n_8_0_6773), 
      .C2(n_8_0_6181), .ZN(n_8_0_3363));
   AOI211_X1 i_8_0_3479 (.A(n_8_0_746), .B(n_8_0_3640), .C1(n_8_0_4127), 
      .C2(n_8_0_6182), .ZN(n_8_0_3364));
   AOI211_X1 i_8_0_3481 (.A(n_8_0_738), .B(n_8_0_3646), .C1(n_8_0_4561), 
      .C2(n_8_0_6196), .ZN(n_8_0_3366));
   OAI221_X1 i_8_0_3482 (.A(n_8_0_4058), .B1(n_8_0_6795), .B2(n_8_0_6190), 
      .C1(n_8_0_3368), .C2(n_8_0_742), .ZN(n_8_0_3367));
   AOI21_X1 i_8_0_3483 (.A(n_8_0_3559), .B1(n_8_0_3406), .B2(n_8_0_6191), 
      .ZN(n_8_0_3368));
   AOI21_X1 i_8_0_3484 (.A(n_8_0_3370), .B1(n_8_0_4310), .B2(n_8_0_6215), 
      .ZN(n_8_0_3369));
   OAI21_X1 i_8_0_3485 (.A(n_8_0_3683), .B1(n_8_0_3371), .B2(n_8_0_744), 
      .ZN(n_8_0_3370));
   AOI21_X1 i_8_0_3486 (.A(n_8_0_3674), .B1(n_8_0_3403), .B2(n_8_0_6215), 
      .ZN(n_8_0_3371));
   OAI21_X1 i_8_0_3488 (.A(n_8_0_3803), .B1(n_8_0_3374), .B2(n_8_0_740), 
      .ZN(n_8_0_3373));
   AOI21_X1 i_8_0_3489 (.A(n_8_0_3620), .B1(n_8_0_3619), .B2(n_8_0_6210), 
      .ZN(n_8_0_3374));
   AOI21_X1 i_8_0_3493 (.A(n_8_0_6853), .B1(n_8_0_3382), .B2(n_8_0_3378), 
      .ZN(n_122));
   NOR3_X1 i_8_0_3494 (.A1(n_8_0_3388), .A2(n_8_0_3379), .A3(n_8_0_3404), 
      .ZN(n_8_0_3378));
   NAND4_X1 i_8_0_3495 (.A1(n_8_0_3385), .A2(n_8_0_3383), .A3(n_8_0_3381), 
      .A4(n_8_0_3380), .ZN(n_8_0_3379));
   AOI21_X1 i_8_0_3496 (.A(n_8_0_4133), .B1(n_8_0_6233), .B2(n_8_0_3397), 
      .ZN(n_8_0_3380));
   NOR2_X1 i_8_0_3497 (.A1(n_8_0_3394), .A2(n_8_0_3398), .ZN(n_8_0_3381));
   NOR2_X1 i_8_0_3498 (.A1(n_8_0_3391), .A2(n_8_0_3400), .ZN(n_8_0_3382));
   OAI21_X1 i_8_0_3499 (.A(n_8_0_3384), .B1(n_8_0_3696), .B2(n_8_0_6253), 
      .ZN(n_8_0_3383));
   OAI22_X1 i_8_0_3500 (.A1(n_8_0_6811), .A2(n_8_0_6252), .B1(n_8_0_3643), 
      .B2(n_8_0_734), .ZN(n_8_0_3384));
   NOR2_X1 i_8_0_3501 (.A1(n_8_0_3387), .A2(n_8_0_3386), .ZN(n_8_0_3385));
   AOI21_X1 i_8_0_3502 (.A(n_8_0_6755), .B1(n_8_0_6226), .B2(n_8_0_4563), 
      .ZN(n_8_0_3386));
   AOI211_X1 i_8_0_3503 (.A(n_8_0_722), .B(n_8_0_3646), .C1(n_8_0_4561), 
      .C2(n_8_0_6226), .ZN(n_8_0_3387));
   OR2_X1 i_8_0_3504 (.A1(\out_as[6] [5]), .A2(n_8_0_722), .ZN(n_8_0_1381));
   AOI21_X1 i_8_0_3505 (.A(n_8_0_3389), .B1(n_8_0_6824), .B2(n_8_0_724), 
      .ZN(n_8_0_3388));
   NAND2_X1 i_8_0_3506 (.A1(n_8_0_3663), .A2(n_8_0_3390), .ZN(n_8_0_3389));
   OAI221_X1 i_8_0_3507 (.A(n_8_0_4110), .B1(n_8_0_6301), .B2(n_8_0_7022), 
      .C1(n_8_0_3662), .C2(n_8_0_724), .ZN(n_8_0_3390));
   AND2_X1 i_8_0_3508 (.A1(n_8_0_3393), .A2(n_8_0_3392), .ZN(n_8_0_3391));
   OAI211_X1 i_8_0_3509 (.A(n_8_0_6287), .B(n_8_0_4367), .C1(n_8_0_3638), 
      .C2(n_8_0_730), .ZN(n_8_0_3392));
   OAI21_X1 i_8_0_3510 (.A(n_8_0_6772), .B1(n_8_0_3640), .B2(n_8_0_730), 
      .ZN(n_8_0_3393));
   OR2_X1 i_8_0_3511 (.A1(\out_as[2] [5]), .A2(n_8_0_730), .ZN(n_8_0_1382));
   OAI211_X1 i_8_0_3512 (.A(n_8_0_4231), .B(n_8_0_3395), .C1(n_8_0_6782), 
      .C2(n_8_0_6270), .ZN(n_8_0_3394));
   OR3_X1 i_8_0_3513 (.A1(n_8_0_732), .A2(n_8_0_3396), .A3(n_8_0_3653), .ZN(
      n_8_0_3395));
   OR2_X1 i_8_0_3514 (.A1(\out_as[1] [5]), .A2(n_8_0_732), .ZN(n_8_0_1383));
   NOR3_X1 i_8_0_3515 (.A1(n_8_0_5394), .A2(n_8_0_6271), .A3(\out_bs[1] [5]), 
      .ZN(n_8_0_3396));
   OAI21_X1 i_8_0_3516 (.A(n_8_0_3399), .B1(n_8_0_3658), .B2(n_8_0_720), 
      .ZN(n_8_0_3397));
   NOR3_X1 i_8_0_3517 (.A1(n_8_0_720), .A2(n_8_0_3399), .A3(n_8_0_3658), 
      .ZN(n_8_0_3398));
   OR2_X1 i_8_0_3518 (.A1(\out_as[7] [5]), .A2(n_8_0_720), .ZN(n_8_0_1384));
   AOI21_X1 i_8_0_3519 (.A(n_8_0_4423), .B1(n_8_0_6237), .B2(\out_bs[7] [4]), 
      .ZN(n_8_0_3399));
   OAI221_X1 i_8_0_3520 (.A(n_8_0_3683), .B1(n_8_0_3401), .B2(n_8_0_728), 
      .C1(n_8_0_4309), .C2(n_8_0_6218), .ZN(n_8_0_3400));
   AOI21_X1 i_8_0_3521 (.A(n_8_0_3674), .B1(n_8_0_3403), .B2(n_8_0_6217), 
      .ZN(n_8_0_3401));
   NAND2_X1 i_8_0_3522 (.A1(\out_bs[3] [4]), .A2(n_8_0_3677), .ZN(n_8_0_3402));
   NOR2_X1 i_8_0_3523 (.A1(n_8_0_7045), .A2(n_8_0_3676), .ZN(n_8_0_3403));
   OAI221_X1 i_8_0_3524 (.A(n_8_0_4058), .B1(n_8_0_3405), .B2(n_8_0_726), 
      .C1(n_8_0_6622), .C2(n_8_0_6245), .ZN(n_8_0_3404));
   AOI21_X1 i_8_0_3525 (.A(n_8_0_3559), .B1(n_8_0_3406), .B2(n_8_0_6244), 
      .ZN(n_8_0_3405));
   NOR2_X1 i_8_0_3526 (.A1(n_8_0_7033), .A2(n_8_0_3669), .ZN(n_8_0_3406));
   NOR2_X1 i_8_0_3527 (.A1(n_8_0_3407), .A2(n_8_0_6853), .ZN(n_123));
   NOR3_X1 i_8_0_3528 (.A1(n_8_0_3424), .A2(n_8_0_3409), .A3(n_8_0_3408), 
      .ZN(n_8_0_3407));
   NAND3_X1 i_8_0_3529 (.A1(n_8_0_3421), .A2(n_8_0_3418), .A3(n_8_0_3412), 
      .ZN(n_8_0_3408));
   OAI211_X1 i_8_0_3530 (.A(n_8_0_4422), .B(n_8_0_3410), .C1(n_8_0_3478), 
      .C2(n_8_0_704), .ZN(n_8_0_3409));
   NAND2_X1 i_8_0_3531 (.A1(n_8_0_6278), .A2(n_8_0_3411), .ZN(n_8_0_3410));
   OAI21_X1 i_8_0_3532 (.A(n_8_0_6471), .B1(n_8_0_3477), .B2(n_8_0_704), 
      .ZN(n_8_0_3411));
   NOR3_X1 i_8_0_3533 (.A1(n_8_0_3417), .A2(n_8_0_3416), .A3(n_8_0_3413), 
      .ZN(n_8_0_3412));
   AOI21_X1 i_8_0_3534 (.A(n_8_0_3414), .B1(n_8_0_3415), .B2(n_8_0_716), 
      .ZN(n_8_0_3413));
   OAI21_X1 i_8_0_3535 (.A(n_8_0_3651), .B1(n_8_0_3585), .B2(n_8_0_6268), 
      .ZN(n_8_0_3414));
   OAI21_X1 i_8_0_3536 (.A(n_8_0_6781), .B1(n_8_0_6268), .B2(n_8_0_4324), 
      .ZN(n_8_0_3415));
   AOI21_X1 i_8_0_3537 (.A(n_8_0_6811), .B1(n_8_0_6261), .B2(n_8_0_4604), 
      .ZN(n_8_0_3416));
   AOI211_X1 i_8_0_3538 (.A(n_8_0_718), .B(n_8_0_3643), .C1(n_8_0_3697), 
      .C2(n_8_0_6261), .ZN(n_8_0_3417));
   NOR2_X1 i_8_0_3539 (.A1(n_8_0_4346), .A2(n_8_0_3419), .ZN(n_8_0_3418));
   OAI22_X1 i_8_0_3540 (.A1(n_8_0_6755), .A2(n_8_0_6292), .B1(n_8_0_3420), 
      .B2(n_8_0_706), .ZN(n_8_0_3419));
   OAI211_X1 i_8_0_3541 (.A(n_8_0_7018), .B(n_8_0_7017), .C1(n_8_0_6291), 
      .C2(n_8_0_4560), .ZN(n_8_0_3420));
   AOI21_X1 i_8_0_3542 (.A(n_8_0_3422), .B1(n_8_0_3622), .B2(n_8_0_6299), 
      .ZN(n_8_0_3421));
   OAI21_X1 i_8_0_3543 (.A(n_8_0_3803), .B1(n_8_0_3423), .B2(n_8_0_708), 
      .ZN(n_8_0_3422));
   AOI21_X1 i_8_0_3544 (.A(n_8_0_3620), .B1(n_8_0_3619), .B2(n_8_0_6299), 
      .ZN(n_8_0_3423));
   NAND3_X1 i_8_0_3545 (.A1(n_8_0_3431), .A2(n_8_0_3428), .A3(n_8_0_3425), 
      .ZN(n_8_0_3424));
   OAI21_X1 i_8_0_3546 (.A(n_8_0_3427), .B1(n_8_0_3426), .B2(n_8_0_6285), 
      .ZN(n_8_0_3425));
   OAI21_X1 i_8_0_3547 (.A(n_8_0_4367), .B1(n_8_0_3638), .B2(n_8_0_714), 
      .ZN(n_8_0_3426));
   OAI21_X1 i_8_0_3548 (.A(n_8_0_6772), .B1(n_8_0_3640), .B2(n_8_0_714), 
      .ZN(n_8_0_3427));
   OR2_X1 i_8_0_3549 (.A1(\out_as[2] [5]), .A2(n_8_0_714), .ZN(n_8_0_1385));
   AOI211_X1 i_8_0_3550 (.A(n_8_0_4059), .B(n_8_0_3429), .C1(n_8_0_6794), 
      .C2(n_8_0_6275), .ZN(n_8_0_3428));
   NOR3_X1 i_8_0_3551 (.A1(n_8_0_710), .A2(n_8_0_3430), .A3(n_8_0_3669), 
      .ZN(n_8_0_3429));
   OR2_X1 i_8_0_3552 (.A1(\out_as[4] [5]), .A2(n_8_0_710), .ZN(n_8_0_1386));
   NOR3_X1 i_8_0_3553 (.A1(n_8_0_5459), .A2(\out_bs[4] [5]), .A3(n_8_0_6275), 
      .ZN(n_8_0_3430));
   AOI211_X1 i_8_0_3554 (.A(n_8_0_3432), .B(n_8_0_3449), .C1(n_8_0_4310), 
      .C2(n_8_0_6650), .ZN(n_8_0_3431));
   AOI211_X1 i_8_0_3555 (.A(n_8_0_712), .B(n_8_0_3676), .C1(n_8_0_3452), 
      .C2(n_8_0_4311), .ZN(n_8_0_3432));
   OR2_X1 i_8_0_3556 (.A1(\out_as[3] [5]), .A2(n_8_0_712), .ZN(n_8_0_1387));
   NOR2_X1 i_8_0_3557 (.A1(n_8_0_3433), .A2(n_8_0_6853), .ZN(n_124));
   NOR3_X1 i_8_0_3558 (.A1(n_8_0_3436), .A2(n_8_0_3434), .A3(n_8_0_3457), 
      .ZN(n_8_0_3433));
   NAND4_X1 i_8_0_3559 (.A1(n_8_0_3437), .A2(n_8_0_3435), .A3(n_8_0_3442), 
      .A4(n_8_0_3439), .ZN(n_8_0_3434));
   OAI21_X1 i_8_0_3560 (.A(n_8_0_6810), .B1(n_8_0_6663), .B2(n_8_0_4603), 
      .ZN(n_8_0_3435));
   NAND4_X1 i_8_0_3561 (.A1(n_8_0_3455), .A2(n_8_0_3453), .A3(n_8_0_3447), 
      .A4(n_8_0_3445), .ZN(n_8_0_3436));
   AOI211_X1 i_8_0_3562 (.A(n_8_0_4232), .B(n_8_0_3438), .C1(n_8_0_6781), 
      .C2(n_8_0_6696), .ZN(n_8_0_3437));
   AOI211_X1 i_8_0_3563 (.A(n_8_0_699), .B(n_8_0_3653), .C1(n_8_0_4199), 
      .C2(n_8_0_6695), .ZN(n_8_0_3438));
   OR2_X1 i_8_0_3564 (.A1(\out_as[1] [5]), .A2(n_8_0_699), .ZN(n_8_0_1388));
   NAND2_X1 i_8_0_3565 (.A1(n_8_0_3441), .A2(n_8_0_3440), .ZN(n_8_0_3439));
   OAI21_X1 i_8_0_3566 (.A(n_8_0_6730), .B1(n_8_0_3658), .B2(n_8_0_681), 
      .ZN(n_8_0_3440));
   OAI211_X1 i_8_0_3567 (.A(n_8_0_6721), .B(n_8_0_4424), .C1(n_8_0_3657), 
      .C2(n_8_0_681), .ZN(n_8_0_3441));
   OR2_X1 i_8_0_3568 (.A1(\out_as[7] [5]), .A2(n_8_0_681), .ZN(n_8_0_1389));
   OAI21_X1 i_8_0_3569 (.A(n_8_0_3444), .B1(n_8_0_3443), .B2(n_8_0_6709), 
      .ZN(n_8_0_3442));
   OAI21_X1 i_8_0_3570 (.A(n_8_0_4367), .B1(n_8_0_3638), .B2(n_8_0_696), 
      .ZN(n_8_0_3443));
   OAI21_X1 i_8_0_3571 (.A(n_8_0_6772), .B1(n_8_0_3640), .B2(n_8_0_696), 
      .ZN(n_8_0_3444));
   OR2_X1 i_8_0_3572 (.A1(\out_as[2] [5]), .A2(n_8_0_696), .ZN(n_8_0_1390));
   INV_X1 i_8_0_3573 (.A(n_8_0_3446), .ZN(n_8_0_3445));
   AOI211_X1 i_8_0_3574 (.A(n_8_0_702), .B(n_8_0_3643), .C1(n_8_0_3697), 
      .C2(n_8_0_6662), .ZN(n_8_0_3446));
   NOR2_X1 i_8_0_3575 (.A1(n_8_0_3449), .A2(n_8_0_3450), .ZN(n_8_0_3447));
   INV_X1 i_8_0_3576 (.A(n_8_0_3449), .ZN(n_8_0_3448));
   OAI21_X1 i_8_0_3577 (.A(n_8_0_3683), .B1(n_8_0_6647), .B2(n_8_0_6837), 
      .ZN(n_8_0_3449));
   NOR2_X1 i_8_0_3578 (.A1(n_8_0_693), .A2(n_8_0_3451), .ZN(n_8_0_3450));
   OAI21_X1 i_8_0_3579 (.A(n_8_0_3677), .B1(n_8_0_3675), .B2(n_8_0_6648), 
      .ZN(n_8_0_3451));
   NOR2_X1 i_8_0_3580 (.A1(n_8_0_3675), .A2(\out_as[3] [6]), .ZN(n_8_0_3452));
   AOI211_X1 i_8_0_3581 (.A(n_8_0_4059), .B(n_8_0_3454), .C1(n_8_0_6794), 
      .C2(n_8_0_6633), .ZN(n_8_0_3453));
   AOI211_X1 i_8_0_3582 (.A(n_8_0_690), .B(n_8_0_3669), .C1(n_8_0_4385), 
      .C2(n_8_0_6632), .ZN(n_8_0_3454));
   NOR2_X1 i_8_0_3583 (.A1(n_8_0_3456), .A2(n_8_0_3804), .ZN(n_8_0_3455));
   OAI21_X1 i_8_0_3584 (.A(n_8_0_3621), .B1(n_8_0_3617), .B2(n_8_0_687), 
      .ZN(n_8_0_3456));
   OAI21_X1 i_8_0_3585 (.A(n_8_0_3459), .B1(n_8_0_3458), .B2(n_8_0_684), 
      .ZN(n_8_0_3457));
   OAI21_X1 i_8_0_3586 (.A(n_8_0_3647), .B1(n_8_0_4560), .B2(n_8_0_6751), 
      .ZN(n_8_0_3458));
   OR2_X1 i_8_0_3587 (.A1(\out_as[6] [5]), .A2(n_8_0_684), .ZN(n_8_0_1391));
   OAI21_X1 i_8_0_3588 (.A(n_8_0_6754), .B1(n_8_0_6751), .B2(n_8_0_4562), 
      .ZN(n_8_0_3459));
   AOI211_X1 i_8_0_3592 (.A(n_8_0_3471), .B(n_8_0_3463), .C1(n_8_0_6810), 
      .C2(n_8_0_6343), .ZN(n_8_0_3462));
   OAI21_X1 i_8_0_3593 (.A(n_8_0_3464), .B1(n_8_0_3465), .B2(n_8_0_669), 
      .ZN(n_8_0_3463));
   OAI21_X1 i_8_0_3594 (.A(n_8_0_6838), .B1(n_8_0_6356), .B2(n_8_0_3685), 
      .ZN(n_8_0_3464));
   OAI21_X1 i_8_0_3595 (.A(n_8_0_3677), .B1(n_8_0_3675), .B2(n_8_0_6356), 
      .ZN(n_8_0_3465));
   OAI21_X1 i_8_0_3596 (.A(n_8_0_3467), .B1(n_8_0_3696), .B2(n_8_0_6343), 
      .ZN(n_8_0_3466));
   OAI21_X1 i_8_0_3597 (.A(n_8_0_4132), .B1(n_8_0_3643), .B2(n_8_0_678), 
      .ZN(n_8_0_3467));
   OAI21_X1 i_8_0_3599 (.A(n_8_0_3470), .B1(n_8_0_4126), .B2(n_8_0_6334), 
      .ZN(n_8_0_3469));
   NOR2_X1 i_8_0_3600 (.A1(n_8_0_3640), .A2(n_8_0_672), .ZN(n_8_0_3470));
   OAI211_X1 i_8_0_3601 (.A(n_8_0_4231), .B(n_8_0_3472), .C1(n_8_0_6782), 
      .C2(n_8_0_6339), .ZN(n_8_0_3471));
   OAI21_X1 i_8_0_3602 (.A(n_8_0_3473), .B1(n_8_0_4198), .B2(n_8_0_6340), 
      .ZN(n_8_0_3472));
   NOR2_X1 i_8_0_3603 (.A1(n_8_0_3653), .A2(n_8_0_675), .ZN(n_8_0_3473));
   AOI211_X1 i_8_0_3609 (.A(n_8_0_4059), .B(n_8_0_3480), .C1(n_8_0_6623), 
      .C2(n_8_0_6351), .ZN(n_8_0_3479));
   AOI211_X1 i_8_0_3610 (.A(n_8_0_666), .B(n_8_0_3669), .C1(n_8_0_4385), 
      .C2(n_8_0_6348), .ZN(n_8_0_3480));
   OAI21_X1 i_8_0_3611 (.A(n_8_0_3483), .B1(n_8_0_3482), .B2(n_8_0_6373), 
      .ZN(n_8_0_3481));
   OAI21_X1 i_8_0_3612 (.A(n_8_0_4110), .B1(n_8_0_1392), .B2(n_8_0_4573), 
      .ZN(n_8_0_3482));
   OAI21_X1 i_8_0_3613 (.A(n_8_0_6824), .B1(n_8_0_3664), .B2(n_8_0_663), 
      .ZN(n_8_0_3483));
   OR2_X1 i_8_0_3614 (.A1(\out_as[5] [5]), .A2(n_8_0_663), .ZN(n_8_0_1392));
   OAI21_X1 i_8_0_3616 (.A(n_8_0_3647), .B1(n_8_0_4560), .B2(n_8_0_6367), 
      .ZN(n_8_0_3485));
   OR2_X1 i_8_0_3617 (.A1(\out_as[6] [5]), .A2(n_8_0_660), .ZN(n_8_0_1393));
   OAI21_X1 i_8_0_3618 (.A(n_8_0_6754), .B1(n_8_0_6367), .B2(n_8_0_4562), 
      .ZN(n_8_0_3486));
   AOI21_X1 i_8_0_3619 (.A(n_8_0_6853), .B1(n_8_0_3509), .B2(n_8_0_3487), 
      .ZN(n_125));
   NOR2_X1 i_8_0_3620 (.A1(n_8_0_3506), .A2(n_8_0_3488), .ZN(n_8_0_3487));
   NAND4_X1 i_8_0_3621 (.A1(n_8_0_3491), .A2(n_8_0_3489), .A3(n_8_0_3503), 
      .A4(n_8_0_3494), .ZN(n_8_0_3488));
   NAND3_X1 i_8_0_3622 (.A1(n_8_0_3490), .A2(n_8_0_6663), .A3(n_8_0_6420), 
      .ZN(n_8_0_3489));
   OAI21_X1 i_8_0_3623 (.A(n_8_0_6811), .B1(n_8_0_3643), .B2(n_8_0_654), 
      .ZN(n_8_0_3490));
   OAI21_X1 i_8_0_3624 (.A(n_8_0_3492), .B1(n_8_0_4126), .B2(n_8_0_6398), 
      .ZN(n_8_0_3491));
   OAI21_X1 i_8_0_3625 (.A(n_8_0_3493), .B1(n_8_0_3640), .B2(n_8_0_648), 
      .ZN(n_8_0_3492));
   OAI21_X1 i_8_0_3626 (.A(n_8_0_6773), .B1(n_8_0_6398), .B2(n_8_0_4366), 
      .ZN(n_8_0_3493));
   NOR2_X1 i_8_0_3627 (.A1(n_8_0_3500), .A2(n_8_0_3495), .ZN(n_8_0_3494));
   AOI21_X1 i_8_0_3628 (.A(n_8_0_3496), .B1(n_8_0_3497), .B2(n_8_0_6232), 
      .ZN(n_8_0_3495));
   NOR2_X1 i_8_0_3629 (.A1(n_8_0_3499), .A2(n_8_0_3498), .ZN(n_8_0_3496));
   NAND2_X1 i_8_0_3630 (.A1(n_8_0_3499), .A2(n_8_0_3498), .ZN(n_8_0_3497));
   OAI21_X1 i_8_0_3631 (.A(n_8_0_4424), .B1(n_8_0_6405), .B2(n_8_0_6721), 
      .ZN(n_8_0_3498));
   NOR2_X1 i_8_0_3632 (.A1(n_8_0_3658), .A2(n_8_0_633), .ZN(n_8_0_3499));
   OR2_X1 i_8_0_3633 (.A1(\out_as[7] [5]), .A2(n_8_0_633), .ZN(n_8_0_1394));
   OAI211_X1 i_8_0_3634 (.A(n_8_0_4231), .B(n_8_0_3501), .C1(n_8_0_6782), 
      .C2(n_8_0_6392), .ZN(n_8_0_3500));
   INV_X1 i_8_0_3635 (.A(n_8_0_3502), .ZN(n_8_0_3501));
   AOI211_X1 i_8_0_3636 (.A(n_8_0_651), .B(n_8_0_3653), .C1(n_8_0_4199), 
      .C2(n_8_0_6392), .ZN(n_8_0_3502));
   OAI21_X1 i_8_0_3637 (.A(n_8_0_3504), .B1(n_8_0_4384), .B2(n_8_0_6380), 
      .ZN(n_8_0_3503));
   OAI21_X1 i_8_0_3638 (.A(n_8_0_3505), .B1(n_8_0_3669), .B2(n_8_0_642), 
      .ZN(n_8_0_3504));
   OR2_X1 i_8_0_3639 (.A1(\out_as[4] [5]), .A2(n_8_0_642), .ZN(n_8_0_1395));
   OAI21_X1 i_8_0_3640 (.A(n_8_0_6794), .B1(n_8_0_6380), .B2(n_8_0_4486), 
      .ZN(n_8_0_3505));
   OAI211_X1 i_8_0_3641 (.A(n_8_0_3803), .B(n_8_0_3508), .C1(n_8_0_3507), 
      .C2(n_8_0_639), .ZN(n_8_0_3506));
   AOI21_X1 i_8_0_3642 (.A(n_8_0_3620), .B1(n_8_0_3619), .B2(n_8_0_6409), 
      .ZN(n_8_0_3507));
   NAND2_X1 i_8_0_3643 (.A1(n_8_0_6409), .A2(n_8_0_3622), .ZN(n_8_0_3508));
   AOI211_X1 i_8_0_3644 (.A(n_8_0_3514), .B(n_8_0_3511), .C1(n_8_0_3510), 
      .C2(n_8_0_3696), .ZN(n_8_0_3509));
   OAI21_X1 i_8_0_3645 (.A(n_8_0_4132), .B1(n_8_0_3643), .B2(n_8_0_654), 
      .ZN(n_8_0_3510));
   OR2_X1 i_8_0_3646 (.A1(\out_as[0] [5]), .A2(n_8_0_654), .ZN(n_8_0_1396));
   OAI21_X1 i_8_0_3647 (.A(n_8_0_3513), .B1(n_8_0_3512), .B2(n_8_0_636), 
      .ZN(n_8_0_3511));
   OAI21_X1 i_8_0_3648 (.A(n_8_0_3647), .B1(n_8_0_4560), .B2(n_8_0_6385), 
      .ZN(n_8_0_3512));
   OR2_X1 i_8_0_3649 (.A1(\out_as[6] [5]), .A2(n_8_0_636), .ZN(n_8_0_1397));
   OAI21_X1 i_8_0_3650 (.A(n_8_0_6754), .B1(n_8_0_6385), .B2(n_8_0_4562), 
      .ZN(n_8_0_3513));
   AND2_X1 i_8_0_3651 (.A1(n_8_0_3516), .A2(n_8_0_3515), .ZN(n_8_0_3514));
   OAI21_X1 i_8_0_3652 (.A(n_8_0_6837), .B1(n_8_0_3676), .B2(n_8_0_645), 
      .ZN(n_8_0_3515));
   OAI221_X1 i_8_0_3653 (.A(n_8_0_3686), .B1(n_8_0_6414), .B2(n_8_0_6647), 
      .C1(n_8_0_3673), .C2(n_8_0_645), .ZN(n_8_0_3516));
   AOI21_X1 i_8_0_3654 (.A(n_8_0_6853), .B1(n_8_0_3524), .B2(n_8_0_3517), 
      .ZN(n_126));
   NOR2_X1 i_8_0_3655 (.A1(n_8_0_3534), .A2(n_8_0_3518), .ZN(n_8_0_3517));
   NAND4_X1 i_8_0_3656 (.A1(n_8_0_3536), .A2(n_8_0_3530), .A3(n_8_0_3527), 
      .A4(n_8_0_3519), .ZN(n_8_0_3518));
   NOR4_X1 i_8_0_3657 (.A1(n_8_0_3541), .A2(n_8_0_3539), .A3(n_8_0_3520), 
      .A4(n_8_0_4133), .ZN(n_8_0_3519));
   NAND2_X1 i_8_0_3658 (.A1(n_8_0_3523), .A2(n_8_0_3521), .ZN(n_8_0_3520));
   OAI21_X1 i_8_0_3659 (.A(n_8_0_3522), .B1(n_8_0_4198), .B2(n_8_0_6446), 
      .ZN(n_8_0_3521));
   NOR2_X1 i_8_0_3660 (.A1(n_8_0_3653), .A2(n_8_0_627), .ZN(n_8_0_3522));
   OR2_X1 i_8_0_3661 (.A1(\out_as[1] [5]), .A2(n_8_0_627), .ZN(n_8_0_1398));
   OAI21_X1 i_8_0_3662 (.A(n_8_0_6781), .B1(n_8_0_6446), .B2(n_8_0_4324), 
      .ZN(n_8_0_3523));
   NOR2_X1 i_8_0_3663 (.A1(n_8_0_3526), .A2(n_8_0_3525), .ZN(n_8_0_3524));
   AOI21_X1 i_8_0_3664 (.A(n_8_0_6772), .B1(n_8_0_5337), .B2(n_8_0_7060), 
      .ZN(n_8_0_3525));
   AOI211_X1 i_8_0_3665 (.A(n_8_0_3640), .B(n_8_0_624), .C1(n_8_0_5428), 
      .C2(n_8_0_5337), .ZN(n_8_0_3526));
   NOR2_X1 i_8_0_3666 (.A1(n_8_0_3529), .A2(n_8_0_3528), .ZN(n_8_0_3527));
   AOI21_X1 i_8_0_3667 (.A(n_8_0_6730), .B1(n_8_0_6473), .B2(n_8_0_4424), 
      .ZN(n_8_0_3528));
   AOI211_X1 i_8_0_3668 (.A(n_8_0_609), .B(n_8_0_3658), .C1(n_8_0_3692), 
      .C2(n_8_0_6473), .ZN(n_8_0_3529));
   OR2_X1 i_8_0_3669 (.A1(\out_as[7] [5]), .A2(n_8_0_609), .ZN(n_8_0_1399));
   OAI21_X1 i_8_0_3670 (.A(n_8_0_3531), .B1(n_8_0_3532), .B2(n_8_0_3533), 
      .ZN(n_8_0_3530));
   OAI21_X1 i_8_0_3671 (.A(n_8_0_6837), .B1(n_8_0_3676), .B2(n_8_0_621), 
      .ZN(n_8_0_3531));
   OAI21_X1 i_8_0_3672 (.A(n_8_0_3686), .B1(n_8_0_6429), .B2(n_8_0_6647), 
      .ZN(n_8_0_3532));
   NOR3_X1 i_8_0_3673 (.A1(n_8_0_621), .A2(n_8_0_6847), .A3(n_8_0_3676), 
      .ZN(n_8_0_3533));
   OR2_X1 i_8_0_3674 (.A1(\out_as[3] [5]), .A2(n_8_0_621), .ZN(n_8_0_1400));
   OAI221_X1 i_8_0_3675 (.A(n_8_0_3803), .B1(n_8_0_3623), .B2(n_8_0_6459), 
      .C1(n_8_0_3535), .C2(n_8_0_615), .ZN(n_8_0_3534));
   AOI21_X1 i_8_0_3676 (.A(n_8_0_3620), .B1(n_8_0_3619), .B2(n_8_0_6460), 
      .ZN(n_8_0_3535));
   NOR2_X1 i_8_0_3677 (.A1(n_8_0_3538), .A2(n_8_0_3537), .ZN(n_8_0_3536));
   AOI21_X1 i_8_0_3678 (.A(n_8_0_6795), .B1(n_8_0_6433), .B2(n_8_0_4487), 
      .ZN(n_8_0_3537));
   AOI211_X1 i_8_0_3679 (.A(n_8_0_618), .B(n_8_0_3669), .C1(n_8_0_4385), 
      .C2(n_8_0_6433), .ZN(n_8_0_3538));
   OR2_X1 i_8_0_3680 (.A1(\out_as[4] [5]), .A2(n_8_0_618), .ZN(n_8_0_1401));
   OAI33_X1 i_8_0_3681 (.A1(n_8_0_6811), .A2(n_8_0_6662), .A3(n_8_0_6442), 
      .B1(n_8_0_3540), .B2(n_8_0_3643), .B3(n_8_0_630), .ZN(n_8_0_3539));
   NOR2_X1 i_8_0_3682 (.A1(n_8_0_3696), .A2(n_8_0_6439), .ZN(n_8_0_3540));
   OAI21_X1 i_8_0_3683 (.A(n_8_0_3542), .B1(n_8_0_3543), .B2(n_8_0_612), 
      .ZN(n_8_0_3541));
   OAI21_X1 i_8_0_3684 (.A(n_8_0_6754), .B1(n_8_0_6479), .B2(n_8_0_4562), 
      .ZN(n_8_0_3542));
   OAI21_X1 i_8_0_3685 (.A(n_8_0_3647), .B1(n_8_0_4560), .B2(n_8_0_6479), 
      .ZN(n_8_0_3543));
   NOR3_X1 i_8_0_3690 (.A1(n_8_0_606), .A2(n_8_0_3697), .A3(n_8_0_3643), 
      .ZN(n_8_0_3547));
   NOR2_X1 i_8_0_3692 (.A1(n_8_0_4197), .A2(n_8_0_1402), .ZN(n_8_0_3549));
   OR2_X1 i_8_0_3693 (.A1(\out_as[1] [5]), .A2(n_8_0_602), .ZN(n_8_0_1402));
   AOI211_X1 i_8_0_3694 (.A(n_8_0_6689), .B(n_8_0_3652), .C1(n_8_0_602), 
      .C2(n_8_0_6782), .ZN(n_8_0_3550));
   OAI21_X1 i_8_0_3695 (.A(n_8_0_3553), .B1(n_8_0_3552), .B2(n_8_0_582), 
      .ZN(n_8_0_3551));
   OAI21_X1 i_8_0_3696 (.A(n_8_0_3647), .B1(n_8_0_4560), .B2(n_8_0_6749), 
      .ZN(n_8_0_3552));
   OAI21_X1 i_8_0_3697 (.A(n_8_0_6754), .B1(n_8_0_6749), .B2(n_8_0_4562), 
      .ZN(n_8_0_3553));
   OR2_X1 i_8_0_3698 (.A1(\out_as[6] [5]), .A2(n_8_0_582), .ZN(n_8_0_1403));
   OR2_X1 i_8_0_3702 (.A1(\out_as[7] [5]), .A2(n_8_0_578), .ZN(n_8_0_1404));
   NOR2_X1 i_8_0_3705 (.A1(n_8_0_4385), .A2(n_8_0_3669), .ZN(n_8_0_3559));
   OR2_X1 i_8_0_3706 (.A1(\out_as[4] [5]), .A2(n_8_0_590), .ZN(n_8_0_1405));
   OAI21_X1 i_8_0_3707 (.A(n_8_0_6795), .B1(n_8_0_3669), .B2(n_8_0_590), 
      .ZN(n_8_0_3560));
   OAI21_X1 i_8_0_3709 (.A(n_8_0_3563), .B1(n_8_0_4126), .B2(n_8_0_6707), 
      .ZN(n_8_0_3562));
   OAI22_X1 i_8_0_3710 (.A1(n_8_0_6772), .A2(n_8_0_6706), .B1(n_8_0_3640), 
      .B2(n_8_0_598), .ZN(n_8_0_3563));
   AND3_X1 i_8_0_3711 (.A1(n_8_0_3565), .A2(n_8_0_6663), .A3(\out_bs[0] [2]), 
      .ZN(n_8_0_3564));
   OAI21_X1 i_8_0_3712 (.A(n_8_0_6811), .B1(n_8_0_3643), .B2(n_8_0_606), 
      .ZN(n_8_0_3565));
   OR2_X1 i_8_0_3713 (.A1(\out_as[0] [5]), .A2(n_8_0_606), .ZN(n_8_0_1406));
   OAI211_X1 i_8_0_3715 (.A(n_8_0_5467), .B(n_8_0_3686), .C1(n_8_0_3673), 
      .C2(n_8_0_594), .ZN(n_8_0_3567));
   OAI21_X1 i_8_0_3716 (.A(n_8_0_6837), .B1(n_8_0_3676), .B2(n_8_0_594), 
      .ZN(n_8_0_3568));
   OR2_X1 i_8_0_3717 (.A1(\out_as[3] [5]), .A2(n_8_0_594), .ZN(n_8_0_1407));
   NAND2_X1 i_8_0_3721 (.A1(n_8_0_6810), .A2(n_8_0_6520), .ZN(n_8_0_3571));
   OAI21_X1 i_8_0_3722 (.A(n_8_0_3590), .B1(n_8_0_3696), .B2(n_8_0_6520), 
      .ZN(n_8_0_3572));
   AOI211_X1 i_8_0_3725 (.A(n_8_0_550), .B(n_8_0_3646), .C1(n_8_0_4561), 
      .C2(n_8_0_6548), .ZN(n_8_0_3575));
   OR2_X1 i_8_0_3726 (.A1(\out_as[6] [5]), .A2(n_8_0_550), .ZN(n_8_0_1408));
   AOI21_X1 i_8_0_3727 (.A(n_8_0_6755), .B1(n_8_0_6548), .B2(n_8_0_4563), 
      .ZN(n_8_0_3576));
   AOI22_X1 i_8_0_3729 (.A1(n_8_0_6794), .A2(n_8_0_6558), .B1(n_8_0_3670), 
      .B2(n_8_0_3579), .ZN(n_8_0_3578));
   AOI21_X1 i_8_0_3730 (.A(n_8_0_558), .B1(n_8_0_5460), .B2(n_8_0_5409), 
      .ZN(n_8_0_3579));
   OR2_X1 i_8_0_3734 (.A1(\out_as[7] [5]), .A2(n_8_0_546), .ZN(n_8_0_1409));
   OAI211_X1 i_8_0_3735 (.A(n_8_0_3651), .B(n_8_0_3584), .C1(n_8_0_6860), 
      .C2(n_8_0_6781), .ZN(n_8_0_3583));
   OAI211_X1 i_8_0_3736 (.A(n_8_0_6530), .B(n_8_0_4325), .C1(n_8_0_3586), 
      .C2(n_8_0_570), .ZN(n_8_0_3584));
   NAND2_X1 i_8_0_3737 (.A1(n_8_0_3586), .A2(n_8_0_4325), .ZN(n_8_0_3585));
   NAND2_X1 i_8_0_3738 (.A1(n_8_0_6788), .A2(n_8_0_3654), .ZN(n_8_0_3586));
   NOR3_X1 i_8_0_3740 (.A1(n_8_0_566), .A2(n_8_0_5428), .A3(n_8_0_3640), 
      .ZN(n_8_0_3588));
   OAI21_X1 i_8_0_3741 (.A(n_8_0_6772), .B1(n_8_0_3640), .B2(n_8_0_566), 
      .ZN(n_8_0_3589));
   NOR2_X1 i_8_0_3742 (.A1(n_8_0_3643), .A2(n_8_0_574), .ZN(n_8_0_3590));
   OAI21_X1 i_8_0_3744 (.A(n_8_0_4494), .B1(n_8_0_3673), .B2(n_8_0_562), 
      .ZN(n_8_0_3592));
   OAI21_X1 i_8_0_3745 (.A(n_8_0_6837), .B1(n_8_0_3676), .B2(n_8_0_562), 
      .ZN(n_8_0_3593));
   OR2_X1 i_8_0_3746 (.A1(\out_as[3] [5]), .A2(n_8_0_562), .ZN(n_8_0_1410));
   AOI21_X1 i_8_0_3748 (.A(n_8_0_3620), .B1(n_8_0_3619), .B2(n_8_0_6516), 
      .ZN(n_8_0_3595));
   AOI21_X1 i_8_0_3749 (.A(n_8_0_3620), .B1(n_8_0_3618), .B2(\out_bs[5] [2]), 
      .ZN(n_8_0_3596));
   NAND3_X1 i_8_0_3750 (.A1(\out_bs[5] [3]), .A2(n_8_0_6517), .A3(n_8_0_3622), 
      .ZN(n_8_0_3597));
   NAND3_X1 i_8_0_3751 (.A1(\out_bs[5] [4]), .A2(n_8_0_6825), .A3(n_8_0_6679), 
      .ZN(n_8_0_3598));
   OR2_X1 i_8_0_3758 (.A1(\out_as[7] [5]), .A2(n_8_0_507), .ZN(n_8_0_1411));
   INV_X1 i_8_0_3761 (.A(n_8_0_3607), .ZN(n_8_0_3606));
   NOR2_X1 i_8_0_3762 (.A1(n_8_0_3609), .A2(n_8_0_3608), .ZN(n_8_0_3607));
   AOI211_X1 i_8_0_3763 (.A(n_8_0_537), .B(n_8_0_3653), .C1(n_8_0_4199), 
      .C2(n_8_0_4524), .ZN(n_8_0_3608));
   OR2_X1 i_8_0_3764 (.A1(\out_as[1] [5]), .A2(n_8_0_537), .ZN(n_8_0_1412));
   AOI21_X1 i_8_0_3765 (.A(n_8_0_6782), .B1(n_8_0_4524), .B2(n_8_0_4325), 
      .ZN(n_8_0_3609));
   INV_X1 i_8_0_3766 (.A(n_8_0_3611), .ZN(n_8_0_3610));
   AOI211_X1 i_8_0_3767 (.A(n_8_0_542), .B(n_8_0_3643), .C1(n_8_0_3697), 
      .C2(n_8_0_6593), .ZN(n_8_0_3611));
   OAI21_X1 i_8_0_3768 (.A(n_8_0_3614), .B1(n_8_0_3613), .B2(n_8_0_6611), 
      .ZN(n_8_0_3612));
   OAI21_X1 i_8_0_3769 (.A(n_8_0_4367), .B1(n_8_0_3638), .B2(n_8_0_532), 
      .ZN(n_8_0_3613));
   OAI21_X1 i_8_0_3770 (.A(n_8_0_6772), .B1(n_8_0_3640), .B2(n_8_0_532), 
      .ZN(n_8_0_3614));
   OR2_X1 i_8_0_3771 (.A1(\out_as[2] [5]), .A2(n_8_0_532), .ZN(n_8_0_1413));
   AOI21_X1 i_8_0_3773 (.A(n_8_0_3620), .B1(n_8_0_3619), .B2(n_8_0_6676), 
      .ZN(n_8_0_3616));
   NOR2_X1 i_8_0_3774 (.A1(n_8_0_3620), .A2(n_8_0_3618), .ZN(n_8_0_3617));
   NOR3_X1 i_8_0_3775 (.A1(n_8_0_7022), .A2(n_8_0_7021), .A3(n_8_0_3664), 
      .ZN(n_8_0_3618));
   NOR2_X1 i_8_0_3776 (.A1(n_8_0_7022), .A2(n_8_0_3664), .ZN(n_8_0_3619));
   AOI21_X1 i_8_0_3777 (.A(n_8_0_3664), .B1(n_8_0_4110), .B2(n_8_0_6828), 
      .ZN(n_8_0_3620));
   NAND2_X1 i_8_0_3778 (.A1(\out_bs[5] [3]), .A2(n_8_0_3622), .ZN(n_8_0_3621));
   INV_X1 i_8_0_3779 (.A(n_8_0_3623), .ZN(n_8_0_3622));
   NAND2_X1 i_8_0_3780 (.A1(\out_bs[5] [4]), .A2(n_8_0_6825), .ZN(n_8_0_3623));
   OAI21_X1 i_8_0_3782 (.A(n_8_0_3626), .B1(n_8_0_3627), .B2(n_8_0_6580), 
      .ZN(n_8_0_3625));
   OAI21_X1 i_8_0_3783 (.A(n_8_0_6837), .B1(n_8_0_3676), .B2(n_8_0_527), 
      .ZN(n_8_0_3626));
   OAI21_X1 i_8_0_3784 (.A(n_8_0_3686), .B1(n_8_0_3673), .B2(n_8_0_527), 
      .ZN(n_8_0_3627));
   AOI221_X1 i_8_0_3785 (.A(n_8_0_4059), .B1(n_8_0_3670), .B2(n_8_0_3629), 
      .C1(n_8_0_6623), .C2(n_8_0_6640), .ZN(n_8_0_3628));
   AOI21_X1 i_8_0_3786 (.A(n_8_0_522), .B1(n_8_0_5460), .B2(n_8_0_5442), 
      .ZN(n_8_0_3629));
   OR2_X1 i_8_0_3787 (.A1(\out_as[4] [5]), .A2(n_8_0_522), .ZN(n_8_0_1414));
   INV_X1 i_8_0_3788 (.A(n_8_0_3631), .ZN(n_8_0_3630));
   NOR2_X1 i_8_0_3789 (.A1(n_8_0_3633), .A2(n_8_0_3632), .ZN(n_8_0_3631));
   AOI211_X1 i_8_0_3790 (.A(n_8_0_512), .B(n_8_0_3646), .C1(n_8_0_4561), 
      .C2(n_8_0_6741), .ZN(n_8_0_3632));
   OR2_X1 i_8_0_3791 (.A1(\out_as[6] [5]), .A2(n_8_0_512), .ZN(n_8_0_1415));
   AOI21_X1 i_8_0_3792 (.A(n_8_0_6755), .B1(n_8_0_6741), .B2(n_8_0_4563), 
      .ZN(n_8_0_3633));
   AOI21_X1 i_8_0_3793 (.A(n_8_0_6853), .B1(n_8_0_3648), .B2(n_8_0_3634), 
      .ZN(n_127));
   NOR4_X1 i_8_0_3794 (.A1(n_8_0_3635), .A2(n_8_0_3636), .A3(n_8_0_3642), 
      .A4(n_8_0_4133), .ZN(n_8_0_3634));
   OAI21_X1 i_8_0_3795 (.A(n_8_0_3644), .B1(n_8_0_3643), .B2(n_8_0_3697), 
      .ZN(n_8_0_3635));
   OAI21_X1 i_8_0_3796 (.A(n_8_0_3638), .B1(n_8_0_3637), .B2(n_8_0_3639), 
      .ZN(n_8_0_3636));
   NOR2_X1 i_8_0_3797 (.A1(n_8_0_6704), .A2(n_8_0_4366), .ZN(n_8_0_3637));
   NAND2_X1 i_8_0_3798 (.A1(n_8_0_6775), .A2(n_8_0_3641), .ZN(n_8_0_3638));
   NOR2_X1 i_8_0_3799 (.A1(n_8_0_6773), .A2(n_8_0_3641), .ZN(n_8_0_3639));
   NAND2_X1 i_8_0_3800 (.A1(n_8_0_7066), .A2(n_8_0_7065), .ZN(n_8_0_3640));
   NOR2_X1 i_8_0_3801 (.A1(\out_as[2] [6]), .A2(\out_as[2] [5]), .ZN(n_8_0_3641));
   AOI211_X1 i_8_0_3802 (.A(n_8_0_6665), .B(n_8_0_6662), .C1(n_8_0_6811), 
      .C2(n_8_0_3643), .ZN(n_8_0_3642));
   NAND2_X1 i_8_0_3803 (.A1(n_8_0_7089), .A2(n_8_0_7088), .ZN(n_8_0_3643));
   OAI22_X1 i_8_0_3804 (.A1(n_8_0_6754), .A2(n_8_0_3647), .B1(n_8_0_3645), 
      .B2(n_8_0_5454), .ZN(n_8_0_3644));
   OAI21_X1 i_8_0_3805 (.A(n_8_0_4563), .B1(n_8_0_3646), .B2(n_8_0_6765), 
      .ZN(n_8_0_3645));
   NAND2_X1 i_8_0_3806 (.A1(n_8_0_7018), .A2(n_8_0_7017), .ZN(n_8_0_3646));
   NOR2_X1 i_8_0_3807 (.A1(\out_as[6] [6]), .A2(\out_as[6] [5]), .ZN(n_8_0_3647));
   NOR4_X1 i_8_0_3808 (.A1(n_8_0_3660), .A2(n_8_0_3655), .A3(n_8_0_3666), 
      .A4(n_8_0_3649), .ZN(n_8_0_3648));
   AOI21_X1 i_8_0_3809 (.A(n_8_0_3652), .B1(n_8_0_3650), .B2(n_8_0_4231), 
      .ZN(n_8_0_3649));
   AOI21_X1 i_8_0_3810 (.A(n_8_0_6688), .B1(n_8_0_4198), .B2(n_8_0_3654), 
      .ZN(n_8_0_3650));
   NAND2_X1 i_8_0_3811 (.A1(n_8_0_6782), .A2(n_8_0_3653), .ZN(n_8_0_3651));
   NOR2_X1 i_8_0_3812 (.A1(n_8_0_6781), .A2(n_8_0_3654), .ZN(n_8_0_3652));
   NAND2_X1 i_8_0_3813 (.A1(n_8_0_7078), .A2(n_8_0_7077), .ZN(n_8_0_3653));
   NOR2_X1 i_8_0_3814 (.A1(\out_as[1] [6]), .A2(\out_as[1] [5]), .ZN(n_8_0_3654));
   NAND2_X1 i_8_0_3815 (.A1(n_8_0_3657), .A2(n_8_0_3656), .ZN(n_8_0_3655));
   OAI22_X1 i_8_0_3816 (.A1(n_8_0_6729), .A2(n_8_0_3659), .B1(n_8_0_4423), 
      .B2(n_8_0_6719), .ZN(n_8_0_3656));
   AOI22_X1 i_8_0_3820 (.A1(n_8_0_6824), .A2(n_8_0_3664), .B1(n_8_0_3662), 
      .B2(n_8_0_3661), .ZN(n_8_0_3660));
   AOI21_X1 i_8_0_3821 (.A(n_8_0_4109), .B1(n_8_0_6674), .B2(\out_bs[5] [4]), 
      .ZN(n_8_0_3661));
   NAND2_X1 i_8_0_3822 (.A1(n_8_0_6832), .A2(n_8_0_3665), .ZN(n_8_0_3662));
   NAND2_X1 i_8_0_3823 (.A1(n_8_0_6824), .A2(n_8_0_3664), .ZN(n_8_0_3663));
   NAND2_X1 i_8_0_3824 (.A1(n_8_0_7030), .A2(n_8_0_7029), .ZN(n_8_0_3664));
   NOR2_X1 i_8_0_3825 (.A1(\out_as[5] [6]), .A2(\out_as[5] [5]), .ZN(n_8_0_3665));
   NAND2_X1 i_8_0_3826 (.A1(n_8_0_3667), .A2(n_8_0_3671), .ZN(n_8_0_3666));
   OAI21_X1 i_8_0_3827 (.A(n_8_0_3668), .B1(n_8_0_3670), .B2(n_8_0_6794), 
      .ZN(n_8_0_3667));
   OAI211_X1 i_8_0_3828 (.A(n_8_0_5462), .B(n_8_0_7035), .C1(n_8_0_6803), 
      .C2(n_8_0_3669), .ZN(n_8_0_3668));
   OR2_X1 i_8_0_3829 (.A1(\out_as[4] [6]), .A2(\out_as[4] [5]), .ZN(n_8_0_3669));
   NOR2_X1 i_8_0_3830 (.A1(\out_as[4] [6]), .A2(\out_as[4] [5]), .ZN(n_8_0_3670));
   OAI22_X1 i_8_0_3831 (.A1(n_8_0_6838), .A2(n_8_0_3677), .B1(n_8_0_3674), 
      .B2(n_8_0_3672), .ZN(n_8_0_3671));
   NAND2_X1 i_8_0_3832 (.A1(n_8_0_5466), .A2(n_8_0_3686), .ZN(n_8_0_3672));
   NAND2_X1 i_8_0_3833 (.A1(n_8_0_3675), .A2(n_8_0_3677), .ZN(n_8_0_3673));
   AOI21_X1 i_8_0_3834 (.A(n_8_0_3676), .B1(n_8_0_3686), .B2(n_8_0_6847), 
      .ZN(n_8_0_3674));
   NAND2_X1 i_8_0_3835 (.A1(n_8_0_6847), .A2(n_8_0_3686), .ZN(n_8_0_3675));
   NAND2_X1 i_8_0_3836 (.A1(n_8_0_7053), .A2(n_8_0_7052), .ZN(n_8_0_3676));
   NOR2_X1 i_8_0_3837 (.A1(\out_as[3] [6]), .A2(\out_as[3] [5]), .ZN(n_8_0_3677));
   NAND2_X1 i_8_0_3844 (.A1(n_8_0_6838), .A2(n_8_0_3685), .ZN(n_8_0_3683));
   NOR2_X1 i_8_0_3845 (.A1(n_8_0_6837), .A2(n_8_0_3686), .ZN(n_8_0_3684));
   NAND2_X1 i_8_0_3846 (.A1(n_8_0_7047), .A2(n_8_0_7046), .ZN(n_8_0_3685));
   NOR2_X1 i_8_0_3847 (.A1(\out_bs[3] [6]), .A2(\out_bs[3] [5]), .ZN(n_8_0_3686));
   AOI21_X1 i_8_0_3849 (.A(n_8_0_4107), .B1(n_8_0_4104), .B2(n_8_0_954), 
      .ZN(n_8_0_3688));
   OAI21_X1 i_8_0_3854 (.A(n_8_0_4231), .B1(n_8_0_4197), .B2(n_8_0_958), 
      .ZN(n_8_0_3693));
   NOR3_X1 i_8_0_3856 (.A1(\out_as[0] [6]), .A2(n_8_0_959), .A3(n_8_0_3697), 
      .ZN(n_8_0_3695));
   NAND2_X1 i_8_0_3857 (.A1(n_8_0_6816), .A2(n_8_0_4604), .ZN(n_8_0_3696));
   NOR2_X1 i_8_0_3858 (.A1(n_8_0_6815), .A2(n_8_0_4603), .ZN(n_8_0_3697));
   AOI21_X1 i_8_0_3862 (.A(n_8_0_4611), .B1(n_8_0_4565), .B2(n_8_0_5522), 
      .ZN(n_8_0_3700));
   OAI21_X1 i_8_0_3863 (.A(n_8_0_4346), .B1(n_8_0_5522), .B2(\out_bs[6] [6]), 
      .ZN(n_8_0_3701));
   AOI21_X1 i_8_0_3865 (.A(n_8_0_6514), .B1(n_8_0_5519), .B2(n_8_0_3704), 
      .ZN(n_8_0_3703));
   OAI21_X1 i_8_0_3866 (.A(n_8_0_4378), .B1(n_8_0_4551), .B2(n_8_0_946), 
      .ZN(n_8_0_3704));
   AOI21_X1 i_8_0_3868 (.A(n_8_0_6578), .B1(n_8_0_3707), .B2(n_8_0_5500), 
      .ZN(n_8_0_3706));
   AOI21_X1 i_8_0_3869 (.A(n_8_0_4592), .B1(n_8_0_6837), .B2(n_8_0_948), 
      .ZN(n_8_0_3707));
   OAI21_X1 i_8_0_3874 (.A(n_8_0_3713), .B1(n_8_0_3717), .B2(n_8_0_951), 
      .ZN(n_8_0_3712));
   AOI21_X1 i_8_0_3875 (.A(n_8_0_3714), .B1(n_8_0_5505), .B2(n_8_0_6597), 
      .ZN(n_8_0_3713));
   OAI211_X1 i_8_0_3876 (.A(n_8_0_6526), .B(n_8_0_3715), .C1(n_8_0_4579), 
      .C2(n_8_0_950), .ZN(n_8_0_3714));
   NAND2_X1 i_8_0_3877 (.A1(n_8_0_5525), .A2(n_8_0_3716), .ZN(n_8_0_3715));
   OAI21_X1 i_8_0_3878 (.A(n_8_0_6321), .B1(n_8_0_4525), .B2(n_8_0_950), 
      .ZN(n_8_0_3716));
   AOI21_X1 i_8_0_3879 (.A(n_8_0_4515), .B1(n_8_0_4513), .B2(n_8_0_5505), 
      .ZN(n_8_0_3717));
   OAI221_X1 i_8_0_3880 (.A(n_8_0_6606), .B1(n_8_0_4587), .B2(n_8_0_949), 
      .C1(n_8_0_3719), .C2(n_8_0_5515), .ZN(n_8_0_3718));
   INV_X1 i_8_0_3881 (.A(n_8_0_3720), .ZN(n_8_0_3719));
   OAI21_X1 i_8_0_3882 (.A(n_8_0_4499), .B1(n_8_0_4519), .B2(n_8_0_949), 
      .ZN(n_8_0_3720));
   OAI22_X1 i_8_0_3883 (.A1(n_8_0_3723), .A2(n_8_0_3722), .B1(n_8_0_947), 
      .B2(n_8_0_4542), .ZN(n_8_0_3721));
   NOR3_X1 i_8_0_3884 (.A1(n_8_0_6557), .A2(n_8_0_6352), .A3(n_8_0_5744), 
      .ZN(n_8_0_3722));
   INV_X1 i_8_0_3885 (.A(n_8_0_3724), .ZN(n_8_0_3723));
   OAI21_X1 i_8_0_3886 (.A(n_8_0_4058), .B1(n_8_0_4540), .B2(n_8_0_947), 
      .ZN(n_8_0_3724));
   AOI21_X1 i_8_0_3887 (.A(n_8_0_6853), .B1(n_8_0_3735), .B2(n_8_0_3725), 
      .ZN(n_128));
   NOR3_X1 i_8_0_3888 (.A1(n_8_0_3732), .A2(n_8_0_3729), .A3(n_8_0_3726), 
      .ZN(n_8_0_3725));
   OAI211_X1 i_8_0_3889 (.A(n_8_0_6556), .B(n_8_0_3727), .C1(n_8_0_4484), 
      .C2(n_8_0_5536), .ZN(n_8_0_3726));
   INV_X1 i_8_0_3890 (.A(n_8_0_3728), .ZN(n_8_0_3727));
   AOI211_X1 i_8_0_3891 (.A(n_8_0_939), .B(n_8_0_4383), .C1(n_8_0_4542), 
      .C2(n_8_0_5536), .ZN(n_8_0_3728));
   OAI221_X1 i_8_0_3892 (.A(n_8_0_6577), .B1(n_8_0_3730), .B2(n_8_0_4592), 
      .C1(n_8_0_940), .C2(n_8_0_4590), .ZN(n_8_0_3729));
   INV_X1 i_8_0_3893 (.A(n_8_0_3731), .ZN(n_8_0_3730));
   AOI21_X1 i_8_0_3894 (.A(n_8_0_5564), .B1(n_8_0_6837), .B2(n_8_0_940), 
      .ZN(n_8_0_3731));
   OAI21_X1 i_8_0_3895 (.A(n_8_0_3733), .B1(n_8_0_4595), .B2(n_8_0_936), 
      .ZN(n_8_0_3732));
   AOI21_X1 i_8_0_3896 (.A(n_8_0_6466), .B1(n_8_0_3734), .B2(n_8_0_5560), 
      .ZN(n_8_0_3733));
   AOI21_X1 i_8_0_3897 (.A(n_8_0_4599), .B1(n_8_0_6469), .B2(n_8_0_936), 
      .ZN(n_8_0_3734));
   NOR4_X1 i_8_0_3898 (.A1(n_8_0_3749), .A2(n_8_0_3742), .A3(n_8_0_3739), 
      .A4(n_8_0_3736), .ZN(n_8_0_3735));
   OAI21_X1 i_8_0_3899 (.A(n_8_0_3738), .B1(n_8_0_3737), .B2(n_8_0_937), 
      .ZN(n_8_0_3736));
   AOI21_X1 i_8_0_3900 (.A(n_8_0_4611), .B1(n_8_0_4565), .B2(n_8_0_5544), 
      .ZN(n_8_0_3737));
   OAI21_X1 i_8_0_3901 (.A(n_8_0_4346), .B1(n_8_0_5544), .B2(\out_bs[6] [6]), 
      .ZN(n_8_0_3738));
   OAI211_X1 i_8_0_3902 (.A(n_8_0_6513), .B(n_8_0_3740), .C1(n_8_0_4571), 
      .C2(n_8_0_938), .ZN(n_8_0_3739));
   OAI21_X1 i_8_0_3903 (.A(n_8_0_3741), .B1(n_8_0_6097), .B2(\out_bs[5] [4]), 
      .ZN(n_8_0_3740));
   OAI21_X1 i_8_0_3904 (.A(n_8_0_4378), .B1(n_8_0_4551), .B2(n_8_0_938), 
      .ZN(n_8_0_3741));
   OAI211_X1 i_8_0_3905 (.A(n_8_0_3746), .B(n_8_0_3743), .C1(n_8_0_5553), 
      .C2(n_8_0_4454), .ZN(n_8_0_3742));
   NAND2_X1 i_8_0_3906 (.A1(n_8_0_3745), .A2(n_8_0_3744), .ZN(n_8_0_3743));
   OAI21_X1 i_8_0_3907 (.A(n_8_0_6249), .B1(n_8_0_943), .B2(\out_as[0] [6]), 
      .ZN(n_8_0_3744));
   OAI21_X1 i_8_0_3908 (.A(n_8_0_5274), .B1(n_8_0_5553), .B2(n_8_0_7084), 
      .ZN(n_8_0_3745));
   NOR2_X1 i_8_0_3909 (.A1(n_8_0_3748), .A2(n_8_0_3747), .ZN(n_8_0_3746));
   OAI21_X1 i_8_0_3910 (.A(n_8_0_6606), .B1(n_8_0_6282), .B2(n_8_0_5552), 
      .ZN(n_8_0_3747));
   AOI211_X1 i_8_0_3911 (.A(n_8_0_941), .B(n_8_0_4125), .C1(n_8_0_4587), 
      .C2(n_8_0_5552), .ZN(n_8_0_3748));
   OAI221_X1 i_8_0_3912 (.A(n_8_0_6526), .B1(n_8_0_6321), .B2(n_8_0_5548), 
      .C1(n_8_0_3750), .C2(n_8_0_942), .ZN(n_8_0_3749));
   AOI21_X1 i_8_0_3913 (.A(n_8_0_4580), .B1(n_8_0_4526), .B2(n_8_0_5547), 
      .ZN(n_8_0_3750));
   INV_X1 i_8_0_3917 (.A(n_8_0_3754), .ZN(n_8_0_3753));
   AOI211_X1 i_8_0_3918 (.A(n_8_0_931), .B(n_8_0_4383), .C1(n_8_0_4542), 
      .C2(n_8_0_5573), .ZN(n_8_0_3754));
   OAI21_X1 i_8_0_3924 (.A(n_8_0_6480), .B1(n_8_0_4346), .B2(n_8_0_3761), 
      .ZN(n_8_0_3760));
   NOR3_X1 i_8_0_3925 (.A1(\out_as[6] [6]), .A2(n_8_0_929), .A3(n_8_0_4563), 
      .ZN(n_8_0_3761));
   OAI22_X1 i_8_0_3927 (.A1(n_8_0_3765), .A2(n_8_0_3764), .B1(n_8_0_930), 
      .B2(n_8_0_4573), .ZN(n_8_0_3763));
   NOR3_X1 i_8_0_3928 (.A1(n_8_0_6136), .A2(\out_bs[5] [4]), .A3(\out_bs[5] [6]), 
      .ZN(n_8_0_3764));
   NOR2_X1 i_8_0_3929 (.A1(n_8_0_3804), .A2(n_8_0_3766), .ZN(n_8_0_3765));
   NOR3_X1 i_8_0_3930 (.A1(\out_as[5] [6]), .A2(n_8_0_930), .A3(n_8_0_4110), 
      .ZN(n_8_0_3766));
   OAI21_X1 i_8_0_3931 (.A(n_8_0_3768), .B1(n_8_0_5581), .B2(n_8_0_6325), 
      .ZN(n_8_0_3767));
   AOI21_X1 i_8_0_3932 (.A(n_8_0_6578), .B1(n_8_0_3769), .B2(n_8_0_3770), 
      .ZN(n_8_0_3768));
   NOR2_X1 i_8_0_3933 (.A1(n_8_0_932), .A2(n_8_0_4472), .ZN(n_8_0_3769));
   NAND2_X1 i_8_0_3934 (.A1(n_8_0_4590), .A2(n_8_0_5581), .ZN(n_8_0_3770));
   OAI21_X1 i_8_0_3935 (.A(n_8_0_3779), .B1(n_8_0_3773), .B2(n_8_0_3772), 
      .ZN(n_8_0_3771));
   AOI211_X1 i_8_0_3936 (.A(\out_bs[0] [6]), .B(n_8_0_3775), .C1(n_8_0_5595), 
      .C2(\out_bs[0] [5]), .ZN(n_8_0_3772));
   INV_X1 i_8_0_3937 (.A(n_8_0_3774), .ZN(n_8_0_3773));
   OAI21_X1 i_8_0_3938 (.A(n_8_0_6811), .B1(n_8_0_935), .B2(\out_as[0] [6]), 
      .ZN(n_8_0_3774));
   NOR3_X1 i_8_0_3939 (.A1(\out_as[0] [6]), .A2(n_8_0_935), .A3(n_8_0_6816), 
      .ZN(n_8_0_3775));
   OAI21_X1 i_8_0_3940 (.A(n_8_0_3778), .B1(n_8_0_3777), .B2(n_8_0_934), 
      .ZN(n_8_0_3776));
   AOI21_X1 i_8_0_3941 (.A(n_8_0_4580), .B1(n_8_0_4526), .B2(n_8_0_5586), 
      .ZN(n_8_0_3777));
   OAI21_X1 i_8_0_3942 (.A(n_8_0_4232), .B1(n_8_0_5586), .B2(\out_bs[1] [6]), 
      .ZN(n_8_0_3778));
   AOI21_X1 i_8_0_3943 (.A(n_8_0_3780), .B1(n_8_0_3781), .B2(n_8_0_5589), 
      .ZN(n_8_0_3779));
   OAI21_X1 i_8_0_3944 (.A(n_8_0_6606), .B1(n_8_0_4587), .B2(n_8_0_933), 
      .ZN(n_8_0_3780));
   OAI21_X1 i_8_0_3945 (.A(n_8_0_4364), .B1(n_8_0_4125), .B2(n_8_0_933), 
      .ZN(n_8_0_3781));
   AOI21_X1 i_8_0_3946 (.A(n_8_0_6853), .B1(n_8_0_3807), .B2(n_8_0_3782), 
      .ZN(n_129));
   NOR4_X1 i_8_0_3947 (.A1(n_8_0_3805), .A2(n_8_0_3800), .A3(n_8_0_3792), 
      .A4(n_8_0_3783), .ZN(n_8_0_3782));
   OAI211_X1 i_8_0_3948 (.A(n_8_0_3784), .B(n_8_0_4131), .C1(n_8_0_927), 
      .C2(n_8_0_3791), .ZN(n_8_0_3783));
   AOI211_X1 i_8_0_3949 (.A(n_8_0_3789), .B(n_8_0_3785), .C1(n_8_0_6953), 
      .C2(n_8_0_3790), .ZN(n_8_0_3784));
   OAI221_X1 i_8_0_3950 (.A(n_8_0_6526), .B1(n_8_0_4579), .B2(n_8_0_926), 
      .C1(n_8_0_3786), .C2(n_8_0_5622), .ZN(n_8_0_3785));
   INV_X1 i_8_0_3951 (.A(n_8_0_3787), .ZN(n_8_0_3786));
   OAI21_X1 i_8_0_3952 (.A(n_8_0_6321), .B1(n_8_0_4525), .B2(n_8_0_926), 
      .ZN(n_8_0_3787));
   AOI21_X1 i_8_0_3953 (.A(n_8_0_3789), .B1(n_8_0_3790), .B2(n_8_0_6953), 
      .ZN(n_8_0_3788));
   OAI21_X1 i_8_0_3954 (.A(n_8_0_6606), .B1(n_8_0_6282), .B2(n_8_0_5615), 
      .ZN(n_8_0_3789));
   OAI21_X1 i_8_0_3955 (.A(n_8_0_4587), .B1(n_8_0_4519), .B2(n_8_0_5615), 
      .ZN(n_8_0_3790));
   AOI21_X1 i_8_0_3956 (.A(n_8_0_4128), .B1(n_8_0_4513), .B2(n_8_0_6175), 
      .ZN(n_8_0_3791));
   NAND3_X1 i_8_0_3957 (.A1(n_8_0_3799), .A2(n_8_0_3795), .A3(n_8_0_3793), 
      .ZN(n_8_0_3792));
   AOI211_X1 i_8_0_3958 (.A(n_8_0_6557), .B(n_8_0_3794), .C1(n_8_0_5606), 
      .C2(n_8_0_6799), .ZN(n_8_0_3793));
   AOI211_X1 i_8_0_3959 (.A(\out_as[4] [6]), .B(n_8_0_923), .C1(n_8_0_5460), 
      .C2(n_8_0_5605), .ZN(n_8_0_3794));
   AOI21_X1 i_8_0_3960 (.A(n_8_0_3796), .B1(n_8_0_3797), .B2(n_8_0_6729), 
      .ZN(n_8_0_3795));
   NOR4_X1 i_8_0_3961 (.A1(\out_as[7] [6]), .A2(n_8_0_920), .A3(n_8_0_4424), 
      .A4(n_8_0_3798), .ZN(n_8_0_3796));
   OAI22_X1 i_8_0_3962 (.A1(\out_as[7] [6]), .A2(n_8_0_920), .B1(n_8_0_4424), 
      .B2(n_8_0_3798), .ZN(n_8_0_3797));
   NOR3_X1 i_8_0_3963 (.A1(n_8_0_5975), .A2(\out_bs[7] [2]), .A3(\out_bs[7] [6]), 
      .ZN(n_8_0_3798));
   NAND2_X1 i_8_0_3964 (.A1(n_8_0_6597), .A2(n_8_0_6175), .ZN(n_8_0_3799));
   OAI21_X1 i_8_0_3965 (.A(n_8_0_3801), .B1(n_8_0_4573), .B2(n_8_0_922), 
      .ZN(n_8_0_3800));
   OAI22_X1 i_8_0_3966 (.A1(n_8_0_3804), .A2(n_8_0_3802), .B1(n_8_0_6165), 
      .B2(n_8_0_4105), .ZN(n_8_0_3801));
   NOR3_X1 i_8_0_3967 (.A1(\out_as[5] [6]), .A2(n_8_0_922), .A3(n_8_0_4110), 
      .ZN(n_8_0_3802));
   NAND2_X1 i_8_0_3968 (.A1(n_8_0_6826), .A2(n_8_0_4108), .ZN(n_8_0_3803));
   NOR2_X1 i_8_0_3969 (.A1(n_8_0_6824), .A2(n_8_0_4110), .ZN(n_8_0_3804));
   OAI221_X1 i_8_0_3970 (.A(n_8_0_6590), .B1(n_8_0_4610), .B2(n_8_0_921), 
      .C1(n_8_0_3806), .C2(n_8_0_5626), .ZN(n_8_0_3805));
   AOI21_X1 i_8_0_3971 (.A(n_8_0_4556), .B1(n_8_0_4565), .B2(n_8_0_6887), 
      .ZN(n_8_0_3806));
   AOI21_X1 i_8_0_3972 (.A(n_8_0_3809), .B1(n_8_0_3808), .B2(n_8_0_6160), 
      .ZN(n_8_0_3807));
   AOI21_X1 i_8_0_3973 (.A(n_8_0_4592), .B1(n_8_0_6325), .B2(n_8_0_924), 
      .ZN(n_8_0_3808));
   OAI211_X1 i_8_0_3974 (.A(n_8_0_6577), .B(n_8_0_4307), .C1(n_8_0_4306), 
      .C2(n_8_0_924), .ZN(n_8_0_3809));
   AOI21_X1 i_8_0_3979 (.A(n_8_0_3814), .B1(n_8_0_3815), .B2(n_8_0_6550), 
      .ZN(n_8_0_3813));
   OAI21_X1 i_8_0_3980 (.A(n_8_0_3916), .B1(n_8_0_3994), .B2(n_8_0_913), 
      .ZN(n_8_0_3814));
   OAI21_X1 i_8_0_3981 (.A(n_8_0_4555), .B1(n_8_0_4564), .B2(n_8_0_913), 
      .ZN(n_8_0_3815));
   OAI211_X1 i_8_0_3982 (.A(n_8_0_6577), .B(n_8_0_3817), .C1(n_8_0_4590), 
      .C2(n_8_0_916), .ZN(n_8_0_3816));
   OAI21_X1 i_8_0_3983 (.A(n_8_0_3818), .B1(n_8_0_6007), .B2(n_8_0_6565), 
      .ZN(n_8_0_3817));
   AOI21_X1 i_8_0_3984 (.A(n_8_0_4592), .B1(n_8_0_6837), .B2(n_8_0_916), 
      .ZN(n_8_0_3818));
   AOI211_X1 i_8_0_3988 (.A(n_8_0_4107), .B(n_8_0_3823), .C1(n_8_0_4104), 
      .C2(n_8_0_914), .ZN(n_8_0_3822));
   NOR2_X1 i_8_0_3989 (.A1(n_8_0_6210), .A2(n_8_0_3824), .ZN(n_8_0_3823));
   OAI21_X1 i_8_0_3990 (.A(n_8_0_4106), .B1(n_8_0_4573), .B2(n_8_0_914), 
      .ZN(n_8_0_3824));
   AOI21_X1 i_8_0_3991 (.A(n_8_0_5653), .B1(n_8_0_3826), .B2(n_8_0_6596), 
      .ZN(n_8_0_3825));
   OR2_X1 i_8_0_3992 (.A1(n_8_0_4512), .A2(n_8_0_919), .ZN(n_8_0_3826));
   NAND3_X1 i_8_0_3993 (.A1(n_8_0_6606), .A2(n_8_0_3830), .A3(n_8_0_3828), 
      .ZN(n_8_0_3827));
   OR2_X1 i_8_0_3994 (.A1(n_8_0_917), .A2(n_8_0_3829), .ZN(n_8_0_3828));
   AOI21_X1 i_8_0_3995 (.A(n_8_0_4588), .B1(n_8_0_4520), .B2(n_8_0_5642), 
      .ZN(n_8_0_3829));
   NAND2_X1 i_8_0_3996 (.A1(n_8_0_4498), .A2(n_8_0_5642), .ZN(n_8_0_3830));
   OAI211_X1 i_8_0_3997 (.A(n_8_0_3832), .B(n_8_0_6249), .C1(n_8_0_919), 
      .C2(n_8_0_4514), .ZN(n_8_0_3831));
   AOI21_X1 i_8_0_3998 (.A(n_8_0_3833), .B1(n_8_0_3834), .B2(n_8_0_5647), 
      .ZN(n_8_0_3832));
   OAI21_X1 i_8_0_3999 (.A(n_8_0_6526), .B1(n_8_0_4579), .B2(n_8_0_918), 
      .ZN(n_8_0_3833));
   OAI21_X1 i_8_0_4000 (.A(n_8_0_6321), .B1(n_8_0_4525), .B2(n_8_0_918), 
      .ZN(n_8_0_3834));
   NAND2_X1 i_8_0_4002 (.A1(n_8_0_3837), .A2(n_8_0_6560), .ZN(n_8_0_3836));
   AOI21_X1 i_8_0_4003 (.A(n_8_0_4487), .B1(n_8_0_6795), .B2(n_8_0_3838), 
      .ZN(n_8_0_3837));
   OR2_X1 i_8_0_4004 (.A1(\out_as[4] [6]), .A2(n_8_0_915), .ZN(n_8_0_3838));
   NOR3_X1 i_8_0_4008 (.A1(n_8_0_3842), .A2(n_8_0_6250), .A3(n_8_0_3851), 
      .ZN(n_8_0_3841));
   OAI21_X1 i_8_0_4009 (.A(n_8_0_3843), .B1(n_8_0_4514), .B2(n_8_0_911), 
      .ZN(n_8_0_3842));
   INV_X1 i_8_0_4010 (.A(n_8_0_3844), .ZN(n_8_0_3843));
   OAI211_X1 i_8_0_4011 (.A(n_8_0_6556), .B(n_8_0_3845), .C1(n_8_0_4484), 
      .C2(n_8_0_5691), .ZN(n_8_0_3844));
   INV_X1 i_8_0_4012 (.A(n_8_0_3846), .ZN(n_8_0_3845));
   AOI211_X1 i_8_0_4013 (.A(n_8_0_907), .B(n_8_0_4383), .C1(n_8_0_5460), 
      .C2(n_8_0_5691), .ZN(n_8_0_3846));
   OAI21_X1 i_8_0_4014 (.A(n_8_0_3848), .B1(n_8_0_5943), .B2(n_8_0_6668), 
      .ZN(n_8_0_3847));
   OAI21_X1 i_8_0_4015 (.A(n_8_0_6596), .B1(n_8_0_4512), .B2(n_8_0_911), 
      .ZN(n_8_0_3848));
   AOI211_X1 i_8_0_4016 (.A(n_8_0_6607), .B(n_8_0_3850), .C1(n_8_0_5664), 
      .C2(n_8_0_6283), .ZN(n_8_0_3849));
   AOI211_X1 i_8_0_4017 (.A(n_8_0_909), .B(n_8_0_4125), .C1(n_8_0_4587), 
      .C2(n_8_0_5665), .ZN(n_8_0_3850));
   OAI221_X1 i_8_0_4018 (.A(n_8_0_6526), .B1(n_8_0_6321), .B2(n_8_0_5669), 
      .C1(n_8_0_3852), .C2(n_8_0_910), .ZN(n_8_0_3851));
   AOI21_X1 i_8_0_4019 (.A(n_8_0_4580), .B1(n_8_0_4526), .B2(n_8_0_5668), 
      .ZN(n_8_0_3852));
   NOR2_X1 i_8_0_4023 (.A1(n_8_0_3857), .A2(n_8_0_6514), .ZN(n_8_0_3856));
   OAI22_X1 i_8_0_4024 (.A1(n_8_0_5682), .A2(n_8_0_3858), .B1(n_8_0_4571), 
      .B2(n_8_0_906), .ZN(n_8_0_3857));
   INV_X1 i_8_0_4025 (.A(n_8_0_3859), .ZN(n_8_0_3858));
   OAI21_X1 i_8_0_4026 (.A(n_8_0_4378), .B1(n_8_0_4551), .B2(n_8_0_906), 
      .ZN(n_8_0_3859));
   AOI21_X1 i_8_0_4027 (.A(n_8_0_3861), .B1(n_8_0_5687), .B2(n_8_0_6326), 
      .ZN(n_8_0_3860));
   OAI21_X1 i_8_0_4028 (.A(n_8_0_6577), .B1(n_8_0_3862), .B2(n_8_0_908), 
      .ZN(n_8_0_3861));
   AOI21_X1 i_8_0_4029 (.A(n_8_0_4591), .B1(n_8_0_4593), .B2(n_8_0_5687), 
      .ZN(n_8_0_3862));
   AOI21_X1 i_8_0_4031 (.A(n_8_0_4611), .B1(n_8_0_4565), .B2(n_8_0_5677), 
      .ZN(n_8_0_3864));
   OAI21_X1 i_8_0_4032 (.A(n_8_0_4346), .B1(n_8_0_5677), .B2(\out_bs[6] [6]), 
      .ZN(n_8_0_3865));
   AOI22_X1 i_8_0_4035 (.A1(n_8_0_3869), .A2(n_8_0_3868), .B1(n_8_0_5727), 
      .B2(n_8_0_5460), .ZN(n_8_0_3867));
   OR2_X1 i_8_0_4036 (.A1(n_8_0_899), .A2(n_8_0_4383), .ZN(n_8_0_3868));
   OAI21_X1 i_8_0_4037 (.A(n_8_0_4059), .B1(n_8_0_5728), .B2(\out_bs[4] [6]), 
      .ZN(n_8_0_3869));
   INV_X1 i_8_0_4038 (.A(n_8_0_3871), .ZN(n_8_0_3870));
   OAI21_X1 i_8_0_4039 (.A(n_8_0_3873), .B1(n_8_0_3872), .B2(n_8_0_897), 
      .ZN(n_8_0_3871));
   OAI21_X1 i_8_0_4040 (.A(n_8_0_4559), .B1(n_8_0_4611), .B2(n_8_0_5722), 
      .ZN(n_8_0_3872));
   OAI21_X1 i_8_0_4041 (.A(n_8_0_4346), .B1(n_8_0_5722), .B2(\out_bs[6] [6]), 
      .ZN(n_8_0_3873));
   OAI221_X1 i_8_0_4042 (.A(n_8_0_6577), .B1(n_8_0_6325), .B2(n_8_0_5696), 
      .C1(n_8_0_3875), .C2(n_8_0_900), .ZN(n_8_0_3874));
   AOI21_X1 i_8_0_4043 (.A(n_8_0_4591), .B1(n_8_0_4593), .B2(n_8_0_5697), 
      .ZN(n_8_0_3875));
   AOI21_X1 i_8_0_4047 (.A(n_8_0_4580), .B1(n_8_0_4526), .B2(n_8_0_5711), 
      .ZN(n_8_0_3879));
   NAND3_X1 i_8_0_4048 (.A1(n_8_0_6781), .A2(n_8_0_5711), .A3(\out_bs[1] [5]), 
      .ZN(n_8_0_3880));
   AOI21_X1 i_8_0_4056 (.A(n_8_0_4588), .B1(n_8_0_4520), .B2(n_8_0_5706), 
      .ZN(n_8_0_3888));
   OAI211_X1 i_8_0_4058 (.A(n_8_0_3891), .B(\out_bs[5] [5]), .C1(\out_bs[5] [4]), 
      .C2(n_8_0_6299), .ZN(n_8_0_3890));
   OAI21_X1 i_8_0_4059 (.A(n_8_0_6824), .B1(n_8_0_898), .B2(\out_as[5] [6]), 
      .ZN(n_8_0_3891));
   AOI211_X1 i_8_0_4063 (.A(n_8_0_6527), .B(n_8_0_4580), .C1(n_8_0_4526), 
      .C2(n_8_0_5983), .ZN(n_8_0_3894));
   AOI21_X1 i_8_0_4065 (.A(n_8_0_6557), .B1(n_8_0_4485), .B2(n_8_0_5744), 
      .ZN(n_8_0_3896));
   OR2_X1 i_8_0_4066 (.A1(\out_as[4] [6]), .A2(n_8_0_891), .ZN(n_8_0_3897));
   AOI21_X1 i_8_0_4067 (.A(n_8_0_5459), .B1(n_8_0_5744), .B2(\out_bs[4] [5]), 
      .ZN(n_8_0_3898));
   NOR2_X1 i_8_0_4069 (.A1(n_8_0_4105), .A2(\out_bs[5] [3]), .ZN(n_8_0_3900));
   INV_X1 i_8_0_4070 (.A(n_8_0_3902), .ZN(n_8_0_3901));
   OAI21_X1 i_8_0_4071 (.A(n_8_0_6824), .B1(n_8_0_890), .B2(\out_as[5] [6]), 
      .ZN(n_8_0_3902));
   OAI221_X1 i_8_0_4077 (.A(n_8_0_6249), .B1(n_8_0_5944), .B2(n_8_0_4454), 
      .C1(n_8_0_3909), .C2(n_8_0_895), .ZN(n_8_0_3908));
   AOI21_X1 i_8_0_4078 (.A(n_8_0_4515), .B1(n_8_0_4513), .B2(n_8_0_5943), 
      .ZN(n_8_0_3909));
   OAI21_X1 i_8_0_4079 (.A(n_8_0_3911), .B1(n_8_0_3912), .B2(n_8_0_893), 
      .ZN(n_8_0_3910));
   OAI21_X1 i_8_0_4080 (.A(n_8_0_4365), .B1(n_8_0_5814), .B2(\out_bs[2] [6]), 
      .ZN(n_8_0_3911));
   AOI21_X1 i_8_0_4081 (.A(n_8_0_4588), .B1(n_8_0_4520), .B2(n_8_0_5814), 
      .ZN(n_8_0_3912));
   OAI221_X1 i_8_0_4082 (.A(n_8_0_6577), .B1(n_8_0_6325), .B2(n_8_0_6008), 
      .C1(n_8_0_3955), .C2(n_8_0_892), .ZN(n_8_0_3913));
   INV_X1 i_8_0_4083 (.A(n_8_0_3915), .ZN(n_8_0_3914));
   OAI21_X1 i_8_0_4084 (.A(n_8_0_3916), .B1(n_8_0_3994), .B2(n_8_0_889), 
      .ZN(n_8_0_3915));
   AOI21_X1 i_8_0_4085 (.A(n_8_0_6591), .B1(n_8_0_4349), .B2(n_8_0_5893), 
      .ZN(n_8_0_3916));
   OAI211_X1 i_8_0_4090 (.A(n_8_0_3925), .B(n_8_0_3938), .C1(n_8_0_887), 
      .C2(n_8_0_3937), .ZN(n_8_0_3920));
   OAI221_X1 i_8_0_4091 (.A(n_8_0_6590), .B1(n_8_0_5768), .B2(n_8_0_4555), 
      .C1(n_8_0_3922), .C2(n_8_0_881), .ZN(n_8_0_3921));
   OAI21_X1 i_8_0_4092 (.A(n_8_0_4559), .B1(n_8_0_4611), .B2(n_8_0_5767), 
      .ZN(n_8_0_3922));
   AOI21_X1 i_8_0_4094 (.A(n_8_0_4591), .B1(n_8_0_4593), .B2(n_8_0_5787), 
      .ZN(n_8_0_3924));
   AOI21_X1 i_8_0_4095 (.A(n_8_0_6527), .B1(n_8_0_3927), .B2(n_8_0_3926), 
      .ZN(n_8_0_3925));
   OAI22_X1 i_8_0_4096 (.A1(n_8_0_4579), .A2(n_8_0_886), .B1(n_8_0_4582), 
      .B2(n_8_0_5758), .ZN(n_8_0_3926));
   NAND2_X1 i_8_0_4097 (.A1(n_8_0_886), .A2(n_8_0_5397), .ZN(n_8_0_3927));
   OAI21_X1 i_8_0_4099 (.A(n_8_0_5782), .B1(n_8_0_4485), .B2(n_8_0_3930), 
      .ZN(n_8_0_3929));
   NOR3_X1 i_8_0_4100 (.A1(\out_as[4] [6]), .A2(n_8_0_883), .A3(n_8_0_4487), 
      .ZN(n_8_0_3930));
   OAI211_X1 i_8_0_4101 (.A(n_8_0_6513), .B(n_8_0_3932), .C1(n_8_0_4571), 
      .C2(n_8_0_882), .ZN(n_8_0_3931));
   OAI21_X1 i_8_0_4102 (.A(n_8_0_3933), .B1(n_8_0_6374), .B2(\out_bs[5] [4]), 
      .ZN(n_8_0_3932));
   OAI22_X1 i_8_0_4103 (.A1(n_8_0_6828), .A2(n_8_0_4576), .B1(n_8_0_4551), 
      .B2(n_8_0_882), .ZN(n_8_0_3933));
   INV_X1 i_8_0_4105 (.A(n_8_0_3936), .ZN(n_8_0_3935));
   OAI21_X1 i_8_0_4106 (.A(n_8_0_6282), .B1(n_8_0_4519), .B2(n_8_0_885), 
      .ZN(n_8_0_3936));
   AOI21_X1 i_8_0_4107 (.A(n_8_0_4515), .B1(n_8_0_4513), .B2(n_8_0_5771), 
      .ZN(n_8_0_3937));
   OAI21_X1 i_8_0_4108 (.A(n_8_0_4133), .B1(n_8_0_5771), .B2(n_8_0_6250), 
      .ZN(n_8_0_3938));
   AOI21_X1 i_8_0_4112 (.A(n_8_0_6853), .B1(n_8_0_3967), .B2(n_8_0_3942), 
      .ZN(n_130));
   NOR3_X1 i_8_0_4113 (.A1(n_8_0_3957), .A2(n_8_0_3953), .A3(n_8_0_3943), 
      .ZN(n_8_0_3942));
   OAI211_X1 i_8_0_4114 (.A(n_8_0_3944), .B(n_8_0_6249), .C1(n_8_0_5804), 
      .C2(n_8_0_4454), .ZN(n_8_0_3943));
   NOR3_X1 i_8_0_4115 (.A1(n_8_0_3950), .A2(n_8_0_3945), .A3(n_8_0_3948), 
      .ZN(n_8_0_3944));
   OAI221_X1 i_8_0_4116 (.A(n_8_0_6526), .B1(n_8_0_3946), .B2(n_8_0_5819), 
      .C1(n_8_0_878), .C2(n_8_0_4579), .ZN(n_8_0_3945));
   INV_X1 i_8_0_4117 (.A(n_8_0_3947), .ZN(n_8_0_3946));
   OAI21_X1 i_8_0_4118 (.A(n_8_0_6321), .B1(n_8_0_4525), .B2(n_8_0_878), 
      .ZN(n_8_0_3947));
   AOI21_X1 i_8_0_4119 (.A(n_8_0_879), .B1(n_8_0_4514), .B2(n_8_0_3949), 
      .ZN(n_8_0_3948));
   NAND2_X1 i_8_0_4120 (.A1(n_8_0_5805), .A2(n_8_0_4513), .ZN(n_8_0_3949));
   OAI21_X1 i_8_0_4121 (.A(n_8_0_3951), .B1(n_8_0_4587), .B2(n_8_0_877), 
      .ZN(n_8_0_3950));
   AOI21_X1 i_8_0_4122 (.A(n_8_0_6607), .B1(n_8_0_5813), .B2(n_8_0_3952), 
      .ZN(n_8_0_3951));
   OAI21_X1 i_8_0_4123 (.A(n_8_0_4499), .B1(n_8_0_4519), .B2(n_8_0_877), 
      .ZN(n_8_0_3952));
   OAI21_X1 i_8_0_4124 (.A(n_8_0_3954), .B1(n_8_0_3956), .B2(n_8_0_876), 
      .ZN(n_8_0_3953));
   AOI21_X1 i_8_0_4125 (.A(n_8_0_6578), .B1(n_8_0_6326), .B2(n_8_0_5793), 
      .ZN(n_8_0_3954));
   AOI21_X1 i_8_0_4126 (.A(n_8_0_4591), .B1(n_8_0_4593), .B2(n_8_0_6007), 
      .ZN(n_8_0_3955));
   AOI21_X1 i_8_0_4127 (.A(n_8_0_4591), .B1(n_8_0_4593), .B2(n_8_0_5793), 
      .ZN(n_8_0_3956));
   NAND3_X1 i_8_0_4128 (.A1(n_8_0_3961), .A2(n_8_0_3958), .A3(n_8_0_3964), 
      .ZN(n_8_0_3957));
   NOR2_X1 i_8_0_4129 (.A1(n_8_0_3960), .A2(n_8_0_3959), .ZN(n_8_0_3958));
   OAI21_X1 i_8_0_4130 (.A(n_8_0_6590), .B1(n_8_0_4348), .B2(n_8_0_5823), 
      .ZN(n_8_0_3959));
   AOI211_X1 i_8_0_4131 (.A(n_8_0_873), .B(n_8_0_4558), .C1(n_8_0_4610), 
      .C2(n_8_0_5823), .ZN(n_8_0_3960));
   OAI21_X1 i_8_0_4132 (.A(n_8_0_3962), .B1(n_8_0_3963), .B2(n_8_0_6409), 
      .ZN(n_8_0_3961));
   AOI21_X1 i_8_0_4133 (.A(n_8_0_4107), .B1(n_8_0_4104), .B2(n_8_0_874), 
      .ZN(n_8_0_3962));
   OAI21_X1 i_8_0_4134 (.A(n_8_0_4106), .B1(n_8_0_4573), .B2(n_8_0_874), 
      .ZN(n_8_0_3963));
   AOI21_X1 i_8_0_4135 (.A(n_8_0_3965), .B1(n_8_0_4485), .B2(n_8_0_5799), 
      .ZN(n_8_0_3964));
   OAI21_X1 i_8_0_4136 (.A(n_8_0_6556), .B1(n_8_0_3966), .B2(n_8_0_875), 
      .ZN(n_8_0_3965));
   AOI21_X1 i_8_0_4137 (.A(n_8_0_4543), .B1(n_8_0_4099), .B2(n_8_0_5799), 
      .ZN(n_8_0_3966));
   AOI21_X1 i_8_0_4138 (.A(n_8_0_4409), .B1(n_8_0_3969), .B2(n_8_0_3968), 
      .ZN(n_8_0_3967));
   OAI21_X1 i_8_0_4139 (.A(n_8_0_872), .B1(n_8_0_6469), .B2(n_8_0_6403), 
      .ZN(n_8_0_3968));
   OAI21_X1 i_8_0_4140 (.A(n_8_0_4503), .B1(n_8_0_4599), .B2(n_8_0_6403), 
      .ZN(n_8_0_3969));
   AOI21_X1 i_8_0_4141 (.A(n_8_0_6853), .B1(n_8_0_3973), .B2(n_8_0_3970), 
      .ZN(n_131));
   NOR4_X1 i_8_0_4142 (.A1(n_8_0_3986), .A2(n_8_0_3981), .A3(n_8_0_3976), 
      .A4(n_8_0_3971), .ZN(n_8_0_3970));
   OR2_X1 i_8_0_4143 (.A1(n_8_0_3992), .A2(n_8_0_3972), .ZN(n_8_0_3971));
   OAI221_X1 i_8_0_4144 (.A(n_8_0_6249), .B1(n_8_0_5854), .B2(n_8_0_4454), 
      .C1(n_8_0_3984), .C2(n_8_0_871), .ZN(n_8_0_3972));
   NOR3_X1 i_8_0_4145 (.A1(n_8_0_3989), .A2(n_8_0_3979), .A3(n_8_0_3974), 
      .ZN(n_8_0_3973));
   OAI221_X1 i_8_0_4146 (.A(n_8_0_6556), .B1(n_8_0_5836), .B2(n_8_0_4484), 
      .C1(n_8_0_3975), .C2(n_8_0_867), .ZN(n_8_0_3974));
   AOI21_X1 i_8_0_4147 (.A(n_8_0_4543), .B1(n_8_0_4099), .B2(n_8_0_5835), 
      .ZN(n_8_0_3975));
   AOI22_X1 i_8_0_4148 (.A1(n_8_0_3977), .A2(n_8_0_6513), .B1(n_8_0_6828), 
      .B2(n_8_0_866), .ZN(n_8_0_3976));
   AOI21_X1 i_8_0_4149 (.A(n_8_0_3978), .B1(n_8_0_4572), .B2(n_8_0_6901), 
      .ZN(n_8_0_3977));
   AOI21_X1 i_8_0_4150 (.A(n_8_0_4576), .B1(n_8_0_6459), .B2(n_8_0_7022), 
      .ZN(n_8_0_3978));
   OAI221_X1 i_8_0_4151 (.A(n_8_0_6577), .B1(n_8_0_6325), .B2(n_8_0_5859), 
      .C1(n_8_0_3980), .C2(n_8_0_868), .ZN(n_8_0_3979));
   AOI21_X1 i_8_0_4152 (.A(n_8_0_4591), .B1(n_8_0_4593), .B2(n_8_0_5858), 
      .ZN(n_8_0_3980));
   OAI211_X1 i_8_0_4153 (.A(n_8_0_6526), .B(n_8_0_3982), .C1(n_8_0_4579), 
      .C2(n_8_0_870), .ZN(n_8_0_3981));
   NAND2_X1 i_8_0_4154 (.A1(n_8_0_3983), .A2(n_8_0_5850), .ZN(n_8_0_3982));
   OAI21_X1 i_8_0_4155 (.A(n_8_0_6321), .B1(n_8_0_4525), .B2(n_8_0_870), 
      .ZN(n_8_0_3983));
   NOR2_X1 i_8_0_4156 (.A1(n_8_0_4515), .A2(n_8_0_3985), .ZN(n_8_0_3984));
   NOR2_X1 i_8_0_4157 (.A1(n_8_0_5854), .A2(n_8_0_4512), .ZN(n_8_0_3985));
   OAI221_X1 i_8_0_4158 (.A(n_8_0_6606), .B1(n_8_0_5846), .B2(n_8_0_4499), 
      .C1(n_8_0_3987), .C2(n_8_0_869), .ZN(n_8_0_3986));
   INV_X1 i_8_0_4159 (.A(n_8_0_3988), .ZN(n_8_0_3987));
   OAI21_X1 i_8_0_4160 (.A(n_8_0_4587), .B1(n_8_0_4519), .B2(n_8_0_5846), 
      .ZN(n_8_0_3988));
   OAI21_X1 i_8_0_4161 (.A(n_8_0_3990), .B1(n_8_0_4595), .B2(n_8_0_864), 
      .ZN(n_8_0_3989));
   AOI21_X1 i_8_0_4162 (.A(n_8_0_6466), .B1(n_8_0_3991), .B2(n_8_0_5842), 
      .ZN(n_8_0_3990));
   AOI21_X1 i_8_0_4163 (.A(n_8_0_4599), .B1(n_8_0_6469), .B2(n_8_0_864), 
      .ZN(n_8_0_3991));
   OAI221_X1 i_8_0_4164 (.A(n_8_0_6590), .B1(n_8_0_5828), .B2(n_8_0_4555), 
      .C1(n_8_0_3993), .C2(n_8_0_865), .ZN(n_8_0_3992));
   AOI21_X1 i_8_0_4165 (.A(n_8_0_4611), .B1(n_8_0_4565), .B2(n_8_0_5827), 
      .ZN(n_8_0_3993));
   OAI21_X1 i_8_0_4166 (.A(n_8_0_4559), .B1(n_8_0_5455), .B2(n_8_0_5893), 
      .ZN(n_8_0_3994));
   OAI211_X1 i_8_0_4170 (.A(n_8_0_4017), .B(n_8_0_4007), .C1(n_8_0_4008), 
      .C2(n_8_0_863), .ZN(n_8_0_3997));
   INV_X1 i_8_0_4172 (.A(n_8_0_4000), .ZN(n_8_0_3999));
   AOI21_X1 i_8_0_4173 (.A(n_8_0_5865), .B1(n_8_0_6325), .B2(n_8_0_860), 
      .ZN(n_8_0_4000));
   OAI211_X1 i_8_0_4177 (.A(n_8_0_6590), .B(n_8_0_4005), .C1(n_8_0_4555), 
      .C2(n_8_0_5970), .ZN(n_8_0_4004));
   INV_X1 i_8_0_4178 (.A(n_8_0_4006), .ZN(n_8_0_4005));
   AOI211_X1 i_8_0_4179 (.A(n_8_0_857), .B(n_8_0_4558), .C1(n_8_0_4610), 
      .C2(n_8_0_5970), .ZN(n_8_0_4006));
   AOI21_X1 i_8_0_4180 (.A(n_8_0_6250), .B1(n_8_0_5942), .B2(n_8_0_6597), 
      .ZN(n_8_0_4007));
   AOI21_X1 i_8_0_4181 (.A(n_8_0_4515), .B1(n_8_0_4513), .B2(n_8_0_5942), 
      .ZN(n_8_0_4008));
   AOI21_X1 i_8_0_4182 (.A(n_8_0_4010), .B1(n_8_0_5460), .B2(n_8_0_5871), 
      .ZN(n_8_0_4009));
   INV_X1 i_8_0_4183 (.A(n_8_0_4011), .ZN(n_8_0_4010));
   OAI22_X1 i_8_0_4184 (.A1(n_8_0_4058), .A2(n_8_0_4012), .B1(n_8_0_859), 
      .B2(n_8_0_4383), .ZN(n_8_0_4011));
   AND2_X1 i_8_0_4185 (.A1(n_8_0_5871), .A2(n_8_0_7035), .ZN(n_8_0_4012));
   NOR2_X1 i_8_0_4187 (.A1(n_8_0_4015), .A2(n_8_0_6679), .ZN(n_8_0_4014));
   OAI21_X1 i_8_0_4188 (.A(n_8_0_4106), .B1(n_8_0_4573), .B2(n_8_0_858), 
      .ZN(n_8_0_4015));
   OAI221_X1 i_8_0_4189 (.A(n_8_0_6606), .B1(n_8_0_5991), .B2(n_8_0_4499), 
      .C1(n_8_0_4095), .C2(n_8_0_861), .ZN(n_8_0_4016));
   AOI21_X1 i_8_0_4190 (.A(n_8_0_6527), .B1(n_8_0_4019), .B2(n_8_0_4018), 
      .ZN(n_8_0_4017));
   OAI22_X1 i_8_0_4191 (.A1(n_8_0_4579), .A2(n_8_0_862), .B1(n_8_0_5980), 
      .B2(n_8_0_4582), .ZN(n_8_0_4018));
   NAND2_X1 i_8_0_4192 (.A1(n_8_0_862), .A2(n_8_0_5397), .ZN(n_8_0_4019));
   NOR2_X1 i_8_0_4200 (.A1(n_8_0_4027), .A2(n_8_0_6557), .ZN(n_8_0_4026));
   OAI21_X1 i_8_0_4201 (.A(n_8_0_4028), .B1(n_8_0_4542), .B2(n_8_0_851), 
      .ZN(n_8_0_4027));
   OAI21_X1 i_8_0_4202 (.A(n_8_0_5897), .B1(n_8_0_4485), .B2(n_8_0_4029), 
      .ZN(n_8_0_4028));
   NOR3_X1 i_8_0_4203 (.A1(\out_as[4] [6]), .A2(n_8_0_851), .A3(n_8_0_4487), 
      .ZN(n_8_0_4029));
   AOI21_X1 i_8_0_4204 (.A(n_8_0_4031), .B1(n_8_0_5917), .B2(n_8_0_6326), 
      .ZN(n_8_0_4030));
   OAI21_X1 i_8_0_4205 (.A(n_8_0_6577), .B1(n_8_0_4032), .B2(n_8_0_852), 
      .ZN(n_8_0_4031));
   AOI21_X1 i_8_0_4206 (.A(n_8_0_4591), .B1(n_8_0_4593), .B2(n_8_0_5917), 
      .ZN(n_8_0_4032));
   AOI211_X1 i_8_0_4208 (.A(n_8_0_853), .B(n_8_0_4095), .C1(n_8_0_4587), 
      .C2(n_8_0_5906), .ZN(n_8_0_4034));
   AOI21_X1 i_8_0_4210 (.A(n_8_0_4580), .B1(n_8_0_4526), .B2(n_8_0_5902), 
      .ZN(n_8_0_4036));
   OAI221_X1 i_8_0_4212 (.A(n_8_0_6249), .B1(n_8_0_5908), .B2(n_8_0_4454), 
      .C1(n_8_0_4039), .C2(n_8_0_855), .ZN(n_8_0_4038));
   AOI21_X1 i_8_0_4213 (.A(n_8_0_4515), .B1(n_8_0_4513), .B2(n_8_0_5907), 
      .ZN(n_8_0_4039));
   NOR3_X1 i_8_0_4215 (.A1(n_8_0_6516), .A2(n_8_0_4042), .A3(n_8_0_4105), 
      .ZN(n_8_0_4041));
   NOR2_X1 i_8_0_4216 (.A1(n_8_0_4573), .A2(n_8_0_850), .ZN(n_8_0_4042));
   OAI21_X1 i_8_0_4218 (.A(n_8_0_4045), .B1(n_8_0_4611), .B2(n_8_0_5891), 
      .ZN(n_8_0_4044));
   OAI22_X1 i_8_0_4219 (.A1(n_8_0_849), .A2(n_8_0_4558), .B1(n_8_0_4348), 
      .B2(n_8_0_5892), .ZN(n_8_0_4045));
   OAI211_X1 i_8_0_4224 (.A(n_8_0_4070), .B(n_8_0_4073), .C1(n_8_0_4514), 
      .C2(n_8_0_847), .ZN(n_8_0_4049));
   INV_X1 i_8_0_4229 (.A(n_8_0_4055), .ZN(n_8_0_4054));
   OAI221_X1 i_8_0_4230 (.A(n_8_0_6577), .B1(n_8_0_4590), .B2(n_8_0_844), 
      .C1(n_8_0_4592), .C2(n_8_0_5932), .ZN(n_8_0_4055));
   OAI21_X1 i_8_0_4232 (.A(n_8_0_4058), .B1(n_8_0_4540), .B2(n_8_0_843), 
      .ZN(n_8_0_4057));
   NAND2_X1 i_8_0_4233 (.A1(n_8_0_6794), .A2(n_8_0_4486), .ZN(n_8_0_4058));
   NOR2_X1 i_8_0_4234 (.A1(n_8_0_6795), .A2(n_8_0_4487), .ZN(n_8_0_4059));
   NAND2_X1 i_8_0_4235 (.A1(n_8_0_6556), .A2(n_8_0_5927), .ZN(n_8_0_4060));
   NOR2_X1 i_8_0_4236 (.A1(n_8_0_4542), .A2(n_8_0_843), .ZN(n_8_0_4061));
   INV_X1 i_8_0_4237 (.A(n_8_0_4063), .ZN(n_8_0_4062));
   OAI221_X1 i_8_0_4238 (.A(n_8_0_6590), .B1(n_8_0_5936), .B2(n_8_0_4555), 
      .C1(n_8_0_4064), .C2(n_8_0_841), .ZN(n_8_0_4063));
   OAI21_X1 i_8_0_4239 (.A(n_8_0_4559), .B1(n_8_0_4611), .B2(n_8_0_5935), 
      .ZN(n_8_0_4064));
   AOI21_X1 i_8_0_4241 (.A(n_8_0_4588), .B1(n_8_0_4520), .B2(n_8_0_5948), 
      .ZN(n_8_0_4066));
   AND2_X1 i_8_0_4242 (.A1(n_8_0_4069), .A2(n_8_0_4068), .ZN(n_8_0_4067));
   OAI221_X1 i_8_0_4243 (.A(n_8_0_6513), .B1(n_8_0_5957), .B2(n_8_0_4576), 
      .C1(n_8_0_4571), .C2(n_8_0_842), .ZN(n_8_0_4068));
   NAND2_X1 i_8_0_4244 (.A1(n_8_0_842), .A2(n_8_0_6828), .ZN(n_8_0_4069));
   AOI211_X1 i_8_0_4245 (.A(n_8_0_6527), .B(n_8_0_4071), .C1(n_8_0_4580), 
      .C2(n_8_0_6971), .ZN(n_8_0_4070));
   AOI21_X1 i_8_0_4246 (.A(n_8_0_5961), .B1(n_8_0_4072), .B2(n_8_0_6321), 
      .ZN(n_8_0_4071));
   NAND2_X1 i_8_0_4247 (.A1(n_8_0_4526), .A2(n_8_0_6971), .ZN(n_8_0_4072));
   NAND2_X1 i_8_0_4248 (.A1(n_8_0_4074), .A2(n_8_0_5940), .ZN(n_8_0_4073));
   OAI21_X1 i_8_0_4249 (.A(n_8_0_6596), .B1(n_8_0_4512), .B2(n_8_0_847), 
      .ZN(n_8_0_4074));
   OAI211_X1 i_8_0_4254 (.A(n_8_0_4086), .B(n_8_0_4131), .C1(n_8_0_839), 
      .C2(n_8_0_4089), .ZN(n_8_0_4078));
   INV_X1 i_8_0_4258 (.A(n_8_0_4083), .ZN(n_8_0_4082));
   AOI21_X1 i_8_0_4260 (.A(n_8_0_6591), .B1(n_8_0_4556), .B2(n_8_0_5969), 
      .ZN(n_8_0_4084));
   AOI21_X1 i_8_0_4261 (.A(n_8_0_4611), .B1(n_8_0_4565), .B2(n_8_0_5969), 
      .ZN(n_8_0_4085));
   AOI21_X1 i_8_0_4262 (.A(n_8_0_4087), .B1(n_8_0_4088), .B2(n_8_0_5979), 
      .ZN(n_8_0_4086));
   OAI21_X1 i_8_0_4263 (.A(n_8_0_6526), .B1(n_8_0_4579), .B2(n_8_0_838), 
      .ZN(n_8_0_4087));
   OAI21_X1 i_8_0_4264 (.A(n_8_0_6321), .B1(n_8_0_4525), .B2(n_8_0_838), 
      .ZN(n_8_0_4088));
   AOI21_X1 i_8_0_4265 (.A(n_8_0_4128), .B1(n_8_0_4513), .B2(n_8_0_6664), 
      .ZN(n_8_0_4089));
   NAND3_X1 i_8_0_4267 (.A1(\out_bs[3] [5]), .A2(n_8_0_4092), .A3(n_8_0_6005), 
      .ZN(n_8_0_4091));
   AOI21_X1 i_8_0_4268 (.A(\out_bs[3] [6]), .B1(n_8_0_836), .B2(n_8_0_6840), 
      .ZN(n_8_0_4092));
   OAI221_X1 i_8_0_4269 (.A(n_8_0_6606), .B1(n_8_0_6282), .B2(n_8_0_5988), 
      .C1(n_8_0_4094), .C2(n_8_0_837), .ZN(n_8_0_4093));
   AOI21_X1 i_8_0_4270 (.A(n_8_0_4588), .B1(n_8_0_4520), .B2(n_8_0_5989), 
      .ZN(n_8_0_4094));
   AOI21_X1 i_8_0_4271 (.A(n_8_0_4588), .B1(n_8_0_4520), .B2(n_8_0_5990), 
      .ZN(n_8_0_4095));
   OAI21_X1 i_8_0_4273 (.A(n_8_0_6556), .B1(n_8_0_5996), .B2(n_8_0_4098), 
      .ZN(n_8_0_4097));
   AOI21_X1 i_8_0_4274 (.A(n_8_0_4485), .B1(n_8_0_4099), .B2(n_8_0_6911), 
      .ZN(n_8_0_4098));
   NOR2_X1 i_8_0_4275 (.A1(\out_as[4] [6]), .A2(n_8_0_4487), .ZN(n_8_0_4099));
   AOI211_X1 i_8_0_4277 (.A(n_8_0_4107), .B(n_8_0_4102), .C1(n_8_0_4104), 
      .C2(n_8_0_834), .ZN(n_8_0_4101));
   NOR2_X1 i_8_0_4278 (.A1(n_8_0_4103), .A2(n_8_0_6674), .ZN(n_8_0_4102));
   OAI21_X1 i_8_0_4279 (.A(n_8_0_4106), .B1(n_8_0_4573), .B2(n_8_0_834), 
      .ZN(n_8_0_4103));
   NAND2_X1 i_8_0_4280 (.A1(n_8_0_6826), .A2(n_8_0_4109), .ZN(n_8_0_4104));
   NAND2_X1 i_8_0_4281 (.A1(n_8_0_7024), .A2(n_8_0_7022), .ZN(n_8_0_4105));
   NOR2_X1 i_8_0_4282 (.A1(\out_bs[5] [6]), .A2(\out_bs[5] [4]), .ZN(n_8_0_4106));
   NOR2_X1 i_8_0_4283 (.A1(n_8_0_4572), .A2(n_8_0_4108), .ZN(n_8_0_4107));
   AOI21_X1 i_8_0_4284 (.A(n_8_0_4110), .B1(n_8_0_6831), .B2(\out_bs[5] [6]), 
      .ZN(n_8_0_4108));
   NAND2_X1 i_8_0_4285 (.A1(n_8_0_7024), .A2(n_8_0_7023), .ZN(n_8_0_4109));
   NOR2_X1 i_8_0_4286 (.A1(\out_bs[5] [6]), .A2(\out_bs[5] [5]), .ZN(n_8_0_4110));
   AOI21_X1 i_8_0_4287 (.A(n_8_0_6853), .B1(n_8_0_4115), .B2(n_8_0_4111), 
      .ZN(n_132));
   NOR4_X1 i_8_0_4288 (.A1(n_8_0_4123), .A2(n_8_0_4119), .A3(n_8_0_4114), 
      .A4(n_8_0_4112), .ZN(n_8_0_4111));
   NAND3_X1 i_8_0_4289 (.A1(n_8_0_4113), .A2(n_8_0_4131), .A3(n_8_0_4129), 
      .ZN(n_8_0_4112));
   AOI21_X1 i_8_0_4290 (.A(n_8_0_4120), .B1(n_8_0_4128), .B2(n_8_0_6982), 
      .ZN(n_8_0_4113));
   NAND2_X1 i_8_0_4291 (.A1(n_8_0_4117), .A2(n_8_0_4134), .ZN(n_8_0_4114));
   AOI21_X1 i_8_0_4294 (.A(n_8_0_4118), .B1(n_8_0_4556), .B2(\out_bs[6] [4]), 
      .ZN(n_8_0_4117));
   OAI21_X1 i_8_0_4295 (.A(n_8_0_6590), .B1(n_8_0_4457), .B2(n_8_0_819), 
      .ZN(n_8_0_4118));
   OAI211_X1 i_8_0_4296 (.A(n_8_0_6577), .B(n_8_0_4307), .C1(n_8_0_4306), 
      .C2(n_8_0_825), .ZN(n_8_0_4119));
   INV_X1 i_8_0_4297 (.A(n_8_0_4121), .ZN(n_8_0_4120));
   OAI21_X1 i_8_0_4298 (.A(n_8_0_4122), .B1(n_8_0_6827), .B2(n_8_0_6899), 
      .ZN(n_8_0_4121));
   OAI211_X1 i_8_0_4299 (.A(n_8_0_6513), .B(n_8_0_4574), .C1(n_8_0_4571), 
      .C2(n_8_0_821), .ZN(n_8_0_4122));
   OAI221_X1 i_8_0_4300 (.A(n_8_0_6606), .B1(n_8_0_4499), .B2(n_8_0_7058), 
      .C1(n_8_0_4124), .C2(n_8_0_827), .ZN(n_8_0_4123));
   AOI21_X1 i_8_0_4301 (.A(n_8_0_4588), .B1(n_8_0_4520), .B2(\out_bs[2] [4]), 
      .ZN(n_8_0_4124));
   NAND2_X1 i_8_0_4302 (.A1(n_8_0_7066), .A2(n_8_0_4126), .ZN(n_8_0_4125));
   NAND2_X1 i_8_0_4303 (.A1(n_8_0_6774), .A2(n_8_0_4367), .ZN(n_8_0_4126));
   NOR2_X1 i_8_0_4304 (.A1(n_8_0_6775), .A2(n_8_0_4366), .ZN(n_8_0_4127));
   AOI21_X1 i_8_0_4305 (.A(\out_as[0] [6]), .B1(n_8_0_6816), .B2(n_8_0_4602), 
      .ZN(n_8_0_4128));
   AOI21_X1 i_8_0_4306 (.A(n_8_0_4229), .B1(n_8_0_4130), .B2(n_8_0_7078), 
      .ZN(n_8_0_4129));
   AOI21_X1 i_8_0_4307 (.A(n_8_0_829), .B1(n_8_0_6786), .B2(n_8_0_4230), 
      .ZN(n_8_0_4130));
   OR2_X1 i_8_0_4308 (.A1(n_8_0_6811), .A2(n_8_0_4602), .ZN(n_8_0_4131));
   NAND2_X1 i_8_0_4309 (.A1(n_8_0_6810), .A2(n_8_0_4603), .ZN(n_8_0_4132));
   NOR2_X1 i_8_0_4310 (.A1(n_8_0_6811), .A2(n_8_0_4604), .ZN(n_8_0_4133));
   OAI22_X1 i_8_0_4311 (.A1(n_8_0_4135), .A2(n_8_0_6557), .B1(n_8_0_6637), 
      .B2(n_8_0_5459), .ZN(n_8_0_4134));
   OAI21_X1 i_8_0_4312 (.A(n_8_0_4338), .B1(n_8_0_823), .B2(\out_as[4] [6]), 
      .ZN(n_8_0_4135));
   NAND3_X1 i_8_0_4316 (.A1(n_8_0_4139), .A2(n_8_0_4142), .A3(n_8_0_4145), 
      .ZN(n_8_0_4138));
   NAND3_X1 i_8_0_4317 (.A1(n_8_0_4261), .A2(n_8_0_4141), .A3(n_8_0_4140), 
      .ZN(n_8_0_4139));
   OAI211_X1 i_8_0_4318 (.A(n_8_0_811), .B(n_8_0_6606), .C1(n_8_0_6282), 
      .C2(n_8_0_6046), .ZN(n_8_0_4140));
   NAND2_X1 i_8_0_4319 (.A1(n_8_0_6336), .A2(n_8_0_4265), .ZN(n_8_0_4141));
   AOI21_X1 i_8_0_4320 (.A(n_8_0_4143), .B1(n_8_0_4545), .B2(n_8_0_6031), 
      .ZN(n_8_0_4142));
   OAI21_X1 i_8_0_4321 (.A(n_8_0_6556), .B1(n_8_0_4144), .B2(n_8_0_807), 
      .ZN(n_8_0_4143));
   AOI21_X1 i_8_0_4322 (.A(n_8_0_4543), .B1(n_8_0_4539), .B2(n_8_0_6031), 
      .ZN(n_8_0_4144));
   AOI21_X1 i_8_0_4323 (.A(n_8_0_4146), .B1(n_8_0_4308), .B2(n_8_0_5086), 
      .ZN(n_8_0_4145));
   OAI21_X1 i_8_0_4324 (.A(n_8_0_6577), .B1(n_8_0_4147), .B2(n_8_0_809), 
      .ZN(n_8_0_4146));
   AOI21_X1 i_8_0_4325 (.A(n_8_0_4591), .B1(n_8_0_4414), .B2(n_8_0_5086), 
      .ZN(n_8_0_4147));
   OAI221_X1 i_8_0_4326 (.A(n_8_0_6249), .B1(n_8_0_6054), .B2(n_8_0_4454), 
      .C1(n_8_0_4149), .C2(n_8_0_815), .ZN(n_8_0_4148));
   AOI21_X1 i_8_0_4327 (.A(n_8_0_4515), .B1(n_8_0_4513), .B2(n_8_0_6053), 
      .ZN(n_8_0_4149));
   OAI21_X1 i_8_0_4328 (.A(n_8_0_4151), .B1(n_8_0_4152), .B2(n_8_0_805), 
      .ZN(n_8_0_4150));
   AOI21_X1 i_8_0_4329 (.A(n_8_0_6514), .B1(n_8_0_6059), .B2(n_8_0_4553), 
      .ZN(n_8_0_4151));
   AOI21_X1 i_8_0_4330 (.A(n_8_0_4572), .B1(n_8_0_4550), .B2(n_8_0_6059), 
      .ZN(n_8_0_4152));
   OAI211_X1 i_8_0_4331 (.A(n_8_0_6526), .B(n_8_0_4154), .C1(n_8_0_4579), 
      .C2(n_8_0_813), .ZN(n_8_0_4153));
   OAI21_X1 i_8_0_4332 (.A(n_8_0_6050), .B1(n_8_0_4229), .B2(n_8_0_4155), 
      .ZN(n_8_0_4154));
   NOR3_X1 i_8_0_4333 (.A1(n_8_0_4230), .A2(n_8_0_813), .A3(\out_as[1] [6]), 
      .ZN(n_8_0_4155));
   OAI211_X1 i_8_0_4335 (.A(n_8_0_6590), .B(n_8_0_4158), .C1(n_8_0_4610), 
      .C2(n_8_0_803), .ZN(n_8_0_4157));
   INV_X1 i_8_0_4336 (.A(n_8_0_4159), .ZN(n_8_0_4158));
   AOI211_X1 i_8_0_4337 (.A(n_8_0_6036), .B(n_8_0_4255), .C1(n_8_0_803), 
      .C2(n_8_0_6755), .ZN(n_8_0_4159));
   NAND3_X1 i_8_0_4344 (.A1(n_8_0_4169), .A2(n_8_0_4166), .A3(n_8_0_4172), 
      .ZN(n_8_0_4165));
   AOI21_X1 i_8_0_4345 (.A(n_8_0_4167), .B1(n_8_0_4168), .B2(n_8_0_6074), 
      .ZN(n_8_0_4166));
   OAI21_X1 i_8_0_4346 (.A(n_8_0_6526), .B1(n_8_0_4579), .B2(n_8_0_797), 
      .ZN(n_8_0_4167));
   OAI21_X1 i_8_0_4347 (.A(n_8_0_6321), .B1(n_8_0_4525), .B2(n_8_0_797), 
      .ZN(n_8_0_4168));
   AOI21_X1 i_8_0_4348 (.A(n_8_0_4170), .B1(n_8_0_4171), .B2(n_8_0_6069), 
      .ZN(n_8_0_4169));
   OAI21_X1 i_8_0_4349 (.A(n_8_0_6606), .B1(n_8_0_4587), .B2(n_8_0_795), 
      .ZN(n_8_0_4170));
   OAI21_X1 i_8_0_4350 (.A(n_8_0_6282), .B1(n_8_0_4519), .B2(n_8_0_795), 
      .ZN(n_8_0_4171));
   NAND2_X1 i_8_0_4351 (.A1(n_8_0_6082), .A2(n_8_0_4173), .ZN(n_8_0_4172));
   OAI21_X1 i_8_0_4352 (.A(n_8_0_4454), .B1(n_8_0_4512), .B2(n_8_0_799), 
      .ZN(n_8_0_4173));
   OAI21_X1 i_8_0_4353 (.A(n_8_0_6249), .B1(n_8_0_4514), .B2(n_8_0_799), 
      .ZN(n_8_0_4174));
   OAI21_X1 i_8_0_4354 (.A(n_8_0_4176), .B1(n_8_0_4571), .B2(n_8_0_789), 
      .ZN(n_8_0_4175));
   AOI21_X1 i_8_0_4355 (.A(n_8_0_6514), .B1(n_8_0_4177), .B2(n_8_0_6097), 
      .ZN(n_8_0_4176));
   AOI21_X1 i_8_0_4356 (.A(n_8_0_4574), .B1(n_8_0_6828), .B2(n_8_0_789), 
      .ZN(n_8_0_4177));
   OAI21_X1 i_8_0_4358 (.A(n_8_0_6556), .B1(n_8_0_4180), .B2(n_8_0_791), 
      .ZN(n_8_0_4179));
   AOI21_X1 i_8_0_4359 (.A(n_8_0_4543), .B1(n_8_0_4539), .B2(n_8_0_6092), 
      .ZN(n_8_0_4180));
   OAI21_X1 i_8_0_4361 (.A(n_8_0_6577), .B1(n_8_0_4183), .B2(n_8_0_793), 
      .ZN(n_8_0_4182));
   AOI21_X1 i_8_0_4362 (.A(n_8_0_4591), .B1(n_8_0_4414), .B2(n_8_0_5116), 
      .ZN(n_8_0_4183));
   NAND2_X1 i_8_0_4365 (.A1(n_8_0_4531), .A2(n_8_0_6080), .ZN(n_8_0_4186));
   OAI21_X1 i_8_0_4367 (.A(n_8_0_6590), .B1(n_8_0_4255), .B2(n_8_0_4189), 
      .ZN(n_8_0_4188));
   OAI21_X1 i_8_0_4368 (.A(n_8_0_6088), .B1(n_8_0_6754), .B2(n_8_0_6878), 
      .ZN(n_8_0_4189));
   NAND4_X1 i_8_0_4371 (.A1(n_8_0_4211), .A2(n_8_0_4196), .A3(n_8_0_4193), 
      .A4(n_8_0_4192), .ZN(n_8_0_4191));
   AOI21_X1 i_8_0_4372 (.A(n_8_0_4203), .B1(n_8_0_4202), .B2(n_8_0_6140), 
      .ZN(n_8_0_4192));
   AOI21_X1 i_8_0_4373 (.A(n_8_0_4194), .B1(n_8_0_4195), .B2(n_8_0_6131), 
      .ZN(n_8_0_4193));
   OAI21_X1 i_8_0_4374 (.A(n_8_0_6606), .B1(n_8_0_4587), .B2(n_8_0_779), 
      .ZN(n_8_0_4194));
   OAI21_X1 i_8_0_4375 (.A(n_8_0_6282), .B1(n_8_0_4519), .B2(n_8_0_779), 
      .ZN(n_8_0_4195));
   AOI21_X1 i_8_0_4376 (.A(n_8_0_4200), .B1(n_8_0_4201), .B2(n_8_0_6127), 
      .ZN(n_8_0_4196));
   NAND2_X1 i_8_0_4377 (.A1(n_8_0_7078), .A2(n_8_0_4198), .ZN(n_8_0_4197));
   NAND2_X1 i_8_0_4378 (.A1(n_8_0_5397), .A2(n_8_0_4325), .ZN(n_8_0_4198));
   NOR2_X1 i_8_0_4379 (.A1(n_8_0_5396), .A2(n_8_0_4324), .ZN(n_8_0_4199));
   OAI21_X1 i_8_0_4380 (.A(n_8_0_6526), .B1(n_8_0_4579), .B2(n_8_0_781), 
      .ZN(n_8_0_4200));
   OAI21_X1 i_8_0_4381 (.A(n_8_0_6321), .B1(n_8_0_4525), .B2(n_8_0_781), 
      .ZN(n_8_0_4201));
   OAI21_X1 i_8_0_4382 (.A(n_8_0_4454), .B1(n_8_0_4512), .B2(n_8_0_783), 
      .ZN(n_8_0_4202));
   OAI21_X1 i_8_0_4383 (.A(n_8_0_6249), .B1(n_8_0_4514), .B2(n_8_0_783), 
      .ZN(n_8_0_4203));
   OAI211_X1 i_8_0_4384 (.A(n_8_0_6513), .B(n_8_0_4205), .C1(n_8_0_4571), 
      .C2(n_8_0_773), .ZN(n_8_0_4204));
   OAI211_X1 i_8_0_4385 (.A(n_8_0_4575), .B(n_8_0_6136), .C1(n_8_0_6827), 
      .C2(n_8_0_6898), .ZN(n_8_0_4205));
   INV_X1 i_8_0_4388 (.A(n_8_0_4209), .ZN(n_8_0_4208));
   OAI221_X1 i_8_0_4389 (.A(n_8_0_6577), .B1(n_8_0_4210), .B2(n_8_0_777), 
      .C1(n_8_0_4307), .C2(n_8_0_6109), .ZN(n_8_0_4209));
   AOI21_X1 i_8_0_4390 (.A(n_8_0_4591), .B1(n_8_0_4414), .B2(n_8_0_6108), 
      .ZN(n_8_0_4210));
   OAI21_X1 i_8_0_4392 (.A(n_8_0_6590), .B1(n_8_0_4348), .B2(n_8_0_6123), 
      .ZN(n_8_0_4212));
   AOI21_X1 i_8_0_4393 (.A(n_8_0_771), .B1(n_8_0_4610), .B2(n_8_0_6123), 
      .ZN(n_8_0_4213));
   INV_X1 i_8_0_4394 (.A(n_8_0_4215), .ZN(n_8_0_4214));
   AOI21_X1 i_8_0_4395 (.A(n_8_0_4216), .B1(n_8_0_4545), .B2(n_8_0_6113), 
      .ZN(n_8_0_4215));
   OAI21_X1 i_8_0_4396 (.A(n_8_0_6556), .B1(n_8_0_4217), .B2(n_8_0_775), 
      .ZN(n_8_0_4216));
   AOI21_X1 i_8_0_4397 (.A(n_8_0_4543), .B1(n_8_0_4539), .B2(n_8_0_6113), 
      .ZN(n_8_0_4217));
   AOI21_X1 i_8_0_4398 (.A(n_8_0_6853), .B1(n_8_0_4233), .B2(n_8_0_4218), 
      .ZN(n_133));
   NOR4_X1 i_8_0_4399 (.A1(n_8_0_4241), .A2(n_8_0_4236), .A3(n_8_0_4219), 
      .A4(n_8_0_6250), .ZN(n_8_0_4218));
   OAI211_X1 i_8_0_4400 (.A(n_8_0_4220), .B(n_8_0_4221), .C1(n_8_0_4454), 
      .C2(n_8_0_6174), .ZN(n_8_0_4219));
   NOR4_X1 i_8_0_4401 (.A1(n_8_0_4243), .A2(n_8_0_4239), .A3(n_8_0_4226), 
      .A4(n_8_0_4223), .ZN(n_8_0_4220));
   NAND2_X1 i_8_0_4402 (.A1(n_8_0_6981), .A2(n_8_0_4222), .ZN(n_8_0_4221));
   OAI21_X1 i_8_0_4403 (.A(n_8_0_4514), .B1(n_8_0_4512), .B2(n_8_0_6174), 
      .ZN(n_8_0_4222));
   OAI21_X1 i_8_0_4404 (.A(n_8_0_4224), .B1(n_8_0_4571), .B2(n_8_0_757), 
      .ZN(n_8_0_4223));
   NOR2_X1 i_8_0_4405 (.A1(n_8_0_6514), .A2(n_8_0_4225), .ZN(n_8_0_4224));
   AOI211_X1 i_8_0_4406 (.A(n_8_0_4574), .B(n_8_0_6166), .C1(n_8_0_6828), 
      .C2(n_8_0_757), .ZN(n_8_0_4225));
   OAI211_X1 i_8_0_4407 (.A(n_8_0_6526), .B(n_8_0_4227), .C1(n_8_0_4579), 
      .C2(n_8_0_765), .ZN(n_8_0_4226));
   OAI22_X1 i_8_0_4408 (.A1(\out_bs[1] [3]), .A2(\out_bs[1] [2]), .B1(n_8_0_4229), 
      .B2(n_8_0_4228), .ZN(n_8_0_4227));
   NOR3_X1 i_8_0_4409 (.A1(n_8_0_4230), .A2(n_8_0_765), .A3(\out_as[1] [6]), 
      .ZN(n_8_0_4228));
   NOR2_X1 i_8_0_4410 (.A1(n_8_0_6782), .A2(n_8_0_4230), .ZN(n_8_0_4229));
   AOI21_X1 i_8_0_4411 (.A(\out_bs[1] [6]), .B1(\out_bs[1] [5]), .B2(
      \out_bs[1] [4]), .ZN(n_8_0_4230));
   NAND2_X1 i_8_0_4412 (.A1(n_8_0_6781), .A2(n_8_0_4324), .ZN(n_8_0_4231));
   NAND2_X1 i_8_0_4413 (.A1(n_8_0_6526), .A2(n_8_0_6321), .ZN(n_8_0_4232));
   NOR2_X1 i_8_0_4414 (.A1(n_8_0_4235), .A2(n_8_0_4234), .ZN(n_8_0_4233));
   OAI21_X1 i_8_0_4415 (.A(n_8_0_6465), .B1(n_8_0_6467), .B2(n_8_0_6157), 
      .ZN(n_8_0_4234));
   AOI211_X1 i_8_0_4416 (.A(n_8_0_753), .B(n_8_0_4503), .C1(n_8_0_4595), 
      .C2(n_8_0_6157), .ZN(n_8_0_4235));
   OAI211_X1 i_8_0_4417 (.A(n_8_0_6590), .B(n_8_0_4237), .C1(n_8_0_4555), 
      .C2(n_8_0_6293), .ZN(n_8_0_4236));
   INV_X1 i_8_0_4418 (.A(n_8_0_4238), .ZN(n_8_0_4237));
   AOI211_X1 i_8_0_4419 (.A(n_8_0_755), .B(n_8_0_4558), .C1(n_8_0_4610), 
      .C2(n_8_0_6293), .ZN(n_8_0_4238));
   OAI221_X1 i_8_0_4420 (.A(n_8_0_6577), .B1(n_8_0_4240), .B2(n_8_0_761), 
      .C1(n_8_0_4307), .C2(n_8_0_6161), .ZN(n_8_0_4239));
   AOI21_X1 i_8_0_4421 (.A(n_8_0_4591), .B1(n_8_0_4414), .B2(n_8_0_6160), 
      .ZN(n_8_0_4240));
   OAI221_X1 i_8_0_4422 (.A(n_8_0_6556), .B1(n_8_0_6171), .B2(n_8_0_4338), 
      .C1(n_8_0_4242), .C2(n_8_0_759), .ZN(n_8_0_4241));
   AOI21_X1 i_8_0_4423 (.A(n_8_0_4543), .B1(n_8_0_4539), .B2(n_8_0_6170), 
      .ZN(n_8_0_4242));
   AOI21_X1 i_8_0_4424 (.A(n_8_0_4244), .B1(n_8_0_4265), .B2(n_8_0_7056), 
      .ZN(n_8_0_4243));
   OAI21_X1 i_8_0_4425 (.A(n_8_0_4261), .B1(n_8_0_4245), .B2(n_8_0_6607), 
      .ZN(n_8_0_4244));
   OAI21_X1 i_8_0_4426 (.A(n_8_0_763), .B1(n_8_0_6282), .B2(n_8_0_6151), 
      .ZN(n_8_0_4245));
   INV_X1 i_8_0_4430 (.A(n_8_0_4249), .ZN(n_8_0_4248));
   AOI211_X1 i_8_0_4431 (.A(n_8_0_743), .B(n_8_0_4383), .C1(n_8_0_4542), 
      .C2(n_8_0_6190), .ZN(n_8_0_4249));
   AOI21_X1 i_8_0_4433 (.A(n_8_0_4572), .B1(n_8_0_4550), .B2(n_8_0_6210), 
      .ZN(n_8_0_4251));
   INV_X1 i_8_0_4435 (.A(n_8_0_4254), .ZN(n_8_0_4253));
   AOI211_X1 i_8_0_4436 (.A(n_8_0_6198), .B(n_8_0_4255), .C1(n_8_0_739), 
      .C2(n_8_0_6755), .ZN(n_8_0_4254));
   OAI21_X1 i_8_0_4437 (.A(\out_bs[6] [4]), .B1(n_8_0_4565), .B2(n_8_0_4556), 
      .ZN(n_8_0_4255));
   NAND2_X1 i_8_0_4441 (.A1(n_8_0_6201), .A2(n_8_0_4531), .ZN(n_8_0_4259));
   NOR2_X1 i_8_0_4443 (.A1(n_8_0_4585), .A2(n_8_0_4262), .ZN(n_8_0_4261));
   AOI21_X1 i_8_0_4444 (.A(n_8_0_4586), .B1(\out_bs[2] [4]), .B2(\out_bs[2] [5]), 
      .ZN(n_8_0_4262));
   OAI211_X1 i_8_0_4445 (.A(n_8_0_747), .B(n_8_0_6606), .C1(n_8_0_6282), 
      .C2(n_8_0_6182), .ZN(n_8_0_4263));
   NAND2_X1 i_8_0_4446 (.A1(n_8_0_6537), .A2(n_8_0_4265), .ZN(n_8_0_4264));
   NOR2_X1 i_8_0_4447 (.A1(n_8_0_4586), .A2(\out_bs[2] [3]), .ZN(n_8_0_4265));
   OAI21_X1 i_8_0_4449 (.A(n_8_0_6249), .B1(n_8_0_4514), .B2(n_8_0_751), 
      .ZN(n_8_0_4267));
   OAI21_X1 i_8_0_4450 (.A(n_8_0_4454), .B1(n_8_0_4512), .B2(n_8_0_751), 
      .ZN(n_8_0_4268));
   OAI221_X1 i_8_0_4451 (.A(n_8_0_6526), .B1(n_8_0_4270), .B2(n_8_0_6206), 
      .C1(n_8_0_749), .C2(n_8_0_4579), .ZN(n_8_0_4269));
   INV_X1 i_8_0_4452 (.A(n_8_0_4271), .ZN(n_8_0_4270));
   OAI21_X1 i_8_0_4453 (.A(n_8_0_6321), .B1(n_8_0_4525), .B2(n_8_0_749), 
      .ZN(n_8_0_4271));
   OAI221_X1 i_8_0_4455 (.A(n_8_0_6577), .B1(n_8_0_4274), .B2(n_8_0_745), 
      .C1(n_8_0_4307), .C2(n_8_0_6216), .ZN(n_8_0_4273));
   AOI21_X1 i_8_0_4456 (.A(n_8_0_4591), .B1(n_8_0_4414), .B2(n_8_0_6215), 
      .ZN(n_8_0_4274));
   NAND2_X1 i_8_0_4461 (.A1(n_8_0_4282), .A2(n_8_0_4279), .ZN(n_8_0_4278));
   AOI21_X1 i_8_0_4462 (.A(n_8_0_4280), .B1(n_8_0_4553), .B2(n_8_0_6300), 
      .ZN(n_8_0_4279));
   OAI21_X1 i_8_0_4463 (.A(n_8_0_6513), .B1(n_8_0_4281), .B2(n_8_0_725), 
      .ZN(n_8_0_4280));
   AOI21_X1 i_8_0_4464 (.A(n_8_0_4572), .B1(n_8_0_4575), .B2(n_8_0_6300), 
      .ZN(n_8_0_4281));
   AOI21_X1 i_8_0_4465 (.A(n_8_0_4283), .B1(n_8_0_4284), .B2(n_8_0_6271), 
      .ZN(n_8_0_4282));
   OAI21_X1 i_8_0_4466 (.A(n_8_0_6526), .B1(n_8_0_4579), .B2(n_8_0_733), 
      .ZN(n_8_0_4283));
   OAI21_X1 i_8_0_4467 (.A(n_8_0_6321), .B1(n_8_0_4525), .B2(n_8_0_733), 
      .ZN(n_8_0_4284));
   OAI21_X1 i_8_0_4468 (.A(n_8_0_4454), .B1(n_8_0_4512), .B2(n_8_0_735), 
      .ZN(n_8_0_4285));
   OAI211_X1 i_8_0_4469 (.A(n_8_0_4287), .B(n_8_0_6249), .C1(n_8_0_735), 
      .C2(n_8_0_4514), .ZN(n_8_0_4286));
   AOI21_X1 i_8_0_4470 (.A(n_8_0_4288), .B1(n_8_0_4289), .B2(n_8_0_6288), 
      .ZN(n_8_0_4287));
   OAI21_X1 i_8_0_4471 (.A(n_8_0_6606), .B1(n_8_0_4587), .B2(n_8_0_731), 
      .ZN(n_8_0_4288));
   OAI21_X1 i_8_0_4472 (.A(n_8_0_6282), .B1(n_8_0_4519), .B2(n_8_0_731), 
      .ZN(n_8_0_4289));
   AOI21_X1 i_8_0_4476 (.A(n_8_0_4591), .B1(n_8_0_4414), .B2(n_8_0_6217), 
      .ZN(n_8_0_4293));
   AOI21_X1 i_8_0_4478 (.A(n_8_0_4296), .B1(n_8_0_4545), .B2(n_8_0_6244), 
      .ZN(n_8_0_4295));
   OAI21_X1 i_8_0_4479 (.A(n_8_0_6556), .B1(n_8_0_4297), .B2(n_8_0_727), 
      .ZN(n_8_0_4296));
   AOI21_X1 i_8_0_4480 (.A(n_8_0_4543), .B1(n_8_0_4539), .B2(n_8_0_6244), 
      .ZN(n_8_0_4297));
   AOI211_X1 i_8_0_4481 (.A(n_8_0_6591), .B(n_8_0_4299), .C1(n_8_0_4349), 
      .C2(n_8_0_6225), .ZN(n_8_0_4298));
   AOI21_X1 i_8_0_4482 (.A(n_8_0_723), .B1(n_8_0_4420), .B2(n_8_0_4300), 
      .ZN(n_8_0_4299));
   NAND3_X1 i_8_0_4483 (.A1(\out_bs[6] [4]), .A2(n_8_0_6744), .A3(n_8_0_4565), 
      .ZN(n_8_0_4300));
   INV_X1 i_8_0_4488 (.A(n_8_0_4305), .ZN(n_8_0_4304));
   AOI211_X1 i_8_0_4489 (.A(n_8_0_713), .B(n_8_0_4306), .C1(n_8_0_4590), 
      .C2(n_8_0_5698), .ZN(n_8_0_4305));
   NOR2_X1 i_8_0_4490 (.A1(n_8_0_4591), .A2(n_8_0_4414), .ZN(n_8_0_4306));
   NAND2_X1 i_8_0_4491 (.A1(\out_bs[3] [4]), .A2(n_8_0_6326), .ZN(n_8_0_4307));
   NOR2_X1 i_8_0_4492 (.A1(n_8_0_7045), .A2(n_8_0_6325), .ZN(n_8_0_4308));
   NAND2_X1 i_8_0_4493 (.A1(\out_bs[3] [4]), .A2(n_8_0_6838), .ZN(n_8_0_4309));
   NOR2_X1 i_8_0_4494 (.A1(n_8_0_7045), .A2(n_8_0_6837), .ZN(n_8_0_4310));
   OAI21_X1 i_8_0_4495 (.A(\out_bs[3] [4]), .B1(\out_bs[3] [3]), .B2(n_8_0_6650), 
      .ZN(n_8_0_4311));
   AOI211_X1 i_8_0_4497 (.A(n_8_0_707), .B(n_8_0_4558), .C1(n_8_0_4610), 
      .C2(n_8_0_6292), .ZN(n_8_0_4313));
   OAI21_X1 i_8_0_4499 (.A(n_8_0_4316), .B1(n_8_0_4317), .B2(n_8_0_709), 
      .ZN(n_8_0_4315));
   AOI21_X1 i_8_0_4500 (.A(n_8_0_6514), .B1(n_8_0_6299), .B2(n_8_0_4553), 
      .ZN(n_8_0_4316));
   AOI21_X1 i_8_0_4501 (.A(n_8_0_4572), .B1(n_8_0_4575), .B2(n_8_0_6299), 
      .ZN(n_8_0_4317));
   OAI211_X1 i_8_0_4503 (.A(n_8_0_4320), .B(n_8_0_6249), .C1(n_8_0_6261), 
      .C2(n_8_0_4454), .ZN(n_8_0_4319));
   AOI22_X1 i_8_0_4504 (.A1(n_8_0_6781), .A2(n_8_0_4322), .B1(n_8_0_4321), 
      .B2(n_8_0_7078), .ZN(n_8_0_4320));
   AOI21_X1 i_8_0_4505 (.A(n_8_0_717), .B1(n_8_0_6786), .B2(n_8_0_4323), 
      .ZN(n_8_0_4321));
   INV_X1 i_8_0_4506 (.A(n_8_0_4323), .ZN(n_8_0_4322));
   OAI21_X1 i_8_0_4507 (.A(n_8_0_4324), .B1(n_8_0_6268), .B2(\out_bs[1] [6]), 
      .ZN(n_8_0_4323));
   NAND2_X1 i_8_0_4508 (.A1(n_8_0_7072), .A2(n_8_0_7071), .ZN(n_8_0_4324));
   NOR2_X1 i_8_0_4509 (.A1(\out_bs[1] [6]), .A2(\out_bs[1] [5]), .ZN(n_8_0_4325));
   OAI21_X1 i_8_0_4510 (.A(n_8_0_4514), .B1(n_8_0_4512), .B2(n_8_0_6261), 
      .ZN(n_8_0_4326));
   INV_X1 i_8_0_4511 (.A(n_8_0_4328), .ZN(n_8_0_4327));
   AOI21_X1 i_8_0_4513 (.A(n_8_0_4543), .B1(n_8_0_4541), .B2(n_8_0_6275), 
      .ZN(n_8_0_4329));
   AOI21_X1 i_8_0_4515 (.A(n_8_0_4588), .B1(n_8_0_4520), .B2(n_8_0_6285), 
      .ZN(n_8_0_4331));
   AOI21_X1 i_8_0_4519 (.A(n_8_0_6853), .B1(n_8_0_4340), .B2(n_8_0_4335), 
      .ZN(n_134));
   NOR3_X1 i_8_0_4520 (.A1(n_8_0_4339), .A2(n_8_0_4337), .A3(n_8_0_4336), 
      .ZN(n_8_0_4335));
   OAI221_X1 i_8_0_4521 (.A(n_8_0_6465), .B1(n_8_0_6467), .B2(n_8_0_6997), 
      .C1(n_8_0_682), .C2(n_8_0_4530), .ZN(n_8_0_4336));
   OAI221_X1 i_8_0_4522 (.A(n_8_0_6556), .B1(n_8_0_4484), .B2(n_8_0_6632), 
      .C1(n_8_0_4538), .C2(n_8_0_691), .ZN(n_8_0_4337));
   NAND2_X1 i_8_0_4523 (.A1(n_8_0_6799), .A2(n_8_0_6637), .ZN(n_8_0_4338));
   OAI221_X1 i_8_0_4524 (.A(n_8_0_6577), .B1(n_8_0_6325), .B2(n_8_0_6647), 
      .C1(n_8_0_4413), .C2(n_8_0_694), .ZN(n_8_0_4339));
   NOR4_X1 i_8_0_4525 (.A1(n_8_0_4350), .A2(n_8_0_4345), .A3(n_8_0_4342), 
      .A4(n_8_0_4341), .ZN(n_8_0_4340));
   OAI21_X1 i_8_0_4526 (.A(n_8_0_6249), .B1(n_8_0_4454), .B2(n_8_0_6662), 
      .ZN(n_8_0_4341));
   AND2_X1 i_8_0_4527 (.A1(n_8_0_4344), .A2(n_8_0_4343), .ZN(n_8_0_4342));
   NAND3_X1 i_8_0_4528 (.A1(n_8_0_6526), .A2(n_8_0_4581), .A3(n_8_0_4579), 
      .ZN(n_8_0_4343));
   OAI211_X1 i_8_0_4529 (.A(n_8_0_6526), .B(n_8_0_700), .C1(n_8_0_4581), 
      .C2(n_8_0_5397), .ZN(n_8_0_4344));
   OAI221_X1 i_8_0_4530 (.A(n_8_0_6590), .B1(n_8_0_4348), .B2(n_8_0_6750), 
      .C1(n_8_0_4420), .C2(n_8_0_685), .ZN(n_8_0_4345));
   NAND2_X1 i_8_0_4531 (.A1(n_8_0_6590), .A2(n_8_0_4348), .ZN(n_8_0_4346));
   NAND2_X1 i_8_0_4532 (.A1(n_8_0_6754), .A2(n_8_0_4562), .ZN(n_8_0_4347));
   NAND2_X1 i_8_0_4533 (.A1(\out_bs[6] [5]), .A2(n_8_0_6757), .ZN(n_8_0_4348));
   NOR2_X1 i_8_0_4534 (.A1(n_8_0_7011), .A2(n_8_0_6756), .ZN(n_8_0_4349));
   OAI211_X1 i_8_0_4535 (.A(n_8_0_4353), .B(n_8_0_4351), .C1(n_8_0_703), 
      .C2(n_8_0_4511), .ZN(n_8_0_4350));
   INV_X1 i_8_0_4536 (.A(n_8_0_4352), .ZN(n_8_0_4351));
   OAI221_X1 i_8_0_4537 (.A(n_8_0_6513), .B1(n_8_0_4552), .B2(n_8_0_7021), 
      .C1(n_8_0_4549), .C2(n_8_0_688), .ZN(n_8_0_4352));
   AOI21_X1 i_8_0_4538 (.A(n_8_0_4354), .B1(n_8_0_6283), .B2(n_8_0_6709), 
      .ZN(n_8_0_4353));
   OAI21_X1 i_8_0_4539 (.A(n_8_0_6606), .B1(n_8_0_4369), .B2(n_8_0_697), 
      .ZN(n_8_0_4354));
   AOI211_X1 i_8_0_4543 (.A(n_8_0_4359), .B(n_8_0_4358), .C1(n_8_0_6343), 
      .C2(n_8_0_4362), .ZN(n_8_0_4357));
   OAI21_X1 i_8_0_4544 (.A(n_8_0_6249), .B1(n_8_0_4514), .B2(n_8_0_679), 
      .ZN(n_8_0_4358));
   OAI211_X1 i_8_0_4545 (.A(n_8_0_6526), .B(n_8_0_4360), .C1(n_8_0_4579), 
      .C2(n_8_0_676), .ZN(n_8_0_4359));
   NAND2_X1 i_8_0_4546 (.A1(n_8_0_4361), .A2(n_8_0_6340), .ZN(n_8_0_4360));
   OAI21_X1 i_8_0_4547 (.A(n_8_0_6321), .B1(n_8_0_4525), .B2(n_8_0_676), 
      .ZN(n_8_0_4361));
   OAI21_X1 i_8_0_4548 (.A(n_8_0_6596), .B1(n_8_0_4512), .B2(n_8_0_679), 
      .ZN(n_8_0_4362));
   NAND2_X1 i_8_0_4550 (.A1(n_8_0_6773), .A2(n_8_0_4366), .ZN(n_8_0_4364));
   NOR2_X1 i_8_0_4551 (.A1(n_8_0_6772), .A2(n_8_0_4367), .ZN(n_8_0_4365));
   NAND2_X1 i_8_0_4552 (.A1(n_8_0_7060), .A2(n_8_0_7059), .ZN(n_8_0_4366));
   NOR2_X1 i_8_0_4553 (.A1(\out_bs[2] [6]), .A2(\out_bs[2] [5]), .ZN(n_8_0_4367));
   AOI21_X1 i_8_0_4554 (.A(n_8_0_4588), .B1(n_8_0_4520), .B2(n_8_0_6334), 
      .ZN(n_8_0_4368));
   AOI21_X1 i_8_0_4555 (.A(n_8_0_4588), .B1(n_8_0_4520), .B2(n_8_0_6709), 
      .ZN(n_8_0_4369));
   AOI211_X1 i_8_0_4559 (.A(n_8_0_6591), .B(n_8_0_4374), .C1(n_8_0_4556), 
      .C2(n_8_0_6367), .ZN(n_8_0_4373));
   AOI211_X1 i_8_0_4560 (.A(n_8_0_661), .B(n_8_0_4558), .C1(n_8_0_4610), 
      .C2(n_8_0_6366), .ZN(n_8_0_4374));
   AOI21_X1 i_8_0_4562 (.A(n_8_0_6514), .B1(n_8_0_4377), .B2(n_8_0_6373), 
      .ZN(n_8_0_4376));
   OAI21_X1 i_8_0_4563 (.A(n_8_0_4378), .B1(n_8_0_4551), .B2(n_8_0_664), 
      .ZN(n_8_0_4377));
   NAND2_X1 i_8_0_4564 (.A1(\out_bs[5] [5]), .A2(n_8_0_6825), .ZN(n_8_0_4378));
   OAI211_X1 i_8_0_4566 (.A(n_8_0_6556), .B(n_8_0_4381), .C1(n_8_0_4544), 
      .C2(n_8_0_6350), .ZN(n_8_0_4380));
   OAI21_X1 i_8_0_4567 (.A(n_8_0_4382), .B1(n_8_0_4543), .B2(n_8_0_6349), 
      .ZN(n_8_0_4381));
   NOR2_X1 i_8_0_4568 (.A1(n_8_0_667), .A2(n_8_0_4383), .ZN(n_8_0_4382));
   NAND2_X1 i_8_0_4569 (.A1(n_8_0_7040), .A2(n_8_0_4384), .ZN(n_8_0_4383));
   NAND2_X1 i_8_0_4570 (.A1(n_8_0_6801), .A2(n_8_0_4487), .ZN(n_8_0_4384));
   NOR2_X1 i_8_0_4571 (.A1(n_8_0_6800), .A2(n_8_0_4486), .ZN(n_8_0_4385));
   OAI221_X1 i_8_0_4572 (.A(n_8_0_6577), .B1(n_8_0_6355), .B2(n_8_0_6325), 
      .C1(n_8_0_4387), .C2(n_8_0_670), .ZN(n_8_0_4386));
   AOI21_X1 i_8_0_4573 (.A(n_8_0_4591), .B1(n_8_0_4593), .B2(n_8_0_6356), 
      .ZN(n_8_0_4387));
   NAND3_X1 i_8_0_4576 (.A1(n_8_0_4411), .A2(n_8_0_4393), .A3(n_8_0_4390), 
      .ZN(n_8_0_4389));
   AOI21_X1 i_8_0_4577 (.A(n_8_0_4391), .B1(n_8_0_4392), .B2(n_8_0_6398), 
      .ZN(n_8_0_4390));
   OAI21_X1 i_8_0_4578 (.A(n_8_0_6606), .B1(n_8_0_4587), .B2(n_8_0_649), 
      .ZN(n_8_0_4391));
   OAI21_X1 i_8_0_4579 (.A(n_8_0_6282), .B1(n_8_0_4519), .B2(n_8_0_649), 
      .ZN(n_8_0_4392));
   OAI21_X1 i_8_0_4580 (.A(n_8_0_4394), .B1(n_8_0_4396), .B2(n_8_0_6794), 
      .ZN(n_8_0_4393));
   INV_X1 i_8_0_4581 (.A(n_8_0_4395), .ZN(n_8_0_4394));
   AOI221_X1 i_8_0_4582 (.A(\out_bs[4] [6]), .B1(\out_bs[4] [5]), .B2(n_8_0_6380), 
      .C1(n_8_0_6800), .C2(n_8_0_4396), .ZN(n_8_0_4395));
   NOR2_X1 i_8_0_4583 (.A1(\out_as[4] [6]), .A2(n_8_0_643), .ZN(n_8_0_4396));
   AOI211_X1 i_8_0_4584 (.A(n_8_0_655), .B(n_8_0_4511), .C1(n_8_0_4514), 
      .C2(n_8_0_6421), .ZN(n_8_0_4397));
   OR4_X1 i_8_0_4585 (.A1(n_8_0_4401), .A2(n_8_0_4399), .A3(n_8_0_6419), 
      .A4(n_8_0_6250), .ZN(n_8_0_4398));
   OAI221_X1 i_8_0_4586 (.A(n_8_0_6526), .B1(n_8_0_6392), .B2(n_8_0_6321), 
      .C1(n_8_0_4400), .C2(n_8_0_652), .ZN(n_8_0_4399));
   AOI21_X1 i_8_0_4587 (.A(n_8_0_4580), .B1(n_8_0_4526), .B2(n_8_0_6393), 
      .ZN(n_8_0_4400));
   OAI21_X1 i_8_0_4588 (.A(n_8_0_4402), .B1(n_8_0_4403), .B2(n_8_0_640), 
      .ZN(n_8_0_4401));
   AOI21_X1 i_8_0_4589 (.A(n_8_0_6514), .B1(n_8_0_6409), .B2(n_8_0_4553), 
      .ZN(n_8_0_4402));
   AOI21_X1 i_8_0_4590 (.A(n_8_0_4572), .B1(n_8_0_4550), .B2(n_8_0_6409), 
      .ZN(n_8_0_4403));
   OAI211_X1 i_8_0_4592 (.A(n_8_0_6590), .B(n_8_0_4407), .C1(n_8_0_4406), 
      .C2(n_8_0_637), .ZN(n_8_0_4405));
   OAI21_X1 i_8_0_4593 (.A(n_8_0_4559), .B1(n_8_0_4611), .B2(n_8_0_6385), 
      .ZN(n_8_0_4406));
   NAND2_X1 i_8_0_4594 (.A1(n_8_0_6385), .A2(n_8_0_4556), .ZN(n_8_0_4407));
   AOI211_X1 i_8_0_4598 (.A(n_8_0_6578), .B(n_8_0_4412), .C1(n_8_0_6326), 
      .C2(n_8_0_6412), .ZN(n_8_0_4411));
   AOI211_X1 i_8_0_4599 (.A(n_8_0_646), .B(n_8_0_4413), .C1(n_8_0_4590), 
      .C2(n_8_0_6414), .ZN(n_8_0_4412));
   AOI21_X1 i_8_0_4600 (.A(n_8_0_4591), .B1(n_8_0_4414), .B2(\out_bs[3] [3]), 
      .ZN(n_8_0_4413));
   NOR3_X1 i_8_0_4601 (.A1(n_8_0_7046), .A2(n_8_0_7045), .A3(\out_as[3] [6]), 
      .ZN(n_8_0_4414));
   AOI21_X1 i_8_0_4602 (.A(n_8_0_6853), .B1(n_8_0_4427), .B2(n_8_0_4415), 
      .ZN(n_135));
   NOR3_X1 i_8_0_4603 (.A1(n_8_0_4437), .A2(n_8_0_4421), .A3(n_8_0_4416), 
      .ZN(n_8_0_4415));
   NAND4_X1 i_8_0_4604 (.A1(n_8_0_4418), .A2(n_8_0_4440), .A3(n_8_0_4434), 
      .A4(n_8_0_4417), .ZN(n_8_0_4416));
   AOI211_X1 i_8_0_4605 (.A(n_8_0_6250), .B(n_8_0_4443), .C1(n_8_0_6597), 
      .C2(n_8_0_6439), .ZN(n_8_0_4417));
   AOI211_X1 i_8_0_4606 (.A(n_8_0_6591), .B(n_8_0_4419), .C1(n_8_0_4556), 
      .C2(n_8_0_6479), .ZN(n_8_0_4418));
   AOI211_X1 i_8_0_4607 (.A(n_8_0_613), .B(n_8_0_4420), .C1(n_8_0_4610), 
      .C2(n_8_0_6481), .ZN(n_8_0_4419));
   AOI21_X1 i_8_0_4608 (.A(n_8_0_4611), .B1(n_8_0_4565), .B2(n_8_0_6751), 
      .ZN(n_8_0_4420));
   OAI211_X1 i_8_0_4609 (.A(n_8_0_6465), .B(n_8_0_4425), .C1(n_8_0_6473), 
      .C2(n_8_0_6469), .ZN(n_8_0_4421));
   OAI21_X1 i_8_0_4613 (.A(n_8_0_6864), .B1(n_8_0_4596), .B2(n_8_0_4426), 
      .ZN(n_8_0_4425));
   NOR3_X1 i_8_0_4614 (.A1(n_8_0_6473), .A2(\out_as[7] [6]), .A3(n_8_0_6999), 
      .ZN(n_8_0_4426));
   NOR2_X1 i_8_0_4615 (.A1(n_8_0_4431), .A2(n_8_0_4428), .ZN(n_8_0_4427));
   OAI211_X1 i_8_0_4616 (.A(n_8_0_6577), .B(n_8_0_4429), .C1(n_8_0_4590), 
      .C2(n_8_0_622), .ZN(n_8_0_4428));
   NAND4_X1 i_8_0_4617 (.A1(n_8_0_4430), .A2(n_8_0_6427), .A3(\out_bs[3] [4]), 
      .A4(\out_bs[3] [5]), .ZN(n_8_0_4429));
   OAI21_X1 i_8_0_4618 (.A(n_8_0_6837), .B1(n_8_0_622), .B2(\out_bs[3] [6]), 
      .ZN(n_8_0_4430));
   INV_X1 i_8_0_4619 (.A(n_8_0_4432), .ZN(n_8_0_4431));
   AOI221_X1 i_8_0_4620 (.A(n_8_0_6557), .B1(n_8_0_4433), .B2(n_8_0_6907), 
      .C1(n_8_0_4545), .C2(n_8_0_6434), .ZN(n_8_0_4432));
   OAI21_X1 i_8_0_4621 (.A(n_8_0_4542), .B1(n_8_0_4540), .B2(n_8_0_6433), 
      .ZN(n_8_0_4433));
   AOI21_X1 i_8_0_4622 (.A(n_8_0_4435), .B1(n_8_0_4553), .B2(n_8_0_6460), 
      .ZN(n_8_0_4434));
   OAI21_X1 i_8_0_4623 (.A(n_8_0_6513), .B1(n_8_0_4436), .B2(n_8_0_616), 
      .ZN(n_8_0_4435));
   AOI21_X1 i_8_0_4624 (.A(n_8_0_4572), .B1(n_8_0_4550), .B2(n_8_0_6460), 
      .ZN(n_8_0_4436));
   OAI21_X1 i_8_0_4625 (.A(n_8_0_4438), .B1(n_8_0_4587), .B2(n_8_0_625), 
      .ZN(n_8_0_4437));
   AOI21_X1 i_8_0_4626 (.A(n_8_0_6607), .B1(n_8_0_6451), .B2(n_8_0_4439), 
      .ZN(n_8_0_4438));
   OAI21_X1 i_8_0_4627 (.A(n_8_0_4499), .B1(n_8_0_4519), .B2(n_8_0_625), 
      .ZN(n_8_0_4439));
   OAI21_X1 i_8_0_4628 (.A(n_8_0_4441), .B1(n_8_0_5396), .B2(n_8_0_6964), 
      .ZN(n_8_0_4440));
   OAI21_X1 i_8_0_4629 (.A(n_8_0_4442), .B1(n_8_0_4581), .B2(n_8_0_6448), 
      .ZN(n_8_0_4441));
   OAI22_X1 i_8_0_4630 (.A1(n_8_0_6527), .A2(n_8_0_4580), .B1(\out_as[1] [6]), 
      .B2(n_8_0_6964), .ZN(n_8_0_4442));
   AOI211_X1 i_8_0_4631 (.A(n_8_0_631), .B(n_8_0_4511), .C1(n_8_0_4514), 
      .C2(n_8_0_6442), .ZN(n_8_0_4443));
   AOI21_X1 i_8_0_4634 (.A(n_8_0_4446), .B1(n_8_0_6828), .B2(n_8_0_587), 
      .ZN(n_8_0_4445));
   INV_X1 i_8_0_4635 (.A(n_8_0_4447), .ZN(n_8_0_4446));
   OAI221_X1 i_8_0_4636 (.A(n_8_0_6513), .B1(n_8_0_4574), .B2(n_8_0_6678), 
      .C1(n_8_0_4571), .C2(n_8_0_587), .ZN(n_8_0_4447));
   OAI21_X1 i_8_0_4637 (.A(n_8_0_4449), .B1(n_8_0_4544), .B2(n_8_0_6641), 
      .ZN(n_8_0_4448));
   AOI21_X1 i_8_0_4638 (.A(n_8_0_6557), .B1(n_8_0_4451), .B2(n_8_0_4450), 
      .ZN(n_8_0_4449));
   NOR2_X1 i_8_0_4639 (.A1(\out_as[4] [6]), .A2(n_8_0_591), .ZN(n_8_0_4450));
   OAI21_X1 i_8_0_4640 (.A(n_8_0_5460), .B1(n_8_0_6638), .B2(n_8_0_6641), 
      .ZN(n_8_0_4451));
   AND3_X1 i_8_0_4641 (.A1(n_8_0_4453), .A2(n_8_0_6663), .A3(\out_bs[0] [2]), 
      .ZN(n_8_0_4452));
   OAI21_X1 i_8_0_4642 (.A(n_8_0_4454), .B1(n_8_0_4512), .B2(n_8_0_607), 
      .ZN(n_8_0_4453));
   NAND2_X1 i_8_0_4643 (.A1(\out_bs[0] [5]), .A2(n_8_0_6814), .ZN(n_8_0_4454));
   OAI211_X1 i_8_0_4644 (.A(n_8_0_6590), .B(n_8_0_4458), .C1(n_8_0_4456), 
      .C2(n_8_0_583), .ZN(n_8_0_4455));
   OAI21_X1 i_8_0_4645 (.A(n_8_0_4559), .B1(n_8_0_4611), .B2(n_8_0_6749), 
      .ZN(n_8_0_4456));
   AOI21_X1 i_8_0_4646 (.A(n_8_0_4611), .B1(n_8_0_4565), .B2(\out_bs[6] [4]), 
      .ZN(n_8_0_4457));
   NAND2_X1 i_8_0_4647 (.A1(n_8_0_6749), .A2(n_8_0_4556), .ZN(n_8_0_4458));
   OAI22_X1 i_8_0_4650 (.A1(n_8_0_4462), .A2(\out_bs[2] [6]), .B1(n_8_0_6773), 
      .B2(n_8_0_4464), .ZN(n_8_0_4461));
   INV_X1 i_8_0_4651 (.A(n_8_0_4463), .ZN(n_8_0_4462));
   AOI22_X1 i_8_0_4652 (.A1(n_8_0_6775), .A2(n_8_0_4464), .B1(n_8_0_6707), 
      .B2(\out_bs[2] [5]), .ZN(n_8_0_4463));
   NOR2_X1 i_8_0_4653 (.A1(\out_as[2] [6]), .A2(n_8_0_599), .ZN(n_8_0_4464));
   INV_X1 i_8_0_4655 (.A(n_8_0_4467), .ZN(n_8_0_4466));
   OAI21_X1 i_8_0_4656 (.A(n_8_0_4579), .B1(n_8_0_4525), .B2(n_8_0_6689), 
      .ZN(n_8_0_4467));
   NOR2_X1 i_8_0_4661 (.A1(n_8_0_4593), .A2(n_8_0_4591), .ZN(n_8_0_4472));
   AOI21_X1 i_8_0_4662 (.A(n_8_0_4591), .B1(n_8_0_4593), .B2(n_8_0_5468), 
      .ZN(n_8_0_4473));
   NOR4_X1 i_8_0_4667 (.A1(n_8_0_4488), .A2(n_8_0_6250), .A3(n_8_0_4491), 
      .A4(n_8_0_4478), .ZN(n_8_0_4477));
   OAI211_X1 i_8_0_4668 (.A(n_8_0_6526), .B(n_8_0_4479), .C1(n_8_0_4579), 
      .C2(n_8_0_571), .ZN(n_8_0_4478));
   INV_X1 i_8_0_4669 (.A(n_8_0_4480), .ZN(n_8_0_4479));
   AOI211_X1 i_8_0_4670 (.A(n_8_0_6532), .B(n_8_0_4581), .C1(n_8_0_5397), 
      .C2(n_8_0_571), .ZN(n_8_0_4480));
   AOI21_X1 i_8_0_4671 (.A(n_8_0_4482), .B1(n_8_0_4483), .B2(n_8_0_6558), 
      .ZN(n_8_0_4481));
   OAI21_X1 i_8_0_4672 (.A(n_8_0_6556), .B1(n_8_0_4542), .B2(n_8_0_559), 
      .ZN(n_8_0_4482));
   OAI21_X1 i_8_0_4673 (.A(n_8_0_4484), .B1(n_8_0_4540), .B2(n_8_0_559), 
      .ZN(n_8_0_4483));
   NAND2_X1 i_8_0_4674 (.A1(n_8_0_6799), .A2(n_8_0_4486), .ZN(n_8_0_4484));
   NOR2_X1 i_8_0_4675 (.A1(n_8_0_6798), .A2(n_8_0_4487), .ZN(n_8_0_4485));
   NAND2_X1 i_8_0_4676 (.A1(n_8_0_7035), .A2(n_8_0_7034), .ZN(n_8_0_4486));
   NOR2_X1 i_8_0_4677 (.A1(\out_bs[4] [6]), .A2(\out_bs[4] [5]), .ZN(n_8_0_4487));
   OAI21_X1 i_8_0_4678 (.A(n_8_0_4489), .B1(n_8_0_4490), .B2(n_8_0_555), 
      .ZN(n_8_0_4488));
   AOI21_X1 i_8_0_4679 (.A(n_8_0_6514), .B1(n_8_0_4553), .B2(n_8_0_6516), 
      .ZN(n_8_0_4489));
   AOI21_X1 i_8_0_4680 (.A(n_8_0_4572), .B1(n_8_0_4550), .B2(n_8_0_6516), 
      .ZN(n_8_0_4490));
   OAI211_X1 i_8_0_4681 (.A(n_8_0_6577), .B(n_8_0_4492), .C1(n_8_0_4590), 
      .C2(n_8_0_563), .ZN(n_8_0_4491));
   INV_X1 i_8_0_4682 (.A(n_8_0_4493), .ZN(n_8_0_4492));
   AOI211_X1 i_8_0_4683 (.A(n_8_0_4494), .B(n_8_0_4592), .C1(n_8_0_6325), 
      .C2(n_8_0_563), .ZN(n_8_0_4493));
   NAND2_X1 i_8_0_4684 (.A1(n_8_0_6565), .A2(n_8_0_6648), .ZN(n_8_0_4494));
   AOI21_X1 i_8_0_4685 (.A(n_8_0_4496), .B1(n_8_0_4497), .B2(n_8_0_6535), 
      .ZN(n_8_0_4495));
   OAI21_X1 i_8_0_4686 (.A(n_8_0_6606), .B1(n_8_0_4587), .B2(n_8_0_567), 
      .ZN(n_8_0_4496));
   OAI21_X1 i_8_0_4687 (.A(n_8_0_4499), .B1(n_8_0_4519), .B2(n_8_0_567), 
      .ZN(n_8_0_4497));
   INV_X1 i_8_0_4688 (.A(n_8_0_4499), .ZN(n_8_0_4498));
   NAND3_X1 i_8_0_4689 (.A1(n_8_0_7060), .A2(n_8_0_6775), .A3(\out_bs[2] [5]), 
      .ZN(n_8_0_4499));
   OAI21_X1 i_8_0_4695 (.A(n_8_0_6590), .B1(n_8_0_4506), .B2(n_8_0_551), 
      .ZN(n_8_0_4505));
   AOI21_X1 i_8_0_4696 (.A(n_8_0_4611), .B1(n_8_0_4565), .B2(n_8_0_6549), 
      .ZN(n_8_0_4506));
   AOI21_X1 i_8_0_4697 (.A(n_8_0_6853), .B1(n_8_0_4527), .B2(n_8_0_4507), 
      .ZN(n_136));
   AND4_X1 i_8_0_4698 (.A1(n_8_0_4554), .A2(n_8_0_4536), .A3(n_8_0_4516), 
      .A4(n_8_0_4508), .ZN(n_8_0_4507));
   NOR4_X1 i_8_0_4699 (.A1(n_8_0_4546), .A2(n_8_0_4521), .A3(n_8_0_4510), 
      .A4(n_8_0_4509), .ZN(n_8_0_4508));
   OAI211_X1 i_8_0_4700 (.A(n_8_0_4533), .B(n_8_0_6249), .C1(n_8_0_6593), 
      .C2(n_8_0_6596), .ZN(n_8_0_4509));
   AOI211_X1 i_8_0_4701 (.A(n_8_0_543), .B(n_8_0_4511), .C1(n_8_0_4514), 
      .C2(n_8_0_6667), .ZN(n_8_0_4510));
   AOI21_X1 i_8_0_4702 (.A(n_8_0_4515), .B1(n_8_0_4513), .B2(n_8_0_6663), 
      .ZN(n_8_0_4511));
   NAND2_X1 i_8_0_4703 (.A1(n_8_0_7089), .A2(\out_bs[0] [5]), .ZN(n_8_0_4512));
   NOR2_X1 i_8_0_4704 (.A1(n_8_0_7084), .A2(\out_as[0] [6]), .ZN(n_8_0_4513));
   NOR2_X1 i_8_0_4706 (.A1(\out_as[0] [6]), .A2(n_8_0_5274), .ZN(n_8_0_4515));
   AOI21_X1 i_8_0_4707 (.A(n_8_0_4517), .B1(n_8_0_4518), .B2(n_8_0_6611), 
      .ZN(n_8_0_4516));
   OAI21_X1 i_8_0_4708 (.A(n_8_0_6606), .B1(n_8_0_4587), .B2(n_8_0_533), 
      .ZN(n_8_0_4517));
   OAI21_X1 i_8_0_4709 (.A(n_8_0_6282), .B1(n_8_0_4519), .B2(n_8_0_533), 
      .ZN(n_8_0_4518));
   NAND2_X1 i_8_0_4710 (.A1(n_8_0_7066), .A2(\out_bs[2] [5]), .ZN(n_8_0_4519));
   NOR2_X1 i_8_0_4711 (.A1(n_8_0_7059), .A2(\out_as[2] [6]), .ZN(n_8_0_4520));
   OAI21_X1 i_8_0_4712 (.A(n_8_0_4522), .B1(n_8_0_4524), .B2(n_8_0_6321), 
      .ZN(n_8_0_4521));
   AOI21_X1 i_8_0_4713 (.A(n_8_0_6527), .B1(n_8_0_4523), .B2(n_8_0_6962), 
      .ZN(n_8_0_4522));
   OAI21_X1 i_8_0_4714 (.A(n_8_0_4579), .B1(n_8_0_4525), .B2(n_8_0_4524), 
      .ZN(n_8_0_4523));
   NAND2_X1 i_8_0_4715 (.A1(n_8_0_6700), .A2(n_8_0_6696), .ZN(n_8_0_4524));
   NAND2_X1 i_8_0_4716 (.A1(n_8_0_7078), .A2(\out_bs[1] [5]), .ZN(n_8_0_4525));
   NOR2_X1 i_8_0_4717 (.A1(n_8_0_7071), .A2(\out_as[1] [6]), .ZN(n_8_0_4526));
   NOR3_X1 i_8_0_4718 (.A1(n_8_0_6466), .A2(n_8_0_4529), .A3(n_8_0_4528), 
      .ZN(n_8_0_4527));
   NOR3_X1 i_8_0_4719 (.A1(n_8_0_6724), .A2(n_8_0_6721), .A3(n_8_0_6469), 
      .ZN(n_8_0_4528));
   AOI211_X1 i_8_0_4720 (.A(n_8_0_508), .B(n_8_0_4530), .C1(n_8_0_4595), 
      .C2(n_8_0_6724), .ZN(n_8_0_4529));
   AOI21_X1 i_8_0_4721 (.A(n_8_0_4596), .B1(n_8_0_4531), .B2(\out_bs[7] [3]), 
      .ZN(n_8_0_4530));
   AOI21_X1 i_8_0_4724 (.A(n_8_0_6578), .B1(n_8_0_4535), .B2(n_8_0_4534), 
      .ZN(n_8_0_4533));
   OAI22_X1 i_8_0_4725 (.A1(n_8_0_6579), .A2(n_8_0_4592), .B1(n_8_0_4590), 
      .B2(n_8_0_528), .ZN(n_8_0_4534));
   NAND2_X1 i_8_0_4726 (.A1(n_8_0_6325), .A2(n_8_0_528), .ZN(n_8_0_4535));
   AOI211_X1 i_8_0_4727 (.A(n_8_0_6557), .B(n_8_0_4537), .C1(n_8_0_4545), 
      .C2(n_8_0_6640), .ZN(n_8_0_4536));
   AOI211_X1 i_8_0_4728 (.A(n_8_0_523), .B(n_8_0_4538), .C1(n_8_0_4542), 
      .C2(n_8_0_6642), .ZN(n_8_0_4537));
   AOI21_X1 i_8_0_4729 (.A(n_8_0_4543), .B1(n_8_0_4539), .B2(\out_bs[4] [3]), 
      .ZN(n_8_0_4538));
   NOR2_X1 i_8_0_4730 (.A1(n_8_0_6638), .A2(\out_as[4] [6]), .ZN(n_8_0_4539));
   NAND2_X1 i_8_0_4731 (.A1(n_8_0_7040), .A2(\out_bs[4] [5]), .ZN(n_8_0_4540));
   NOR2_X1 i_8_0_4732 (.A1(n_8_0_7034), .A2(\out_as[4] [6]), .ZN(n_8_0_4541));
   NAND2_X1 i_8_0_4733 (.A1(n_8_0_7040), .A2(n_8_0_5459), .ZN(n_8_0_4542));
   NOR2_X1 i_8_0_4734 (.A1(\out_as[4] [6]), .A2(n_8_0_5460), .ZN(n_8_0_4543));
   INV_X1 i_8_0_4735 (.A(n_8_0_4545), .ZN(n_8_0_4544));
   NOR2_X1 i_8_0_4736 (.A1(n_8_0_6795), .A2(n_8_0_6638), .ZN(n_8_0_4545));
   NAND2_X1 i_8_0_4737 (.A1(n_8_0_6513), .A2(n_8_0_4547), .ZN(n_8_0_4546));
   OAI21_X1 i_8_0_4738 (.A(n_8_0_4548), .B1(n_8_0_4572), .B2(n_8_0_6682), 
      .ZN(n_8_0_4547));
   OAI22_X1 i_8_0_4739 (.A1(n_8_0_518), .A2(n_8_0_4549), .B1(n_8_0_4552), 
      .B2(n_8_0_6675), .ZN(n_8_0_4548));
   AOI21_X1 i_8_0_4740 (.A(n_8_0_4572), .B1(n_8_0_4550), .B2(\out_bs[5] [3]), 
      .ZN(n_8_0_4549));
   NOR2_X1 i_8_0_4741 (.A1(n_8_0_7022), .A2(n_8_0_4551), .ZN(n_8_0_4550));
   NAND2_X1 i_8_0_4742 (.A1(n_8_0_7030), .A2(\out_bs[5] [5]), .ZN(n_8_0_4551));
   NAND2_X1 i_8_0_4743 (.A1(n_8_0_6827), .A2(n_8_0_4575), .ZN(n_8_0_4552));
   NOR2_X1 i_8_0_4744 (.A1(n_8_0_6828), .A2(n_8_0_4574), .ZN(n_8_0_4553));
   AOI211_X1 i_8_0_4745 (.A(n_8_0_6591), .B(n_8_0_4557), .C1(n_8_0_4556), 
      .C2(n_8_0_6742), .ZN(n_8_0_4554));
   NAND2_X1 i_8_0_4746 (.A1(n_8_0_6754), .A2(\out_bs[6] [5]), .ZN(n_8_0_4555));
   NOR2_X1 i_8_0_4747 (.A1(n_8_0_6755), .A2(n_8_0_7011), .ZN(n_8_0_4556));
   AOI211_X1 i_8_0_4748 (.A(n_8_0_513), .B(n_8_0_4558), .C1(n_8_0_4610), 
      .C2(n_8_0_6741), .ZN(n_8_0_4557));
   NAND2_X1 i_8_0_4749 (.A1(n_8_0_7018), .A2(n_8_0_4560), .ZN(n_8_0_4558));
   NOR2_X1 i_8_0_4750 (.A1(\out_as[6] [6]), .A2(n_8_0_4561), .ZN(n_8_0_4559));
   NAND2_X1 i_8_0_4751 (.A1(n_8_0_6761), .A2(n_8_0_4563), .ZN(n_8_0_4560));
   NOR2_X1 i_8_0_4752 (.A1(n_8_0_6760), .A2(n_8_0_4562), .ZN(n_8_0_4561));
   NAND2_X1 i_8_0_4753 (.A1(n_8_0_7012), .A2(n_8_0_7011), .ZN(n_8_0_4562));
   NOR2_X1 i_8_0_4754 (.A1(\out_bs[6] [6]), .A2(\out_bs[6] [5]), .ZN(n_8_0_4563));
   NAND2_X1 i_8_0_4755 (.A1(n_8_0_7018), .A2(\out_bs[6] [5]), .ZN(n_8_0_4564));
   NOR2_X1 i_8_0_4756 (.A1(n_8_0_7011), .A2(\out_as[6] [6]), .ZN(n_8_0_4565));
   OAI221_X1 i_8_0_4762 (.A(n_8_0_4571), .B1(n_8_0_4574), .B2(n_8_0_6673), 
      .C1(n_8_0_7024), .C2(n_8_0_6831), .ZN(n_8_0_4570));
   OAI21_X1 i_8_0_4763 (.A(n_8_0_7030), .B1(n_8_0_6830), .B2(\out_bs[5] [6]), 
      .ZN(n_8_0_4571));
   NOR2_X1 i_8_0_4764 (.A1(\out_as[5] [6]), .A2(n_8_0_5302), .ZN(n_8_0_4572));
   NAND2_X1 i_8_0_4765 (.A1(n_8_0_7030), .A2(n_8_0_6830), .ZN(n_8_0_4573));
   NAND2_X1 i_8_0_4766 (.A1(\out_bs[5] [4]), .A2(n_8_0_4577), .ZN(n_8_0_4574));
   NOR2_X1 i_8_0_4767 (.A1(n_8_0_7022), .A2(n_8_0_4576), .ZN(n_8_0_4575));
   INV_X1 i_8_0_4768 (.A(n_8_0_4577), .ZN(n_8_0_4576));
   NOR2_X1 i_8_0_4769 (.A1(n_8_0_7023), .A2(\out_bs[5] [6]), .ZN(n_8_0_4577));
   OAI211_X1 i_8_0_4770 (.A(n_8_0_6526), .B(n_8_0_4579), .C1(n_8_0_4581), 
      .C2(n_8_0_6697), .ZN(n_8_0_4578));
   NAND2_X1 i_8_0_4771 (.A1(n_8_0_7078), .A2(n_8_0_5394), .ZN(n_8_0_4579));
   NOR2_X1 i_8_0_4772 (.A1(\out_as[1] [6]), .A2(n_8_0_5395), .ZN(n_8_0_4580));
   NAND3_X1 i_8_0_4773 (.A1(n_8_0_6696), .A2(n_8_0_7072), .A3(\out_bs[1] [5]), 
      .ZN(n_8_0_4581));
   NAND2_X1 i_8_0_4774 (.A1(n_8_0_7072), .A2(\out_bs[1] [5]), .ZN(n_8_0_4582));
   NOR2_X1 i_8_0_4776 (.A1(n_8_0_4585), .A2(n_8_0_6703), .ZN(n_8_0_4584));
   NOR2_X1 i_8_0_4777 (.A1(n_8_0_7066), .A2(n_8_0_6775), .ZN(n_8_0_4585));
   NAND2_X1 i_8_0_4778 (.A1(n_8_0_6606), .A2(n_8_0_4587), .ZN(n_8_0_4586));
   NAND2_X1 i_8_0_4779 (.A1(n_8_0_7066), .A2(n_8_0_5427), .ZN(n_8_0_4587));
   NOR2_X1 i_8_0_4780 (.A1(\out_as[2] [6]), .A2(n_8_0_5428), .ZN(n_8_0_4588));
   NAND2_X1 i_8_0_4782 (.A1(n_8_0_7053), .A2(n_8_0_4621), .ZN(n_8_0_4590));
   NOR2_X1 i_8_0_4783 (.A1(\out_as[3] [6]), .A2(n_8_0_4622), .ZN(n_8_0_4591));
   AOI21_X1 i_8_0_4784 (.A(n_8_0_4593), .B1(n_8_0_6839), .B2(\out_bs[3] [5]), 
      .ZN(n_8_0_4592));
   NOR2_X1 i_8_0_4785 (.A1(n_8_0_7046), .A2(\out_as[3] [6]), .ZN(n_8_0_4593));
   AOI22_X1 i_8_0_4793 (.A1(n_8_0_4606), .A2(n_8_0_4605), .B1(\out_as[0] [6]), 
      .B2(n_8_0_6816), .ZN(n_8_0_4601));
   AOI21_X1 i_8_0_4794 (.A(\out_bs[0] [6]), .B1(\out_bs[0] [5]), .B2(
      \out_bs[0] [4]), .ZN(n_8_0_4602));
   NAND2_X1 i_8_0_4795 (.A1(n_8_0_7085), .A2(n_8_0_7084), .ZN(n_8_0_4603));
   NOR2_X1 i_8_0_4796 (.A1(\out_bs[0] [6]), .A2(\out_bs[0] [5]), .ZN(n_8_0_4604));
   AOI21_X1 i_8_0_4797 (.A(\out_bs[0] [6]), .B1(n_8_0_6817), .B2(n_8_0_7089), 
      .ZN(n_8_0_4605));
   NAND3_X1 i_8_0_4798 (.A1(\out_bs[0] [5]), .A2(n_8_0_6666), .A3(n_8_0_6663), 
      .ZN(n_8_0_4606));
   AOI21_X1 i_8_0_4799 (.A(n_8_0_4608), .B1(n_8_0_6801), .B2(\out_as[4] [6]), 
      .ZN(n_8_0_4607));
   AOI22_X1 i_8_0_4800 (.A1(n_8_0_6809), .A2(n_8_0_5459), .B1(n_8_0_6628), 
      .B2(\out_bs[4] [5]), .ZN(n_8_0_4608));
   OAI211_X1 i_8_0_4801 (.A(n_8_0_4612), .B(n_8_0_4610), .C1(n_8_0_7012), 
      .C2(n_8_0_6761), .ZN(n_8_0_4609));
   NAND2_X1 i_8_0_4802 (.A1(n_8_0_7018), .A2(n_8_0_5455), .ZN(n_8_0_4610));
   NOR2_X1 i_8_0_4803 (.A1(\out_as[6] [6]), .A2(n_8_0_5456), .ZN(n_8_0_4611));
   OAI211_X1 i_8_0_4804 (.A(\out_bs[6] [5]), .B(n_8_0_5454), .C1(n_8_0_6760), 
      .C2(n_8_0_7018), .ZN(n_8_0_4612));
   AOI21_X1 i_8_0_4813 (.A(n_8_0_189), .B1(n_8_0_4622), .B2(n_8_0_7053), 
      .ZN(n_8_0_4620));
   INV_X1 i_8_0_4814 (.A(n_8_0_4622), .ZN(n_8_0_4621));
   NOR2_X1 i_8_0_4815 (.A1(\out_bs[3] [6]), .A2(n_8_0_6846), .ZN(n_8_0_4622));
   AOI21_X1 i_8_0_4819 (.A(n_8_0_6853), .B1(n_8_0_4626), .B2(n_8_0_4647), 
      .ZN(n_137));
   NOR3_X1 i_8_0_4820 (.A1(n_8_0_4644), .A2(n_8_0_4633), .A3(n_8_0_4627), 
      .ZN(n_8_0_4626));
   NAND4_X1 i_8_0_4821 (.A1(n_8_0_4628), .A2(n_8_0_4639), .A3(n_8_0_4650), 
      .A4(n_8_0_4629), .ZN(n_8_0_4627));
   AOI21_X1 i_8_0_4822 (.A(n_8_0_4636), .B1(n_8_0_4642), .B2(n_8_0_4643), 
      .ZN(n_8_0_4628));
   AOI21_X1 i_8_0_4823 (.A(n_8_0_4631), .B1(n_8_0_6233), .B2(n_8_0_4630), 
      .ZN(n_8_0_4629));
   NAND2_X1 i_8_0_4824 (.A1(n_8_0_4632), .A2(n_8_0_442), .ZN(n_8_0_4630));
   NOR2_X1 i_8_0_4825 (.A1(n_8_0_4632), .A2(n_8_0_442), .ZN(n_8_0_4631));
   OAI21_X1 i_8_0_4826 (.A(\out_bs[7] [6]), .B1(n_8_0_6042), .B2(n_8_0_5056), 
      .ZN(n_8_0_4632));
   OAI21_X1 i_8_0_4827 (.A(n_8_0_4634), .B1(n_8_0_6772), .B2(n_8_0_127), 
      .ZN(n_8_0_4633));
   OAI211_X1 i_8_0_4828 (.A(n_8_0_4635), .B(\out_bs[2] [6]), .C1(n_8_0_6335), 
      .C2(n_8_0_4834), .ZN(n_8_0_4634));
   NAND2_X1 i_8_0_4829 (.A1(n_8_0_6772), .A2(n_8_0_127), .ZN(n_8_0_4635));
   OAI21_X1 i_8_0_4830 (.A(n_8_0_4637), .B1(n_8_0_6824), .B2(n_8_0_316), 
      .ZN(n_8_0_4636));
   OAI21_X1 i_8_0_4831 (.A(n_8_0_4638), .B1(n_8_0_5519), .B2(\out_bs[5] [5]), 
      .ZN(n_8_0_4637));
   AOI21_X1 i_8_0_4832 (.A(n_8_0_7024), .B1(n_8_0_6619), .B2(n_8_0_316), 
      .ZN(n_8_0_4638));
   OAI21_X1 i_8_0_4833 (.A(n_8_0_4640), .B1(n_8_0_5262), .B2(n_8_0_5525), 
      .ZN(n_8_0_4639));
   AOI21_X1 i_8_0_4834 (.A(n_8_0_5395), .B1(n_8_0_4641), .B2(n_8_0_64), .ZN(
      n_8_0_4640));
   OAI21_X1 i_8_0_4835 (.A(n_8_0_6527), .B1(n_8_0_5525), .B2(\out_bs[1] [5]), 
      .ZN(n_8_0_4641));
   OAI21_X1 i_8_0_4836 (.A(n_8_0_6249), .B1(n_8_0_5274), .B2(n_8_0_4), .ZN(
      n_8_0_4642));
   OAI211_X1 i_8_0_4837 (.A(n_8_0_7084), .B(n_8_0_5506), .C1(n_8_0_6811), 
      .C2(n_8_0_4), .ZN(n_8_0_4643));
   OAI21_X1 i_8_0_4838 (.A(n_8_0_4645), .B1(n_8_0_6837), .B2(n_8_0_190), 
      .ZN(n_8_0_4644));
   OAI211_X1 i_8_0_4839 (.A(n_8_0_4646), .B(\out_bs[3] [6]), .C1(\out_bs[3] [5]), 
      .C2(n_8_0_5500), .ZN(n_8_0_4645));
   NAND2_X1 i_8_0_4840 (.A1(n_8_0_6844), .A2(n_8_0_190), .ZN(n_8_0_4646));
   OAI21_X1 i_8_0_4841 (.A(n_8_0_4648), .B1(n_8_0_4649), .B2(n_8_0_6031), 
      .ZN(n_8_0_4647));
   OAI21_X1 i_8_0_4842 (.A(n_8_0_6556), .B1(n_8_0_5460), .B2(n_8_0_253), 
      .ZN(n_8_0_4648));
   OAI21_X1 i_8_0_4843 (.A(n_8_0_5224), .B1(n_8_0_6795), .B2(n_8_0_253), 
      .ZN(n_8_0_4649));
   OAI21_X1 i_8_0_4844 (.A(n_8_0_4652), .B1(n_8_0_4651), .B2(n_8_0_6369), 
      .ZN(n_8_0_4650));
   OAI211_X1 i_8_0_4845 (.A(n_8_0_7011), .B(n_8_0_5894), .C1(n_8_0_6755), 
      .C2(n_8_0_379), .ZN(n_8_0_4651));
   AOI21_X1 i_8_0_4846 (.A(n_8_0_5456), .B1(n_8_0_6590), .B2(n_8_0_379), 
      .ZN(n_8_0_4652));
   AOI21_X1 i_8_0_4847 (.A(n_8_0_6853), .B1(n_8_0_4657), .B2(n_8_0_4653), 
      .ZN(n_138));
   NOR4_X1 i_8_0_4848 (.A1(n_8_0_4654), .A2(n_8_0_4655), .A3(n_8_0_4667), 
      .A4(n_8_0_4672), .ZN(n_8_0_4653));
   NAND4_X1 i_8_0_4849 (.A1(n_8_0_4670), .A2(n_8_0_4664), .A3(n_8_0_4661), 
      .A4(n_8_0_4674), .ZN(n_8_0_4654));
   AOI221_X1 i_8_0_4850 (.A(n_8_0_5395), .B1(n_8_0_5263), .B2(n_8_0_5548), 
      .C1(n_8_0_4656), .C2(n_8_0_65), .ZN(n_8_0_4655));
   OAI21_X1 i_8_0_4851 (.A(n_8_0_6527), .B1(n_8_0_5547), .B2(\out_bs[1] [5]), 
      .ZN(n_8_0_4656));
   AOI21_X1 i_8_0_4852 (.A(n_8_0_4658), .B1(n_8_0_6233), .B2(n_8_0_4659), 
      .ZN(n_8_0_4657));
   NOR2_X1 i_8_0_4853 (.A1(n_8_0_443), .A2(n_8_0_4660), .ZN(n_8_0_4658));
   NAND2_X1 i_8_0_4854 (.A1(n_8_0_443), .A2(n_8_0_4660), .ZN(n_8_0_4659));
   OAI21_X1 i_8_0_4855 (.A(\out_bs[7] [6]), .B1(n_8_0_5560), .B2(\out_bs[7] [5]), 
      .ZN(n_8_0_4660));
   OAI21_X1 i_8_0_4856 (.A(n_8_0_4663), .B1(n_8_0_4662), .B2(n_8_0_6399), 
      .ZN(n_8_0_4661));
   OAI21_X1 i_8_0_4857 (.A(n_8_0_4835), .B1(n_8_0_6772), .B2(n_8_0_128), 
      .ZN(n_8_0_4662));
   AOI21_X1 i_8_0_4858 (.A(n_8_0_5428), .B1(n_8_0_6606), .B2(n_8_0_128), 
      .ZN(n_8_0_4663));
   OAI21_X1 i_8_0_4859 (.A(n_8_0_4665), .B1(n_8_0_4666), .B2(n_8_0_5554), 
      .ZN(n_8_0_4664));
   OAI21_X1 i_8_0_4860 (.A(n_8_0_6249), .B1(n_8_0_5274), .B2(n_8_0_0), .ZN(
      n_8_0_4665));
   OAI21_X1 i_8_0_4861 (.A(n_8_0_7084), .B1(n_8_0_0), .B2(n_8_0_6811), .ZN(
      n_8_0_4666));
   OAI21_X1 i_8_0_4862 (.A(n_8_0_4668), .B1(n_8_0_6837), .B2(n_8_0_191), 
      .ZN(n_8_0_4667));
   OAI211_X1 i_8_0_4863 (.A(n_8_0_4669), .B(\out_bs[3] [6]), .C1(n_8_0_6413), 
      .C2(n_8_0_4829), .ZN(n_8_0_4668));
   NAND2_X1 i_8_0_4864 (.A1(n_8_0_6844), .A2(n_8_0_191), .ZN(n_8_0_4669));
   AOI22_X1 i_8_0_4865 (.A1(n_8_0_6903), .A2(n_8_0_6825), .B1(n_8_0_4671), 
      .B2(\out_bs[5] [6]), .ZN(n_8_0_4670));
   AOI22_X1 i_8_0_4866 (.A1(n_8_0_6619), .A2(n_8_0_317), .B1(n_8_0_5054), 
      .B2(n_8_0_6098), .ZN(n_8_0_4671));
   AOI221_X1 i_8_0_4867 (.A(n_8_0_5460), .B1(n_8_0_254), .B2(n_8_0_6556), 
      .C1(n_8_0_4673), .C2(n_8_0_6093), .ZN(n_8_0_4672));
   AOI21_X1 i_8_0_4868 (.A(n_8_0_5223), .B1(n_8_0_6794), .B2(n_8_0_6918), 
      .ZN(n_8_0_4673));
   AOI22_X1 i_8_0_4869 (.A1(n_8_0_6894), .A2(n_8_0_6754), .B1(n_8_0_4676), 
      .B2(n_8_0_4675), .ZN(n_8_0_4674));
   OAI21_X1 i_8_0_4870 (.A(n_8_0_6590), .B1(n_8_0_5456), .B2(n_8_0_380), 
      .ZN(n_8_0_4675));
   NAND2_X1 i_8_0_4871 (.A1(n_8_0_5543), .A2(n_8_0_7011), .ZN(n_8_0_4676));
   NOR2_X1 i_8_0_4872 (.A1(n_8_0_4677), .A2(n_8_0_6853), .ZN(n_139));
   NOR3_X1 i_8_0_4873 (.A1(n_8_0_4678), .A2(n_8_0_4692), .A3(n_8_0_4679), 
      .ZN(n_8_0_4677));
   NAND4_X1 i_8_0_4874 (.A1(n_8_0_4701), .A2(n_8_0_4698), .A3(n_8_0_4695), 
      .A4(n_8_0_4683), .ZN(n_8_0_4678));
   OAI221_X1 i_8_0_4875 (.A(n_8_0_4680), .B1(n_8_0_6232), .B2(n_8_0_444), 
      .C1(n_8_0_3), .C2(n_8_0_6811), .ZN(n_8_0_4679));
   NOR3_X1 i_8_0_4876 (.A1(n_8_0_4689), .A2(n_8_0_4682), .A3(n_8_0_4681), 
      .ZN(n_8_0_4680));
   AOI21_X1 i_8_0_4877 (.A(n_8_0_4686), .B1(n_8_0_6232), .B2(n_8_0_444), 
      .ZN(n_8_0_4681));
   AOI21_X1 i_8_0_4878 (.A(n_8_0_4687), .B1(n_8_0_6812), .B2(n_8_0_3), .ZN(
      n_8_0_4682));
   OAI21_X1 i_8_0_4879 (.A(n_8_0_5394), .B1(n_8_0_4685), .B2(n_8_0_4684), 
      .ZN(n_8_0_4683));
   AOI22_X1 i_8_0_4880 (.A1(n_8_0_6526), .A2(n_8_0_66), .B1(n_8_0_4840), 
      .B2(n_8_0_6448), .ZN(n_8_0_4684));
   NOR2_X1 i_8_0_4881 (.A1(n_8_0_66), .A2(n_8_0_6782), .ZN(n_8_0_4685));
   OAI21_X1 i_8_0_4882 (.A(\out_bs[7] [6]), .B1(n_8_0_6475), .B2(n_8_0_4823), 
      .ZN(n_8_0_4686));
   AOI21_X1 i_8_0_4883 (.A(n_8_0_6671), .B1(n_8_0_5595), .B2(\out_bs[0] [6]), 
      .ZN(n_8_0_4687));
   INV_X1 i_8_0_4884 (.A(n_8_0_4689), .ZN(n_8_0_4688));
   OAI21_X1 i_8_0_4885 (.A(n_8_0_4690), .B1(n_8_0_6837), .B2(n_8_0_192), 
      .ZN(n_8_0_4689));
   OAI211_X1 i_8_0_4886 (.A(n_8_0_4691), .B(\out_bs[3] [6]), .C1(n_8_0_6428), 
      .C2(n_8_0_4829), .ZN(n_8_0_4690));
   NAND2_X1 i_8_0_4887 (.A1(n_8_0_6844), .A2(n_8_0_192), .ZN(n_8_0_4691));
   AOI211_X1 i_8_0_4888 (.A(n_8_0_5428), .B(n_8_0_4693), .C1(n_8_0_129), 
      .C2(n_8_0_6606), .ZN(n_8_0_4692));
   INV_X1 i_8_0_4889 (.A(n_8_0_4694), .ZN(n_8_0_4693));
   OAI211_X1 i_8_0_4890 (.A(n_8_0_6453), .B(n_8_0_4835), .C1(n_8_0_6772), 
      .C2(n_8_0_129), .ZN(n_8_0_4694));
   OAI21_X1 i_8_0_4891 (.A(n_8_0_4697), .B1(n_8_0_4696), .B2(n_8_0_6113), 
      .ZN(n_8_0_4695));
   OAI21_X1 i_8_0_4892 (.A(n_8_0_5224), .B1(n_8_0_6795), .B2(n_8_0_255), 
      .ZN(n_8_0_4696));
   OAI21_X1 i_8_0_4893 (.A(n_8_0_6556), .B1(n_8_0_5460), .B2(n_8_0_255), 
      .ZN(n_8_0_4697));
   OAI21_X1 i_8_0_4894 (.A(n_8_0_4700), .B1(n_8_0_4699), .B2(n_8_0_6136), 
      .ZN(n_8_0_4698));
   OAI21_X1 i_8_0_4895 (.A(n_8_0_5054), .B1(n_8_0_6824), .B2(n_8_0_318), 
      .ZN(n_8_0_4699));
   AOI21_X1 i_8_0_4896 (.A(n_8_0_5302), .B1(n_8_0_6513), .B2(n_8_0_318), 
      .ZN(n_8_0_4700));
   OAI21_X1 i_8_0_4897 (.A(n_8_0_4703), .B1(n_8_0_4702), .B2(n_8_0_4826), 
      .ZN(n_8_0_4701));
   OAI21_X1 i_8_0_4898 (.A(n_8_0_6481), .B1(n_8_0_6755), .B2(n_8_0_381), 
      .ZN(n_8_0_4702));
   OAI21_X1 i_8_0_4899 (.A(n_8_0_6590), .B1(n_8_0_5456), .B2(n_8_0_381), 
      .ZN(n_8_0_4703));
   AOI21_X1 i_8_0_4900 (.A(n_8_0_6853), .B1(n_8_0_4709), .B2(n_8_0_4704), 
      .ZN(n_140));
   NOR4_X1 i_8_0_4901 (.A1(n_8_0_4726), .A2(n_8_0_4705), .A3(n_8_0_4720), 
      .A4(n_8_0_4729), .ZN(n_8_0_4704));
   NAND2_X1 i_8_0_4902 (.A1(n_8_0_4723), .A2(n_8_0_4706), .ZN(n_8_0_4705));
   AOI21_X1 i_8_0_4903 (.A(n_8_0_4707), .B1(n_8_0_6838), .B2(n_8_0_6937), 
      .ZN(n_8_0_4706));
   AOI21_X1 i_8_0_4904 (.A(n_8_0_4708), .B1(n_8_0_6844), .B2(n_8_0_193), 
      .ZN(n_8_0_4707));
   OAI21_X1 i_8_0_4905 (.A(\out_bs[3] [6]), .B1(n_8_0_4829), .B2(\out_bs[3] [2]), 
      .ZN(n_8_0_4708));
   NOR2_X1 i_8_0_4906 (.A1(n_8_0_4717), .A2(n_8_0_4710), .ZN(n_8_0_4709));
   NAND2_X1 i_8_0_4907 (.A1(n_8_0_4714), .A2(n_8_0_4711), .ZN(n_8_0_4710));
   NAND2_X1 i_8_0_4908 (.A1(n_8_0_4713), .A2(n_8_0_4712), .ZN(n_8_0_4711));
   AOI21_X1 i_8_0_4909 (.A(n_8_0_5395), .B1(n_8_0_6526), .B2(n_8_0_67), .ZN(
      n_8_0_4712));
   OAI211_X1 i_8_0_4910 (.A(n_8_0_7068), .B(n_8_0_4840), .C1(n_8_0_6782), 
      .C2(n_8_0_67), .ZN(n_8_0_4713));
   OAI21_X1 i_8_0_4911 (.A(n_8_0_4715), .B1(n_8_0_6729), .B2(n_8_0_6874), 
      .ZN(n_8_0_4714));
   OAI21_X1 i_8_0_4912 (.A(n_8_0_4716), .B1(n_8_0_6730), .B2(n_8_0_445), 
      .ZN(n_8_0_4715));
   OAI21_X1 i_8_0_4913 (.A(\out_bs[7] [6]), .B1(n_8_0_4823), .B2(\out_bs[7] [2]), 
      .ZN(n_8_0_4716));
   OAI21_X1 i_8_0_4914 (.A(n_8_0_4718), .B1(n_8_0_6824), .B2(n_8_0_319), 
      .ZN(n_8_0_4717));
   OAI21_X1 i_8_0_4915 (.A(n_8_0_4719), .B1(n_8_0_5053), .B2(n_8_0_6165), 
      .ZN(n_8_0_4718));
   AOI21_X1 i_8_0_4916 (.A(n_8_0_7024), .B1(n_8_0_6619), .B2(n_8_0_319), 
      .ZN(n_8_0_4719));
   AND2_X1 i_8_0_4917 (.A1(n_8_0_4722), .A2(n_8_0_4721), .ZN(n_8_0_4720));
   OAI211_X1 i_8_0_4918 (.A(n_8_0_7034), .B(n_8_0_5607), .C1(n_8_0_6795), 
      .C2(n_8_0_256), .ZN(n_8_0_4721));
   OAI21_X1 i_8_0_4919 (.A(n_8_0_6556), .B1(n_8_0_5460), .B2(n_8_0_256), 
      .ZN(n_8_0_4722));
   OAI21_X1 i_8_0_4920 (.A(n_8_0_4724), .B1(n_8_0_4725), .B2(\out_bs[2] [2]), 
      .ZN(n_8_0_4723));
   AOI21_X1 i_8_0_4921 (.A(n_8_0_5428), .B1(n_8_0_6606), .B2(n_8_0_130), 
      .ZN(n_8_0_4724));
   OAI21_X1 i_8_0_4922 (.A(n_8_0_4835), .B1(n_8_0_6772), .B2(n_8_0_130), 
      .ZN(n_8_0_4725));
   AOI211_X1 i_8_0_4923 (.A(n_8_0_5456), .B(n_8_0_4727), .C1(n_8_0_382), 
      .C2(n_8_0_6590), .ZN(n_8_0_4726));
   AOI21_X1 i_8_0_4924 (.A(n_8_0_4728), .B1(n_8_0_6754), .B2(n_8_0_6893), 
      .ZN(n_8_0_4727));
   NAND2_X1 i_8_0_4925 (.A1(n_8_0_5626), .A2(n_8_0_7011), .ZN(n_8_0_4728));
   AOI211_X1 i_8_0_4926 (.A(n_8_0_5274), .B(n_8_0_4730), .C1(n_8_0_1), .C2(
      n_8_0_6249), .ZN(n_8_0_4729));
   NOR2_X1 i_8_0_4927 (.A1(n_8_0_4731), .A2(\out_bs[0] [2]), .ZN(n_8_0_4730));
   OAI211_X1 i_8_0_4928 (.A(n_8_0_7084), .B(n_8_0_5944), .C1(n_8_0_6811), 
      .C2(n_8_0_1), .ZN(n_8_0_4731));
   AOI21_X1 i_8_0_4929 (.A(n_8_0_6853), .B1(n_8_0_4732), .B2(n_8_0_4738), 
      .ZN(n_141));
   AOI211_X1 i_8_0_4930 (.A(n_8_0_4745), .B(n_8_0_4733), .C1(n_8_0_4744), 
      .C2(n_8_0_6233), .ZN(n_8_0_4732));
   NAND3_X1 i_8_0_4931 (.A1(n_8_0_4734), .A2(n_8_0_4747), .A3(n_8_0_4750), 
      .ZN(n_8_0_4733));
   NOR3_X1 i_8_0_4932 (.A1(n_8_0_4760), .A2(n_8_0_4753), .A3(n_8_0_4735), 
      .ZN(n_8_0_4734));
   NAND3_X1 i_8_0_4933 (.A1(n_8_0_4736), .A2(n_8_0_4741), .A3(n_8_0_4836), 
      .ZN(n_8_0_4735));
   AOI21_X1 i_8_0_4934 (.A(n_8_0_4756), .B1(n_8_0_4737), .B2(\out_bs[0] [6]), 
      .ZN(n_8_0_4736));
   AOI21_X1 i_8_0_4935 (.A(n_8_0_6523), .B1(n_8_0_6812), .B2(n_8_0_2), .ZN(
      n_8_0_4737));
   OAI21_X1 i_8_0_4936 (.A(n_8_0_4739), .B1(n_8_0_4740), .B2(n_8_0_6536), 
      .ZN(n_8_0_4738));
   OAI21_X1 i_8_0_4937 (.A(n_8_0_6606), .B1(n_8_0_5428), .B2(n_8_0_131), 
      .ZN(n_8_0_4739));
   OAI21_X1 i_8_0_4938 (.A(n_8_0_4835), .B1(n_8_0_6772), .B2(n_8_0_131), 
      .ZN(n_8_0_4740));
   NAND2_X1 i_8_0_4939 (.A1(n_8_0_4743), .A2(n_8_0_4742), .ZN(n_8_0_4741));
   OAI211_X1 i_8_0_4940 (.A(n_8_0_4773), .B(n_8_0_6698), .C1(n_8_0_6782), 
      .C2(n_8_0_68), .ZN(n_8_0_4742));
   AOI21_X1 i_8_0_4941 (.A(n_8_0_5395), .B1(n_8_0_6526), .B2(n_8_0_68), .ZN(
      n_8_0_4743));
   NAND2_X1 i_8_0_4942 (.A1(n_8_0_4746), .A2(n_8_0_446), .ZN(n_8_0_4744));
   NOR2_X1 i_8_0_4943 (.A1(n_8_0_4746), .A2(n_8_0_446), .ZN(n_8_0_4745));
   OAI21_X1 i_8_0_4944 (.A(\out_bs[7] [6]), .B1(n_8_0_6542), .B2(n_8_0_4823), 
      .ZN(n_8_0_4746));
   AOI21_X1 i_8_0_4945 (.A(n_8_0_4748), .B1(n_8_0_6838), .B2(n_8_0_6936), 
      .ZN(n_8_0_4747));
   AOI21_X1 i_8_0_4946 (.A(n_8_0_4749), .B1(n_8_0_6844), .B2(n_8_0_194), 
      .ZN(n_8_0_4748));
   OAI21_X1 i_8_0_4947 (.A(\out_bs[3] [6]), .B1(n_8_0_6565), .B2(n_8_0_4829), 
      .ZN(n_8_0_4749));
   OAI21_X1 i_8_0_4948 (.A(n_8_0_4752), .B1(n_8_0_4751), .B2(n_8_0_6191), 
      .ZN(n_8_0_4750));
   OAI21_X1 i_8_0_4949 (.A(n_8_0_5224), .B1(n_8_0_6795), .B2(n_8_0_257), 
      .ZN(n_8_0_4751));
   OAI21_X1 i_8_0_4950 (.A(n_8_0_6556), .B1(n_8_0_5460), .B2(n_8_0_257), 
      .ZN(n_8_0_4752));
   OAI21_X1 i_8_0_4951 (.A(n_8_0_4754), .B1(n_8_0_6824), .B2(n_8_0_320), 
      .ZN(n_8_0_4753));
   OAI211_X1 i_8_0_4952 (.A(n_8_0_4755), .B(\out_bs[5] [6]), .C1(n_8_0_6210), 
      .C2(n_8_0_5053), .ZN(n_8_0_4754));
   NAND2_X1 i_8_0_4953 (.A1(n_8_0_6619), .A2(n_8_0_320), .ZN(n_8_0_4755));
   INV_X1 i_8_0_4954 (.A(n_8_0_4757), .ZN(n_8_0_4756));
   OAI21_X1 i_8_0_4955 (.A(n_8_0_4759), .B1(n_8_0_4758), .B2(n_8_0_4826), 
      .ZN(n_8_0_4757));
   OAI21_X1 i_8_0_4956 (.A(n_8_0_6551), .B1(n_8_0_6755), .B2(n_8_0_383), 
      .ZN(n_8_0_4758));
   OAI21_X1 i_8_0_4957 (.A(n_8_0_6590), .B1(n_8_0_5456), .B2(n_8_0_383), 
      .ZN(n_8_0_4759));
   AOI21_X1 i_8_0_4958 (.A(n_8_0_2), .B1(n_8_0_6595), .B2(n_8_0_5803), .ZN(
      n_8_0_4760));
   AOI21_X1 i_8_0_4959 (.A(n_8_0_6853), .B1(n_8_0_4777), .B2(n_8_0_4761), 
      .ZN(n_142));
   AND3_X1 i_8_0_4960 (.A1(n_8_0_4762), .A2(n_8_0_4771), .A3(n_8_0_4774), 
      .ZN(n_8_0_4761));
   AOI211_X1 i_8_0_4961 (.A(n_8_0_4767), .B(n_8_0_4763), .C1(n_8_0_4766), 
      .C2(\out_bs[0] [6]), .ZN(n_8_0_4762));
   AOI221_X1 i_8_0_4962 (.A(n_8_0_5428), .B1(n_8_0_6606), .B2(n_8_0_132), 
      .C1(n_8_0_6612), .C2(n_8_0_4764), .ZN(n_8_0_4763));
   INV_X1 i_8_0_4963 (.A(n_8_0_4765), .ZN(n_8_0_4764));
   OAI21_X1 i_8_0_4964 (.A(n_8_0_4835), .B1(n_8_0_6772), .B2(n_8_0_132), 
      .ZN(n_8_0_4765));
   AOI21_X1 i_8_0_4965 (.A(n_8_0_6667), .B1(n_8_0_6812), .B2(n_8_0_6), .ZN(
      n_8_0_4766));
   OAI211_X1 i_8_0_4966 (.A(n_8_0_4836), .B(n_8_0_4768), .C1(n_8_0_6232), 
      .C2(n_8_0_4769), .ZN(n_8_0_4767));
   OR2_X1 i_8_0_4967 (.A1(n_8_0_447), .A2(n_8_0_4770), .ZN(n_8_0_4768));
   AND2_X1 i_8_0_4968 (.A1(n_8_0_447), .A2(n_8_0_4770), .ZN(n_8_0_4769));
   OAI21_X1 i_8_0_4969 (.A(\out_bs[7] [6]), .B1(n_8_0_6237), .B2(n_8_0_5056), 
      .ZN(n_8_0_4770));
   OAI211_X1 i_8_0_4970 (.A(n_8_0_5394), .B(n_8_0_4772), .C1(n_8_0_5262), 
      .C2(n_8_0_5668), .ZN(n_8_0_4771));
   OAI21_X1 i_8_0_4971 (.A(n_8_0_69), .B1(n_8_0_6526), .B2(n_8_0_4773), .ZN(
      n_8_0_4772));
   NOR2_X1 i_8_0_4972 (.A1(n_8_0_5668), .A2(\out_bs[1] [5]), .ZN(n_8_0_4773));
   AOI21_X1 i_8_0_4973 (.A(n_8_0_4775), .B1(n_8_0_6838), .B2(n_8_0_6935), 
      .ZN(n_8_0_4774));
   AOI21_X1 i_8_0_4974 (.A(n_8_0_4776), .B1(n_8_0_6844), .B2(n_8_0_195), 
      .ZN(n_8_0_4775));
   OAI21_X1 i_8_0_4975 (.A(\out_bs[3] [6]), .B1(n_8_0_4829), .B2(n_8_0_6653), 
      .ZN(n_8_0_4776));
   NOR4_X1 i_8_0_4976 (.A1(n_8_0_4787), .A2(n_8_0_4784), .A3(n_8_0_4781), 
      .A4(n_8_0_4778), .ZN(n_8_0_4777));
   INV_X1 i_8_0_4977 (.A(n_8_0_4779), .ZN(n_8_0_4778));
   OAI211_X1 i_8_0_4978 (.A(n_8_0_5459), .B(n_8_0_4780), .C1(n_8_0_5458), 
      .C2(n_8_0_5690), .ZN(n_8_0_4779));
   OAI211_X1 i_8_0_4979 (.A(n_8_0_258), .B(n_8_0_6554), .C1(n_8_0_6556), 
      .C2(n_8_0_5691), .ZN(n_8_0_4780));
   OAI21_X1 i_8_0_4980 (.A(n_8_0_4782), .B1(n_8_0_6755), .B2(n_8_0_384), 
      .ZN(n_8_0_4781));
   OAI211_X1 i_8_0_4981 (.A(n_8_0_5455), .B(n_8_0_4783), .C1(\out_bs[6] [5]), 
      .C2(n_8_0_5677), .ZN(n_8_0_4782));
   NAND2_X1 i_8_0_4982 (.A1(n_8_0_6590), .A2(n_8_0_384), .ZN(n_8_0_4783));
   AOI221_X1 i_8_0_4983 (.A(n_8_0_5302), .B1(n_8_0_6513), .B2(n_8_0_321), 
      .C1(n_8_0_7023), .C2(n_8_0_4785), .ZN(n_8_0_4784));
   INV_X1 i_8_0_4984 (.A(n_8_0_4786), .ZN(n_8_0_4785));
   OAI21_X1 i_8_0_4985 (.A(n_8_0_5682), .B1(n_8_0_6824), .B2(n_8_0_321), 
      .ZN(n_8_0_4786));
   AOI21_X1 i_8_0_4986 (.A(n_8_0_6), .B1(n_8_0_6595), .B2(n_8_0_5803), .ZN(
      n_8_0_4787));
   AOI21_X1 i_8_0_4987 (.A(n_8_0_6853), .B1(n_8_0_4788), .B2(n_8_0_4811), 
      .ZN(n_143));
   NOR4_X1 i_8_0_4988 (.A1(n_8_0_4808), .A2(n_8_0_4799), .A3(n_8_0_4796), 
      .A4(n_8_0_4789), .ZN(n_8_0_4788));
   NAND4_X1 i_8_0_4989 (.A1(n_8_0_4805), .A2(n_8_0_4790), .A3(n_8_0_4801), 
      .A4(n_8_0_4793), .ZN(n_8_0_4789));
   OAI211_X1 i_8_0_4990 (.A(n_8_0_5455), .B(n_8_0_4791), .C1(n_8_0_5451), 
      .C2(n_8_0_5722), .ZN(n_8_0_4790));
   OAI21_X1 i_8_0_4991 (.A(n_8_0_385), .B1(n_8_0_6590), .B2(n_8_0_4792), 
      .ZN(n_8_0_4791));
   NOR2_X1 i_8_0_4992 (.A1(n_8_0_5722), .A2(\out_bs[6] [5]), .ZN(n_8_0_4792));
   OAI21_X1 i_8_0_4993 (.A(n_8_0_4795), .B1(n_8_0_4794), .B2(n_8_0_6666), 
      .ZN(n_8_0_4793));
   OAI211_X1 i_8_0_4994 (.A(n_8_0_7084), .B(n_8_0_5944), .C1(n_8_0_6811), 
      .C2(n_8_0_7), .ZN(n_8_0_4794));
   AOI21_X1 i_8_0_4995 (.A(n_8_0_5274), .B1(n_8_0_6249), .B2(n_8_0_7), .ZN(
      n_8_0_4795));
   OAI21_X1 i_8_0_4996 (.A(n_8_0_4797), .B1(n_8_0_6837), .B2(n_8_0_196), 
      .ZN(n_8_0_4796));
   OAI211_X1 i_8_0_4997 (.A(n_8_0_4798), .B(\out_bs[3] [6]), .C1(\out_bs[3] [5]), 
      .C2(n_8_0_5697), .ZN(n_8_0_4797));
   NAND2_X1 i_8_0_4998 (.A1(n_8_0_6844), .A2(n_8_0_196), .ZN(n_8_0_4798));
   AOI221_X1 i_8_0_4999 (.A(n_8_0_5428), .B1(n_8_0_5426), .B2(n_8_0_5707), 
      .C1(n_8_0_4800), .C2(n_8_0_133), .ZN(n_8_0_4799));
   OAI21_X1 i_8_0_5000 (.A(n_8_0_6607), .B1(n_8_0_5706), .B2(\out_bs[2] [5]), 
      .ZN(n_8_0_4800));
   AOI21_X1 i_8_0_5001 (.A(n_8_0_4803), .B1(n_8_0_6731), .B2(n_8_0_4802), 
      .ZN(n_8_0_4801));
   NAND2_X1 i_8_0_5002 (.A1(n_8_0_4804), .A2(n_8_0_448), .ZN(n_8_0_4802));
   NOR2_X1 i_8_0_5003 (.A1(n_8_0_4804), .A2(n_8_0_448), .ZN(n_8_0_4803));
   OAI21_X1 i_8_0_5004 (.A(\out_bs[7] [6]), .B1(n_8_0_6723), .B2(n_8_0_4823), 
      .ZN(n_8_0_4804));
   OAI21_X1 i_8_0_5005 (.A(n_8_0_4806), .B1(n_8_0_5262), .B2(n_8_0_5711), 
      .ZN(n_8_0_4805));
   AOI21_X1 i_8_0_5006 (.A(n_8_0_5395), .B1(n_8_0_4807), .B2(n_8_0_70), .ZN(
      n_8_0_4806));
   OAI21_X1 i_8_0_5007 (.A(n_8_0_6527), .B1(n_8_0_5711), .B2(\out_bs[1] [5]), 
      .ZN(n_8_0_4807));
   AOI211_X1 i_8_0_5008 (.A(n_8_0_5460), .B(n_8_0_4809), .C1(n_8_0_259), 
      .C2(n_8_0_6556), .ZN(n_8_0_4808));
   NOR3_X1 i_8_0_5009 (.A1(\out_bs[4] [5]), .A2(n_8_0_4810), .A3(n_8_0_5728), 
      .ZN(n_8_0_4809));
   NOR2_X1 i_8_0_5010 (.A1(n_8_0_259), .A2(n_8_0_6795), .ZN(n_8_0_4810));
   OAI21_X1 i_8_0_5011 (.A(n_8_0_4812), .B1(n_8_0_4813), .B2(n_8_0_6299), 
      .ZN(n_8_0_4811));
   OAI21_X1 i_8_0_5012 (.A(n_8_0_6513), .B1(n_8_0_5302), .B2(n_8_0_322), 
      .ZN(n_8_0_4812));
   OAI21_X1 i_8_0_5013 (.A(n_8_0_5054), .B1(n_8_0_6824), .B2(n_8_0_322), 
      .ZN(n_8_0_4813));
   OAI21_X1 i_8_0_5018 (.A(n_8_0_323), .B1(n_8_0_6619), .B2(n_8_0_4818), 
      .ZN(n_8_0_4817));
   INV_X1 i_8_0_5019 (.A(n_8_0_4819), .ZN(n_8_0_4818));
   AOI21_X1 i_8_0_5020 (.A(n_8_0_7024), .B1(n_8_0_5054), .B2(n_8_0_7021), 
      .ZN(n_8_0_4819));
   OAI211_X1 i_8_0_5026 (.A(\out_bs[6] [6]), .B(n_8_0_4826), .C1(n_8_0_6759), 
      .C2(n_8_0_6892), .ZN(n_8_0_4825));
   NAND2_X1 i_8_0_5027 (.A1(n_8_0_5894), .A2(n_8_0_7011), .ZN(n_8_0_4826));
   OAI211_X1 i_8_0_5029 (.A(\out_bs[3] [6]), .B(n_8_0_4829), .C1(n_8_0_6843), 
      .C2(n_8_0_6934), .ZN(n_8_0_4828));
   NAND2_X1 i_8_0_5030 (.A1(n_8_0_6008), .A2(n_8_0_7046), .ZN(n_8_0_4829));
   NAND2_X1 i_8_0_5032 (.A1(n_8_0_4836), .A2(n_8_0_4832), .ZN(n_8_0_4831));
   OAI21_X1 i_8_0_5033 (.A(n_8_0_4833), .B1(n_8_0_6773), .B2(n_8_0_6961), 
      .ZN(n_8_0_4832));
   OAI22_X1 i_8_0_5034 (.A1(n_8_0_134), .A2(n_8_0_6772), .B1(n_8_0_4835), 
      .B2(n_8_0_7060), .ZN(n_8_0_4833));
   NAND2_X1 i_8_0_5035 (.A1(n_8_0_5815), .A2(n_8_0_7059), .ZN(n_8_0_4834));
   NOR2_X1 i_8_0_5036 (.A1(n_8_0_5814), .A2(\out_bs[2] [5]), .ZN(n_8_0_4835));
   OAI21_X1 i_8_0_5037 (.A(n_8_0_6250), .B1(n_8_0_5943), .B2(\out_bs[0] [5]), 
      .ZN(n_8_0_4836));
   OAI22_X1 i_8_0_5038 (.A1(n_8_0_71), .A2(n_8_0_6782), .B1(n_8_0_4838), 
      .B2(n_8_0_7072), .ZN(n_8_0_4837));
   INV_X1 i_8_0_5039 (.A(n_8_0_4839), .ZN(n_8_0_4838));
   AOI21_X1 i_8_0_5040 (.A(n_8_0_4840), .B1(n_8_0_6784), .B2(n_8_0_71), .ZN(
      n_8_0_4839));
   NOR2_X1 i_8_0_5041 (.A1(n_8_0_5983), .A2(\out_bs[1] [5]), .ZN(n_8_0_4840));
   AOI21_X1 i_8_0_5042 (.A(n_8_0_8), .B1(n_8_0_6595), .B2(n_8_0_5803), .ZN(
      n_8_0_4841));
   AOI221_X1 i_8_0_5043 (.A(n_8_0_5460), .B1(n_8_0_6556), .B2(n_8_0_260), 
      .C1(n_8_0_4843), .C2(n_8_0_7032), .ZN(n_8_0_4842));
   AOI21_X1 i_8_0_5044 (.A(n_8_0_5223), .B1(n_8_0_6794), .B2(n_8_0_6917), 
      .ZN(n_8_0_4843));
   INV_X1 i_8_0_5054 (.A(n_8_0_4853), .ZN(n_8_0_4852));
   OAI21_X1 i_8_0_5055 (.A(n_8_0_5779), .B1(n_8_0_6772), .B2(n_8_0_135), 
      .ZN(n_8_0_4853));
   AOI21_X1 i_8_0_5056 (.A(n_8_0_4855), .B1(n_8_0_6526), .B2(n_8_0_72), .ZN(
      n_8_0_4854));
   OAI21_X1 i_8_0_5057 (.A(n_8_0_5394), .B1(n_8_0_4856), .B2(\out_bs[1] [5]), 
      .ZN(n_8_0_4855));
   OAI21_X1 i_8_0_5058 (.A(n_8_0_5758), .B1(n_8_0_6782), .B2(n_8_0_72), .ZN(
      n_8_0_4856));
   OAI21_X1 i_8_0_5059 (.A(n_8_0_4859), .B1(n_8_0_4858), .B2(n_8_0_387), 
      .ZN(n_8_0_4857));
   OAI21_X1 i_8_0_5060 (.A(n_8_0_5455), .B1(n_8_0_5451), .B2(n_8_0_5767), 
      .ZN(n_8_0_4858));
   OAI21_X1 i_8_0_5061 (.A(n_8_0_6591), .B1(n_8_0_5767), .B2(\out_bs[6] [5]), 
      .ZN(n_8_0_4859));
   INV_X1 i_8_0_5062 (.A(n_8_0_4861), .ZN(n_8_0_4860));
   OAI21_X1 i_8_0_5064 (.A(n_8_0_4863), .B1(n_8_0_5787), .B2(\out_bs[3] [5]), 
      .ZN(n_8_0_4862));
   AOI21_X1 i_8_0_5065 (.A(n_8_0_7047), .B1(n_8_0_6844), .B2(n_8_0_198), 
      .ZN(n_8_0_4863));
   OAI21_X1 i_8_0_5067 (.A(n_8_0_6350), .B1(n_8_0_6795), .B2(n_8_0_261), 
      .ZN(n_8_0_4865));
   OAI21_X1 i_8_0_5068 (.A(n_8_0_6556), .B1(n_8_0_5460), .B2(n_8_0_261), 
      .ZN(n_8_0_4866));
   OAI211_X1 i_8_0_5070 (.A(n_8_0_4869), .B(\out_bs[5] [6]), .C1(n_8_0_6374), 
      .C2(n_8_0_5053), .ZN(n_8_0_4868));
   NAND2_X1 i_8_0_5071 (.A1(n_8_0_6619), .A2(n_8_0_324), .ZN(n_8_0_4869));
   AOI22_X1 i_8_0_5072 (.A1(n_8_0_9), .A2(n_8_0_4872), .B1(n_8_0_4871), .B2(
      n_8_0_6811), .ZN(n_8_0_4870));
   OAI21_X1 i_8_0_5073 (.A(\out_bs[0] [6]), .B1(\out_bs[0] [5]), .B2(n_8_0_5771), 
      .ZN(n_8_0_4871));
   OAI21_X1 i_8_0_5074 (.A(n_8_0_6250), .B1(n_8_0_5771), .B2(\out_bs[0] [5]), 
      .ZN(n_8_0_4872));
   AOI21_X1 i_8_0_5075 (.A(n_8_0_6853), .B1(n_8_0_4873), .B2(n_8_0_4878), 
      .ZN(n_144));
   AND3_X1 i_8_0_5076 (.A1(n_8_0_4874), .A2(n_8_0_4882), .A3(n_8_0_4894), 
      .ZN(n_8_0_4873));
   AOI211_X1 i_8_0_5077 (.A(n_8_0_4888), .B(n_8_0_4876), .C1(n_8_0_4875), 
      .C2(\out_bs[0] [6]), .ZN(n_8_0_4874));
   AOI22_X1 i_8_0_5078 (.A1(n_8_0_6812), .A2(n_8_0_10), .B1(n_8_0_7084), 
      .B2(n_8_0_5804), .ZN(n_8_0_4875));
   OAI211_X1 i_8_0_5079 (.A(n_8_0_4877), .B(n_8_0_4891), .C1(n_8_0_6811), 
      .C2(n_8_0_10), .ZN(n_8_0_4876));
   NOR3_X1 i_8_0_5080 (.A1(n_8_0_4887), .A2(n_8_0_4886), .A3(n_8_0_4879), 
      .ZN(n_8_0_4877));
   OAI21_X1 i_8_0_5081 (.A(n_8_0_4898), .B1(n_8_0_4897), .B2(n_8_0_6233), 
      .ZN(n_8_0_4878));
   AOI21_X1 i_8_0_5082 (.A(n_8_0_4880), .B1(n_8_0_6590), .B2(n_8_0_388), 
      .ZN(n_8_0_4879));
   OAI21_X1 i_8_0_5083 (.A(n_8_0_5455), .B1(n_8_0_4881), .B2(\out_bs[6] [5]), 
      .ZN(n_8_0_4880));
   OAI21_X1 i_8_0_5084 (.A(n_8_0_5823), .B1(n_8_0_6755), .B2(n_8_0_388), 
      .ZN(n_8_0_4881));
   OAI21_X1 i_8_0_5085 (.A(n_8_0_4883), .B1(n_8_0_4884), .B2(n_8_0_6381), 
      .ZN(n_8_0_4882));
   OAI21_X1 i_8_0_5086 (.A(n_8_0_6556), .B1(n_8_0_5460), .B2(n_8_0_262), 
      .ZN(n_8_0_4883));
   OAI21_X1 i_8_0_5087 (.A(n_8_0_5224), .B1(n_8_0_6795), .B2(n_8_0_262), 
      .ZN(n_8_0_4884));
   NOR2_X1 i_8_0_5088 (.A1(n_8_0_4887), .A2(n_8_0_4886), .ZN(n_8_0_4885));
   AOI221_X1 i_8_0_5089 (.A(n_8_0_7024), .B1(n_8_0_6408), .B2(n_8_0_5054), 
      .C1(n_8_0_6619), .C2(n_8_0_325), .ZN(n_8_0_4886));
   NOR2_X1 i_8_0_5090 (.A1(n_8_0_6824), .A2(n_8_0_325), .ZN(n_8_0_4887));
   OAI21_X1 i_8_0_5091 (.A(n_8_0_4889), .B1(n_8_0_6837), .B2(n_8_0_199), 
      .ZN(n_8_0_4888));
   OAI211_X1 i_8_0_5092 (.A(n_8_0_4890), .B(\out_bs[3] [6]), .C1(\out_bs[3] [5]), 
      .C2(n_8_0_5793), .ZN(n_8_0_4889));
   NAND2_X1 i_8_0_5093 (.A1(n_8_0_6844), .A2(n_8_0_199), .ZN(n_8_0_4890));
   AOI21_X1 i_8_0_5094 (.A(n_8_0_4892), .B1(n_8_0_6773), .B2(n_8_0_6960), 
      .ZN(n_8_0_4891));
   AOI21_X1 i_8_0_5095 (.A(n_8_0_4893), .B1(n_8_0_6772), .B2(n_8_0_136), 
      .ZN(n_8_0_4892));
   AOI21_X1 i_8_0_5096 (.A(n_8_0_6712), .B1(n_8_0_5813), .B2(\out_bs[2] [6]), 
      .ZN(n_8_0_4893));
   OAI21_X1 i_8_0_5097 (.A(n_8_0_4896), .B1(n_8_0_4895), .B2(\out_bs[1] [5]), 
      .ZN(n_8_0_4894));
   OAI21_X1 i_8_0_5098 (.A(n_8_0_5819), .B1(n_8_0_6782), .B2(n_8_0_73), .ZN(
      n_8_0_4895));
   AOI21_X1 i_8_0_5099 (.A(n_8_0_5395), .B1(n_8_0_6526), .B2(n_8_0_73), .ZN(
      n_8_0_4896));
   NOR2_X1 i_8_0_5100 (.A1(n_8_0_4899), .A2(n_8_0_451), .ZN(n_8_0_4897));
   NAND2_X1 i_8_0_5101 (.A1(n_8_0_4899), .A2(n_8_0_451), .ZN(n_8_0_4898));
   OAI21_X1 i_8_0_5102 (.A(\out_bs[7] [6]), .B1(n_8_0_6404), .B2(n_8_0_5056), 
      .ZN(n_8_0_4899));
   AOI21_X1 i_8_0_5103 (.A(n_8_0_6853), .B1(n_8_0_4900), .B2(n_8_0_4908), 
      .ZN(n_145));
   AOI211_X1 i_8_0_5104 (.A(n_8_0_4901), .B(n_8_0_4902), .C1(n_8_0_4904), 
      .C2(n_8_0_4912), .ZN(n_8_0_4900));
   AOI221_X1 i_8_0_5105 (.A(n_8_0_7085), .B1(n_8_0_7084), .B2(n_8_0_5854), 
      .C1(n_8_0_6812), .C2(n_8_0_11), .ZN(n_8_0_4901));
   OAI211_X1 i_8_0_5106 (.A(n_8_0_4903), .B(n_8_0_4905), .C1(n_8_0_6811), 
      .C2(n_8_0_11), .ZN(n_8_0_4902));
   NOR4_X1 i_8_0_5107 (.A1(n_8_0_4923), .A2(n_8_0_4920), .A3(n_8_0_4917), 
      .A4(n_8_0_4914), .ZN(n_8_0_4903));
   OAI21_X1 i_8_0_5108 (.A(n_8_0_6232), .B1(n_8_0_4913), .B2(n_8_0_452), 
      .ZN(n_8_0_4904));
   OAI21_X1 i_8_0_5109 (.A(n_8_0_4906), .B1(n_8_0_4907), .B2(\out_bs[1] [5]), 
      .ZN(n_8_0_4905));
   AOI21_X1 i_8_0_5110 (.A(n_8_0_5395), .B1(n_8_0_6526), .B2(n_8_0_74), .ZN(
      n_8_0_4906));
   OAI21_X1 i_8_0_5111 (.A(n_8_0_5849), .B1(n_8_0_6782), .B2(n_8_0_74), .ZN(
      n_8_0_4907));
   OAI21_X1 i_8_0_5112 (.A(n_8_0_4910), .B1(n_8_0_4909), .B2(n_8_0_6607), 
      .ZN(n_8_0_4908));
   NOR2_X1 i_8_0_5113 (.A1(n_8_0_137), .A2(n_8_0_5428), .ZN(n_8_0_4909));
   OAI211_X1 i_8_0_5114 (.A(n_8_0_7059), .B(n_8_0_5846), .C1(n_8_0_6772), 
      .C2(n_8_0_137), .ZN(n_8_0_4910));
   NOR2_X1 i_8_0_5115 (.A1(n_8_0_4913), .A2(n_8_0_452), .ZN(n_8_0_4911));
   NAND2_X1 i_8_0_5116 (.A1(n_8_0_4913), .A2(n_8_0_452), .ZN(n_8_0_4912));
   OAI21_X1 i_8_0_5117 (.A(\out_bs[7] [6]), .B1(n_8_0_6474), .B2(n_8_0_5056), 
      .ZN(n_8_0_4913));
   OAI21_X1 i_8_0_5118 (.A(n_8_0_4915), .B1(n_8_0_6837), .B2(n_8_0_200), 
      .ZN(n_8_0_4914));
   OAI211_X1 i_8_0_5119 (.A(n_8_0_4916), .B(\out_bs[3] [6]), .C1(\out_bs[3] [5]), 
      .C2(n_8_0_5858), .ZN(n_8_0_4915));
   NAND2_X1 i_8_0_5120 (.A1(n_8_0_6844), .A2(n_8_0_200), .ZN(n_8_0_4916));
   AOI22_X1 i_8_0_5121 (.A1(n_8_0_4918), .A2(n_8_0_7034), .B1(n_8_0_6556), 
      .B2(n_8_0_4919), .ZN(n_8_0_4917));
   AOI21_X1 i_8_0_5122 (.A(n_8_0_5835), .B1(n_8_0_6794), .B2(n_8_0_6916), 
      .ZN(n_8_0_4918));
   NAND2_X1 i_8_0_5123 (.A1(n_8_0_6916), .A2(n_8_0_5459), .ZN(n_8_0_4919));
   AOI21_X1 i_8_0_5124 (.A(n_8_0_4921), .B1(n_8_0_6590), .B2(n_8_0_389), 
      .ZN(n_8_0_4920));
   OAI21_X1 i_8_0_5125 (.A(n_8_0_5455), .B1(n_8_0_4922), .B2(\out_bs[6] [5]), 
      .ZN(n_8_0_4921));
   OAI21_X1 i_8_0_5126 (.A(n_8_0_5828), .B1(n_8_0_6755), .B2(n_8_0_389), 
      .ZN(n_8_0_4922));
   OAI21_X1 i_8_0_5127 (.A(n_8_0_4924), .B1(n_8_0_6824), .B2(n_8_0_326), 
      .ZN(n_8_0_4923));
   OAI211_X1 i_8_0_5128 (.A(n_8_0_4925), .B(\out_bs[5] [6]), .C1(n_8_0_6460), 
      .C2(n_8_0_5053), .ZN(n_8_0_4924));
   NAND2_X1 i_8_0_5129 (.A1(n_8_0_6619), .A2(n_8_0_326), .ZN(n_8_0_4925));
   AOI21_X1 i_8_0_5130 (.A(n_8_0_6853), .B1(n_8_0_4926), .B2(n_8_0_4945), 
      .ZN(n_146));
   NOR4_X1 i_8_0_5131 (.A1(n_8_0_4927), .A2(n_8_0_4938), .A3(n_8_0_4942), 
      .A4(n_8_0_4931), .ZN(n_8_0_4926));
   NAND4_X1 i_8_0_5132 (.A1(n_8_0_4935), .A2(n_8_0_4928), .A3(n_8_0_4948), 
      .A4(n_8_0_4940), .ZN(n_8_0_4927));
   OAI21_X1 i_8_0_5133 (.A(n_8_0_4930), .B1(n_8_0_4929), .B2(n_8_0_6607), 
      .ZN(n_8_0_4928));
   NOR2_X1 i_8_0_5134 (.A1(n_8_0_138), .A2(n_8_0_5428), .ZN(n_8_0_4929));
   OAI211_X1 i_8_0_5135 (.A(n_8_0_7059), .B(n_8_0_5991), .C1(n_8_0_6772), 
      .C2(n_8_0_138), .ZN(n_8_0_4930));
   OAI21_X1 i_8_0_5136 (.A(n_8_0_4932), .B1(n_8_0_4934), .B2(n_8_0_453), 
      .ZN(n_8_0_4931));
   NAND2_X1 i_8_0_5137 (.A1(n_8_0_6731), .A2(n_8_0_4933), .ZN(n_8_0_4932));
   NAND2_X1 i_8_0_5138 (.A1(n_8_0_4934), .A2(n_8_0_453), .ZN(n_8_0_4933));
   OAI21_X1 i_8_0_5139 (.A(\out_bs[7] [6]), .B1(n_8_0_5953), .B2(\out_bs[7] [5]), 
      .ZN(n_8_0_4934));
   AOI21_X1 i_8_0_5140 (.A(n_8_0_4937), .B1(n_8_0_4936), .B2(\out_bs[5] [6]), 
      .ZN(n_8_0_4935));
   AOI22_X1 i_8_0_5141 (.A1(n_8_0_327), .A2(n_8_0_6824), .B1(n_8_0_6678), 
      .B2(n_8_0_5054), .ZN(n_8_0_4936));
   NOR2_X1 i_8_0_5142 (.A1(n_8_0_6824), .A2(n_8_0_327), .ZN(n_8_0_4937));
   AOI221_X1 i_8_0_5143 (.A(n_8_0_5395), .B1(n_8_0_5263), .B2(n_8_0_5980), 
      .C1(n_8_0_4939), .C2(n_8_0_75), .ZN(n_8_0_4938));
   OAI21_X1 i_8_0_5144 (.A(n_8_0_6527), .B1(n_8_0_5981), .B2(\out_bs[1] [5]), 
      .ZN(n_8_0_4939));
   AOI22_X1 i_8_0_5145 (.A1(\out_bs[3] [6]), .A2(n_8_0_4941), .B1(n_8_0_6838), 
      .B2(n_8_0_6933), .ZN(n_8_0_4940));
   AOI22_X1 i_8_0_5146 (.A1(n_8_0_201), .A2(n_8_0_6844), .B1(n_8_0_5865), 
      .B2(n_8_0_7046), .ZN(n_8_0_4941));
   AOI211_X1 i_8_0_5147 (.A(n_8_0_5274), .B(n_8_0_4943), .C1(n_8_0_12), .C2(
      n_8_0_6249), .ZN(n_8_0_4942));
   NOR2_X1 i_8_0_5148 (.A1(n_8_0_4944), .A2(\out_bs[0] [5]), .ZN(n_8_0_4943));
   OAI21_X1 i_8_0_5149 (.A(n_8_0_5941), .B1(n_8_0_6811), .B2(n_8_0_12), .ZN(
      n_8_0_4944));
   OAI21_X1 i_8_0_5150 (.A(n_8_0_4947), .B1(n_8_0_4946), .B2(\out_bs[6] [5]), 
      .ZN(n_8_0_4945));
   OAI21_X1 i_8_0_5151 (.A(n_8_0_5970), .B1(n_8_0_6755), .B2(n_8_0_390), 
      .ZN(n_8_0_4946));
   OAI21_X1 i_8_0_5152 (.A(n_8_0_6590), .B1(n_8_0_5456), .B2(n_8_0_390), 
      .ZN(n_8_0_4947));
   NAND2_X1 i_8_0_5153 (.A1(n_8_0_4950), .A2(n_8_0_4949), .ZN(n_8_0_4948));
   OAI211_X1 i_8_0_5154 (.A(n_8_0_5224), .B(n_8_0_6641), .C1(n_8_0_6795), 
      .C2(n_8_0_264), .ZN(n_8_0_4949));
   OAI21_X1 i_8_0_5155 (.A(n_8_0_6556), .B1(n_8_0_5460), .B2(n_8_0_264), 
      .ZN(n_8_0_4950));
   AOI21_X1 i_8_0_5156 (.A(n_8_0_6853), .B1(n_8_0_4951), .B2(n_8_0_4959), 
      .ZN(n_147));
   AND4_X1 i_8_0_5157 (.A1(n_8_0_4952), .A2(n_8_0_4967), .A3(n_8_0_4974), 
      .A4(n_8_0_4955), .ZN(n_8_0_4951));
   NOR4_X1 i_8_0_5158 (.A1(n_8_0_4964), .A2(n_8_0_4953), .A3(n_8_0_4954), 
      .A4(n_8_0_4970), .ZN(n_8_0_4952));
   OAI21_X1 i_8_0_5159 (.A(n_8_0_4961), .B1(n_8_0_6811), .B2(n_8_0_13), .ZN(
      n_8_0_4953));
   AOI221_X1 i_8_0_5160 (.A(n_8_0_7085), .B1(n_8_0_7084), .B2(n_8_0_5908), 
      .C1(n_8_0_6812), .C2(n_8_0_13), .ZN(n_8_0_4954));
   OAI21_X1 i_8_0_5161 (.A(n_8_0_4956), .B1(n_8_0_4957), .B2(n_8_0_6233), 
      .ZN(n_8_0_4955));
   NAND2_X1 i_8_0_5162 (.A1(n_8_0_4958), .A2(n_8_0_454), .ZN(n_8_0_4956));
   NOR2_X1 i_8_0_5163 (.A1(n_8_0_4958), .A2(n_8_0_454), .ZN(n_8_0_4957));
   OAI21_X1 i_8_0_5164 (.A(\out_bs[7] [6]), .B1(n_8_0_6541), .B2(n_8_0_5056), 
      .ZN(n_8_0_4958));
   OAI211_X1 i_8_0_5165 (.A(n_8_0_5394), .B(n_8_0_4960), .C1(n_8_0_5262), 
      .C2(n_8_0_5902), .ZN(n_8_0_4959));
   OAI211_X1 i_8_0_5166 (.A(n_8_0_6525), .B(n_8_0_76), .C1(n_8_0_6526), .C2(
      n_8_0_5901), .ZN(n_8_0_4960));
   OAI211_X1 i_8_0_5167 (.A(n_8_0_5427), .B(n_8_0_4962), .C1(n_8_0_5425), 
      .C2(n_8_0_5905), .ZN(n_8_0_4961));
   OAI21_X1 i_8_0_5168 (.A(n_8_0_139), .B1(n_8_0_6606), .B2(n_8_0_4963), 
      .ZN(n_8_0_4962));
   NOR2_X1 i_8_0_5169 (.A1(\out_bs[2] [5]), .A2(n_8_0_5905), .ZN(n_8_0_4963));
   OAI21_X1 i_8_0_5170 (.A(n_8_0_4965), .B1(n_8_0_6755), .B2(n_8_0_391), 
      .ZN(n_8_0_4964));
   OAI21_X1 i_8_0_5171 (.A(n_8_0_4966), .B1(n_8_0_5891), .B2(\out_bs[6] [5]), 
      .ZN(n_8_0_4965));
   AOI21_X1 i_8_0_5172 (.A(n_8_0_7012), .B1(n_8_0_6758), .B2(n_8_0_391), 
      .ZN(n_8_0_4966));
   OAI21_X1 i_8_0_5173 (.A(n_8_0_4968), .B1(n_8_0_6843), .B2(n_8_0_6932), 
      .ZN(n_8_0_4967));
   OAI21_X1 i_8_0_5174 (.A(n_8_0_4969), .B1(n_8_0_6837), .B2(n_8_0_202), 
      .ZN(n_8_0_4968));
   AOI21_X1 i_8_0_5175 (.A(n_8_0_6659), .B1(n_8_0_5917), .B2(\out_bs[3] [6]), 
      .ZN(n_8_0_4969));
   OAI21_X1 i_8_0_5176 (.A(n_8_0_4971), .B1(n_8_0_6824), .B2(n_8_0_328), 
      .ZN(n_8_0_4970));
   OAI211_X1 i_8_0_5177 (.A(n_8_0_4972), .B(\out_bs[5] [6]), .C1(n_8_0_6516), 
      .C2(n_8_0_5053), .ZN(n_8_0_4971));
   NAND2_X1 i_8_0_5178 (.A1(n_8_0_6619), .A2(n_8_0_328), .ZN(n_8_0_4972));
   INV_X1 i_8_0_5179 (.A(n_8_0_4974), .ZN(n_8_0_4973));
   OAI211_X1 i_8_0_5180 (.A(n_8_0_5459), .B(n_8_0_4975), .C1(n_8_0_5458), 
      .C2(n_8_0_5897), .ZN(n_8_0_4974));
   OAI21_X1 i_8_0_5181 (.A(n_8_0_265), .B1(n_8_0_6556), .B2(n_8_0_4976), 
      .ZN(n_8_0_4975));
   NOR2_X1 i_8_0_5182 (.A1(n_8_0_6559), .A2(n_8_0_5223), .ZN(n_8_0_4976));
   NOR2_X1 i_8_0_5183 (.A1(n_8_0_4977), .A2(n_8_0_6853), .ZN(n_148));
   NOR4_X1 i_8_0_5184 (.A1(n_8_0_4979), .A2(n_8_0_4978), .A3(n_8_0_4998), 
      .A4(n_8_0_4990), .ZN(n_8_0_4977));
   NAND3_X1 i_8_0_5185 (.A1(n_8_0_4981), .A2(n_8_0_4993), .A3(n_8_0_4995), 
      .ZN(n_8_0_4978));
   OAI211_X1 i_8_0_5186 (.A(n_8_0_4980), .B(n_8_0_5001), .C1(n_8_0_6811), 
      .C2(n_8_0_14), .ZN(n_8_0_4979));
   AOI211_X1 i_8_0_5187 (.A(n_8_0_4987), .B(n_8_0_4984), .C1(n_8_0_4985), 
      .C2(n_8_0_6731), .ZN(n_8_0_4980));
   OAI211_X1 i_8_0_5188 (.A(n_8_0_5427), .B(n_8_0_4982), .C1(n_8_0_5425), 
      .C2(n_8_0_5948), .ZN(n_8_0_4981));
   OAI21_X1 i_8_0_5189 (.A(n_8_0_140), .B1(n_8_0_6606), .B2(n_8_0_4983), 
      .ZN(n_8_0_4982));
   NOR2_X1 i_8_0_5190 (.A1(\out_bs[2] [5]), .A2(n_8_0_5948), .ZN(n_8_0_4983));
   NOR2_X1 i_8_0_5191 (.A1(n_8_0_455), .A2(n_8_0_4986), .ZN(n_8_0_4984));
   NAND2_X1 i_8_0_5192 (.A1(n_8_0_455), .A2(n_8_0_4986), .ZN(n_8_0_4985));
   AOI21_X1 i_8_0_5193 (.A(n_8_0_6728), .B1(n_8_0_5952), .B2(\out_bs[7] [6]), 
      .ZN(n_8_0_4986));
   AOI211_X1 i_8_0_5194 (.A(n_8_0_5395), .B(n_8_0_4988), .C1(n_8_0_77), .C2(
      n_8_0_6526), .ZN(n_8_0_4987));
   NOR2_X1 i_8_0_5195 (.A1(n_8_0_4989), .A2(\out_bs[1] [5]), .ZN(n_8_0_4988));
   OAI21_X1 i_8_0_5196 (.A(n_8_0_5961), .B1(n_8_0_6782), .B2(n_8_0_77), .ZN(
      n_8_0_4989));
   OAI21_X1 i_8_0_5197 (.A(n_8_0_4991), .B1(n_8_0_6824), .B2(n_8_0_329), 
      .ZN(n_8_0_4990));
   OAI211_X1 i_8_0_5198 (.A(n_8_0_4992), .B(\out_bs[5] [6]), .C1(n_8_0_6676), 
      .C2(n_8_0_5053), .ZN(n_8_0_4991));
   NAND2_X1 i_8_0_5199 (.A1(n_8_0_6619), .A2(n_8_0_329), .ZN(n_8_0_4992));
   OAI21_X1 i_8_0_5200 (.A(n_8_0_4994), .B1(n_8_0_6843), .B2(n_8_0_6931), 
      .ZN(n_8_0_4993));
   OAI221_X1 i_8_0_5201 (.A(n_8_0_6658), .B1(n_8_0_5932), .B2(n_8_0_7047), 
      .C1(n_8_0_6837), .C2(n_8_0_203), .ZN(n_8_0_4994));
   OAI21_X1 i_8_0_5202 (.A(n_8_0_4996), .B1(n_8_0_4997), .B2(n_8_0_6640), 
      .ZN(n_8_0_4995));
   OAI21_X1 i_8_0_5203 (.A(n_8_0_6556), .B1(n_8_0_5460), .B2(n_8_0_266), 
      .ZN(n_8_0_4996));
   OAI21_X1 i_8_0_5204 (.A(n_8_0_5224), .B1(n_8_0_6795), .B2(n_8_0_266), 
      .ZN(n_8_0_4997));
   AOI211_X1 i_8_0_5205 (.A(n_8_0_5456), .B(n_8_0_4999), .C1(n_8_0_392), 
      .C2(n_8_0_6590), .ZN(n_8_0_4998));
   NOR2_X1 i_8_0_5206 (.A1(n_8_0_5000), .A2(\out_bs[6] [5]), .ZN(n_8_0_4999));
   OAI21_X1 i_8_0_5207 (.A(n_8_0_5936), .B1(n_8_0_6755), .B2(n_8_0_392), 
      .ZN(n_8_0_5000));
   OAI211_X1 i_8_0_5208 (.A(n_8_0_5002), .B(\out_bs[0] [6]), .C1(\out_bs[0] [5]), 
      .C2(n_8_0_5940), .ZN(n_8_0_5001));
   NAND2_X1 i_8_0_5209 (.A1(n_8_0_6812), .A2(n_8_0_14), .ZN(n_8_0_5002));
   AOI21_X1 i_8_0_5210 (.A(n_8_0_6853), .B1(n_8_0_5020), .B2(n_8_0_5003), 
      .ZN(n_149));
   NOR4_X1 i_8_0_5211 (.A1(n_8_0_5017), .A2(n_8_0_5006), .A3(n_8_0_5004), 
      .A4(n_8_0_5014), .ZN(n_8_0_5003));
   AOI211_X1 i_8_0_5212 (.A(n_8_0_5395), .B(n_8_0_5005), .C1(n_8_0_78), .C2(
      n_8_0_6526), .ZN(n_8_0_5004));
   AOI211_X1 i_8_0_5213 (.A(\out_bs[1] [5]), .B(n_8_0_5979), .C1(n_8_0_6781), 
      .C2(n_8_0_6977), .ZN(n_8_0_5005));
   NAND2_X1 i_8_0_5214 (.A1(n_8_0_5012), .A2(n_8_0_5007), .ZN(n_8_0_5006));
   OAI21_X1 i_8_0_5215 (.A(n_8_0_5008), .B1(n_8_0_5009), .B2(n_8_0_6731), 
      .ZN(n_8_0_5007));
   NAND2_X1 i_8_0_5216 (.A1(n_8_0_5011), .A2(n_8_0_456), .ZN(n_8_0_5008));
   INV_X1 i_8_0_5217 (.A(n_8_0_5010), .ZN(n_8_0_5009));
   OR2_X1 i_8_0_5218 (.A1(n_8_0_5011), .A2(n_8_0_456), .ZN(n_8_0_5010));
   OAI21_X1 i_8_0_5219 (.A(\out_bs[7] [6]), .B1(n_8_0_5973), .B2(\out_bs[7] [5]), 
      .ZN(n_8_0_5011));
   AOI21_X1 i_8_0_5220 (.A(n_8_0_5013), .B1(n_8_0_6773), .B2(n_8_0_6959), 
      .ZN(n_8_0_5012));
   AOI221_X1 i_8_0_5221 (.A(n_8_0_7060), .B1(n_8_0_7059), .B2(n_8_0_5988), 
      .C1(n_8_0_6772), .C2(n_8_0_141), .ZN(n_8_0_5013));
   OAI21_X1 i_8_0_5222 (.A(n_8_0_5015), .B1(n_8_0_6824), .B2(n_8_0_330), 
      .ZN(n_8_0_5014));
   OAI211_X1 i_8_0_5223 (.A(n_8_0_5016), .B(\out_bs[5] [6]), .C1(n_8_0_6674), 
      .C2(n_8_0_5053), .ZN(n_8_0_5015));
   NAND2_X1 i_8_0_5224 (.A1(n_8_0_6619), .A2(n_8_0_330), .ZN(n_8_0_5016));
   OAI21_X1 i_8_0_5225 (.A(n_8_0_5018), .B1(n_8_0_6837), .B2(n_8_0_204), 
      .ZN(n_8_0_5017));
   OAI211_X1 i_8_0_5226 (.A(n_8_0_5019), .B(\out_bs[3] [6]), .C1(\out_bs[3] [5]), 
      .C2(n_8_0_6005), .ZN(n_8_0_5018));
   NAND2_X1 i_8_0_5227 (.A1(n_8_0_6844), .A2(n_8_0_204), .ZN(n_8_0_5019));
   NOR3_X1 i_8_0_5228 (.A1(n_8_0_5027), .A2(n_8_0_5024), .A3(n_8_0_5021), 
      .ZN(n_8_0_5020));
   AOI211_X1 i_8_0_5229 (.A(n_8_0_5460), .B(n_8_0_5022), .C1(n_8_0_267), 
      .C2(n_8_0_6556), .ZN(n_8_0_5021));
   NOR2_X1 i_8_0_5230 (.A1(n_8_0_5023), .A2(\out_bs[4] [5]), .ZN(n_8_0_5022));
   OAI21_X1 i_8_0_5231 (.A(n_8_0_5996), .B1(n_8_0_6795), .B2(n_8_0_267), 
      .ZN(n_8_0_5023));
   AOI22_X1 i_8_0_5232 (.A1(n_8_0_15), .A2(n_8_0_5026), .B1(n_8_0_5025), 
      .B2(n_8_0_6811), .ZN(n_8_0_5024));
   OAI21_X1 i_8_0_5233 (.A(\out_bs[0] [6]), .B1(n_8_0_5999), .B2(\out_bs[0] [5]), 
      .ZN(n_8_0_5025));
   OAI21_X1 i_8_0_5234 (.A(n_8_0_6250), .B1(n_8_0_5999), .B2(\out_bs[0] [5]), 
      .ZN(n_8_0_5026));
   AOI211_X1 i_8_0_5235 (.A(n_8_0_5456), .B(n_8_0_5028), .C1(n_8_0_393), 
      .C2(n_8_0_6590), .ZN(n_8_0_5027));
   NOR3_X1 i_8_0_5236 (.A1(\out_bs[6] [5]), .A2(n_8_0_5029), .A3(n_8_0_5969), 
      .ZN(n_8_0_5028));
   NOR2_X1 i_8_0_5237 (.A1(n_8_0_393), .A2(n_8_0_6755), .ZN(n_8_0_5029));
   AOI21_X1 i_8_0_5238 (.A(n_8_0_6853), .B1(n_8_0_5055), .B2(n_8_0_5030), 
      .ZN(n_150));
   NOR3_X1 i_8_0_5239 (.A1(n_8_0_5032), .A2(n_8_0_5031), .A3(n_8_0_5037), 
      .ZN(n_8_0_5030));
   OR4_X1 i_8_0_5240 (.A1(n_8_0_5058), .A2(n_8_0_5045), .A3(n_8_0_5039), 
      .A4(n_8_0_5034), .ZN(n_8_0_5031));
   NAND3_X1 i_8_0_5241 (.A1(n_8_0_5049), .A2(n_8_0_5048), .A3(n_8_0_5043), 
      .ZN(n_8_0_5032));
   INV_X1 i_8_0_5242 (.A(n_8_0_5034), .ZN(n_8_0_5033));
   OAI21_X1 i_8_0_5243 (.A(n_8_0_5035), .B1(n_8_0_6755), .B2(n_8_0_394), 
      .ZN(n_8_0_5034));
   OAI211_X1 i_8_0_5244 (.A(n_8_0_5036), .B(\out_bs[6] [6]), .C1(\out_bs[6] [5]), 
      .C2(\out_bs[6] [4]), .ZN(n_8_0_5035));
   NAND2_X1 i_8_0_5245 (.A1(n_8_0_6758), .A2(n_8_0_394), .ZN(n_8_0_5036));
   AOI21_X1 i_8_0_5246 (.A(n_8_0_16), .B1(n_8_0_6811), .B2(n_8_0_5038), .ZN(
      n_8_0_5037));
   OAI21_X1 i_8_0_5247 (.A(\out_bs[0] [6]), .B1(\out_bs[0] [5]), .B2(
      \out_bs[0] [4]), .ZN(n_8_0_5038));
   OAI22_X1 i_8_0_5248 (.A1(n_8_0_142), .A2(n_8_0_5040), .B1(n_8_0_6606), 
      .B2(n_8_0_5042), .ZN(n_8_0_5039));
   INV_X1 i_8_0_5249 (.A(n_8_0_5041), .ZN(n_8_0_5040));
   AOI21_X1 i_8_0_5250 (.A(n_8_0_5428), .B1(n_8_0_6772), .B2(n_8_0_5042), 
      .ZN(n_8_0_5041));
   NOR2_X1 i_8_0_5251 (.A1(\out_bs[2] [5]), .A2(\out_bs[2] [4]), .ZN(n_8_0_5042));
   OAI21_X1 i_8_0_5252 (.A(n_8_0_5044), .B1(n_8_0_6843), .B2(n_8_0_6930), 
      .ZN(n_8_0_5043));
   OAI211_X1 i_8_0_5253 (.A(n_8_0_6658), .B(n_8_0_6656), .C1(n_8_0_6837), 
      .C2(n_8_0_205), .ZN(n_8_0_5044));
   OAI21_X1 i_8_0_5254 (.A(n_8_0_5046), .B1(n_8_0_6782), .B2(n_8_0_79), .ZN(
      n_8_0_5045));
   OAI211_X1 i_8_0_5255 (.A(n_8_0_5047), .B(\out_bs[1] [6]), .C1(\out_bs[1] [5]), 
      .C2(\out_bs[1] [4]), .ZN(n_8_0_5046));
   NAND2_X1 i_8_0_5256 (.A1(n_8_0_6784), .A2(n_8_0_79), .ZN(n_8_0_5047));
   OAI21_X1 i_8_0_5257 (.A(n_8_0_6250), .B1(\out_bs[0] [4]), .B2(\out_bs[0] [5]), 
      .ZN(n_8_0_5048));
   INV_X1 i_8_0_5258 (.A(n_8_0_5050), .ZN(n_8_0_5049));
   OAI21_X1 i_8_0_5259 (.A(n_8_0_5051), .B1(n_8_0_6824), .B2(n_8_0_331), 
      .ZN(n_8_0_5050));
   NAND3_X1 i_8_0_5260 (.A1(n_8_0_5052), .A2(\out_bs[5] [6]), .A3(n_8_0_5053), 
      .ZN(n_8_0_5051));
   NAND2_X1 i_8_0_5261 (.A1(n_8_0_6824), .A2(n_8_0_331), .ZN(n_8_0_5052));
   NAND2_X1 i_8_0_5262 (.A1(n_8_0_7023), .A2(n_8_0_7022), .ZN(n_8_0_5053));
   NOR2_X1 i_8_0_5263 (.A1(\out_bs[5] [5]), .A2(\out_bs[5] [4]), .ZN(n_8_0_5054));
   AOI21_X1 i_8_0_5264 (.A(n_8_0_5057), .B1(n_8_0_5056), .B2(n_8_0_6466), 
      .ZN(n_8_0_5055));
   AOI21_X1 i_8_0_5266 (.A(n_8_0_457), .B1(n_8_0_6718), .B2(n_8_0_6716), 
      .ZN(n_8_0_5057));
   OAI22_X1 i_8_0_5267 (.A1(n_8_0_268), .A2(n_8_0_5221), .B1(n_8_0_5224), 
      .B2(n_8_0_6556), .ZN(n_8_0_5058));
   NOR2_X1 i_8_0_5276 (.A1(n_8_0_6031), .A2(n_8_0_5928), .ZN(n_8_0_5066));
   NOR2_X1 i_8_0_5277 (.A1(n_8_0_6555), .A2(n_8_0_6031), .ZN(n_8_0_5067));
   OAI221_X1 i_8_0_5279 (.A(n_8_0_6511), .B1(n_8_0_6057), .B2(n_8_0_6513), 
      .C1(n_8_0_5070), .C2(n_8_0_332), .ZN(n_8_0_5069));
   AOI21_X1 i_8_0_5280 (.A(n_8_0_6375), .B1(n_8_0_6059), .B2(n_8_0_6686), 
      .ZN(n_8_0_5070));
   OAI211_X1 i_8_0_5282 (.A(n_8_0_5073), .B(\out_bs[6] [6]), .C1(\out_bs[6] [5]), 
      .C2(n_8_0_6035), .ZN(n_8_0_5072));
   NAND2_X1 i_8_0_5283 (.A1(n_8_0_6758), .A2(n_8_0_395), .ZN(n_8_0_5073));
   OAI21_X1 i_8_0_5285 (.A(n_8_0_6526), .B1(n_8_0_5395), .B2(n_8_0_80), .ZN(
      n_8_0_5075));
   OAI211_X1 i_8_0_5286 (.A(n_8_0_7071), .B(n_8_0_6049), .C1(n_8_0_6782), 
      .C2(n_8_0_80), .ZN(n_8_0_5076));
   AOI21_X1 i_8_0_5288 (.A(n_8_0_5428), .B1(n_8_0_5426), .B2(n_8_0_6046), 
      .ZN(n_8_0_5078));
   OAI21_X1 i_8_0_5289 (.A(n_8_0_143), .B1(n_8_0_6606), .B2(n_8_0_6046), 
      .ZN(n_8_0_5079));
   INV_X1 i_8_0_5290 (.A(n_8_0_5081), .ZN(n_8_0_5080));
   AOI21_X1 i_8_0_5293 (.A(n_8_0_6844), .B1(n_8_0_6658), .B2(n_8_0_5085), 
      .ZN(n_8_0_5083));
   AOI21_X1 i_8_0_5294 (.A(n_8_0_206), .B1(n_8_0_6572), .B2(n_8_0_5085), 
      .ZN(n_8_0_5084));
   NAND2_X1 i_8_0_5295 (.A1(n_8_0_5086), .A2(n_8_0_6657), .ZN(n_8_0_5085));
   INV_X1 i_8_0_5296 (.A(n_8_0_5087), .ZN(n_8_0_5086));
   NOR2_X1 i_8_0_5297 (.A1(n_8_0_6357), .A2(\out_bs[3] [3]), .ZN(n_8_0_5087));
   NOR2_X1 i_8_0_5298 (.A1(n_8_0_5088), .A2(n_8_0_6853), .ZN(n_151));
   NOR2_X1 i_8_0_5299 (.A1(n_8_0_5103), .A2(n_8_0_5089), .ZN(n_8_0_5088));
   NAND4_X1 i_8_0_5300 (.A1(n_8_0_5112), .A2(n_8_0_5091), .A3(n_8_0_5090), 
      .A4(n_8_0_5095), .ZN(n_8_0_5089));
   AOI21_X1 i_8_0_5301 (.A(n_8_0_5109), .B1(n_8_0_5092), .B2(n_8_0_6233), 
      .ZN(n_8_0_5090));
   NOR4_X1 i_8_0_5302 (.A1(n_8_0_5106), .A2(n_8_0_5101), .A3(n_8_0_5099), 
      .A4(n_8_0_5093), .ZN(n_8_0_5091));
   NAND2_X1 i_8_0_5303 (.A1(n_8_0_459), .A2(n_8_0_5094), .ZN(n_8_0_5092));
   NOR2_X1 i_8_0_5304 (.A1(n_8_0_459), .A2(n_8_0_5094), .ZN(n_8_0_5093));
   AOI21_X1 i_8_0_5305 (.A(n_8_0_6728), .B1(n_8_0_6080), .B2(n_8_0_6717), 
      .ZN(n_8_0_5094));
   INV_X1 i_8_0_5306 (.A(n_8_0_5096), .ZN(n_8_0_5095));
   OAI21_X1 i_8_0_5307 (.A(n_8_0_5097), .B1(n_8_0_6772), .B2(n_8_0_144), 
      .ZN(n_8_0_5096));
   OAI211_X1 i_8_0_5308 (.A(n_8_0_5098), .B(\out_bs[2] [6]), .C1(\out_bs[2] [5]), 
      .C2(n_8_0_6069), .ZN(n_8_0_5097));
   NAND2_X1 i_8_0_5309 (.A1(n_8_0_6772), .A2(n_8_0_144), .ZN(n_8_0_5098));
   AOI21_X1 i_8_0_5310 (.A(n_8_0_5100), .B1(n_8_0_6812), .B2(n_8_0_18), .ZN(
      n_8_0_5099));
   AOI221_X1 i_8_0_5311 (.A(n_8_0_6671), .B1(\out_bs[0] [6]), .B2(n_8_0_6082), 
      .C1(n_8_0_6810), .C2(n_8_0_6986), .ZN(n_8_0_5100));
   AOI221_X1 i_8_0_5312 (.A(n_8_0_5456), .B1(n_8_0_5452), .B2(n_8_0_6086), 
      .C1(n_8_0_5102), .C2(n_8_0_396), .ZN(n_8_0_5101));
   OAI21_X1 i_8_0_5313 (.A(n_8_0_6591), .B1(n_8_0_6087), .B2(\out_bs[6] [5]), 
      .ZN(n_8_0_5102));
   OAI211_X1 i_8_0_5314 (.A(n_8_0_6511), .B(n_8_0_5104), .C1(n_8_0_6376), 
      .C2(n_8_0_333), .ZN(n_8_0_5103));
   NAND3_X1 i_8_0_5315 (.A1(n_8_0_5105), .A2(n_8_0_6686), .A3(n_8_0_6097), 
      .ZN(n_8_0_5104));
   NAND2_X1 i_8_0_5316 (.A1(n_8_0_6619), .A2(n_8_0_333), .ZN(n_8_0_5105));
   OAI33_X1 i_8_0_5317 (.A1(n_8_0_270), .A2(n_8_0_5221), .A3(n_8_0_5107), 
      .B1(n_8_0_5108), .B2(n_8_0_6556), .B3(n_8_0_5224), .ZN(n_8_0_5106));
   NOR2_X1 i_8_0_5318 (.A1(n_8_0_6092), .A2(n_8_0_5928), .ZN(n_8_0_5107));
   NOR2_X1 i_8_0_5319 (.A1(n_8_0_6092), .A2(n_8_0_6636), .ZN(n_8_0_5108));
   INV_X1 i_8_0_5320 (.A(n_8_0_5110), .ZN(n_8_0_5109));
   OAI211_X1 i_8_0_5321 (.A(n_8_0_5394), .B(n_8_0_5111), .C1(n_8_0_5262), 
      .C2(n_8_0_6074), .ZN(n_8_0_5110));
   OAI211_X1 i_8_0_5322 (.A(n_8_0_81), .B(n_8_0_6525), .C1(n_8_0_6526), .C2(
      n_8_0_6075), .ZN(n_8_0_5111));
   AOI211_X1 i_8_0_5323 (.A(n_8_0_6576), .B(n_8_0_5113), .C1(n_8_0_5116), 
      .C2(n_8_0_5226), .ZN(n_8_0_5112));
   AOI21_X1 i_8_0_5324 (.A(n_8_0_207), .B1(n_8_0_6572), .B2(n_8_0_5114), 
      .ZN(n_8_0_5113));
   NAND2_X1 i_8_0_5325 (.A1(n_8_0_5116), .A2(n_8_0_6657), .ZN(n_8_0_5114));
   INV_X1 i_8_0_5326 (.A(n_8_0_5116), .ZN(n_8_0_5115));
   NAND2_X1 i_8_0_5327 (.A1(n_8_0_6414), .A2(n_8_0_7044), .ZN(n_8_0_5116));
   AOI21_X1 i_8_0_5328 (.A(n_8_0_6853), .B1(n_8_0_5141), .B2(n_8_0_5117), 
      .ZN(n_152));
   NOR4_X1 i_8_0_5329 (.A1(n_8_0_5120), .A2(n_8_0_5118), .A3(n_8_0_5119), 
      .A4(n_8_0_5132), .ZN(n_8_0_5117));
   NAND3_X1 i_8_0_5330 (.A1(n_8_0_5138), .A2(n_8_0_5126), .A3(n_8_0_5123), 
      .ZN(n_8_0_5118));
   AOI21_X1 i_8_0_5331 (.A(n_8_0_19), .B1(n_8_0_6595), .B2(n_8_0_5131), .ZN(
      n_8_0_5119));
   NAND3_X1 i_8_0_5332 (.A1(n_8_0_5129), .A2(n_8_0_5122), .A3(n_8_0_5121), 
      .ZN(n_8_0_5120));
   OAI21_X1 i_8_0_5333 (.A(n_8_0_5136), .B1(n_8_0_5135), .B2(n_8_0_6233), 
      .ZN(n_8_0_5121));
   OAI21_X1 i_8_0_5334 (.A(n_8_0_6250), .B1(n_8_0_6140), .B2(\out_bs[0] [5]), 
      .ZN(n_8_0_5122));
   NOR3_X1 i_8_0_5335 (.A1(n_8_0_5152), .A2(n_8_0_5125), .A3(n_8_0_5124), 
      .ZN(n_8_0_5123));
   AOI211_X1 i_8_0_5336 (.A(n_8_0_271), .B(n_8_0_5221), .C1(n_8_0_5929), 
      .C2(n_8_0_6114), .ZN(n_8_0_5124));
   NOR3_X1 i_8_0_5337 (.A1(n_8_0_6639), .A2(n_8_0_6556), .A3(n_8_0_5224), 
      .ZN(n_8_0_5125));
   OAI21_X1 i_8_0_5338 (.A(n_8_0_5127), .B1(n_8_0_5128), .B2(n_8_0_6589), 
      .ZN(n_8_0_5126));
   AOI21_X1 i_8_0_5339 (.A(n_8_0_5456), .B1(n_8_0_5452), .B2(n_8_0_6123), 
      .ZN(n_8_0_5127));
   OAI21_X1 i_8_0_5340 (.A(n_8_0_397), .B1(n_8_0_6590), .B2(n_8_0_6123), 
      .ZN(n_8_0_5128));
   OAI211_X1 i_8_0_5341 (.A(n_8_0_5394), .B(n_8_0_5130), .C1(n_8_0_5262), 
      .C2(n_8_0_6127), .ZN(n_8_0_5129));
   OAI211_X1 i_8_0_5342 (.A(n_8_0_6525), .B(n_8_0_82), .C1(n_8_0_6526), .C2(
      n_8_0_6126), .ZN(n_8_0_5130));
   NAND2_X1 i_8_0_5343 (.A1(n_8_0_6140), .A2(\out_bs[0] [6]), .ZN(n_8_0_5131));
   AOI211_X1 i_8_0_5344 (.A(n_8_0_5428), .B(n_8_0_5134), .C1(n_8_0_5133), 
      .C2(n_8_0_145), .ZN(n_8_0_5132));
   OAI21_X1 i_8_0_5345 (.A(n_8_0_6607), .B1(n_8_0_6131), .B2(\out_bs[2] [5]), 
      .ZN(n_8_0_5133));
   NOR2_X1 i_8_0_5346 (.A1(n_8_0_6131), .A2(n_8_0_5425), .ZN(n_8_0_5134));
   NOR2_X1 i_8_0_5347 (.A1(n_8_0_460), .A2(n_8_0_5137), .ZN(n_8_0_5135));
   NAND2_X1 i_8_0_5348 (.A1(n_8_0_460), .A2(n_8_0_5137), .ZN(n_8_0_5136));
   AOI21_X1 i_8_0_5349 (.A(n_8_0_6728), .B1(n_8_0_6118), .B2(n_8_0_6717), 
      .ZN(n_8_0_5137));
   NOR2_X1 i_8_0_5350 (.A1(n_8_0_5139), .A2(n_8_0_6512), .ZN(n_8_0_5138));
   OAI22_X1 i_8_0_5351 (.A1(n_8_0_334), .A2(n_8_0_5140), .B1(n_8_0_5470), 
      .B2(n_8_0_6135), .ZN(n_8_0_5139));
   AOI21_X1 i_8_0_5352 (.A(n_8_0_6375), .B1(n_8_0_6136), .B2(n_8_0_6686), 
      .ZN(n_8_0_5140));
   AOI21_X1 i_8_0_5353 (.A(n_8_0_5142), .B1(n_8_0_5143), .B2(n_8_0_6657), 
      .ZN(n_8_0_5141));
   OAI21_X1 i_8_0_5354 (.A(n_8_0_6575), .B1(n_8_0_6572), .B2(n_8_0_208), 
      .ZN(n_8_0_5142));
   AOI21_X1 i_8_0_5355 (.A(n_8_0_6109), .B1(n_8_0_6844), .B2(n_8_0_208), 
      .ZN(n_8_0_5143));
   AOI21_X1 i_8_0_5356 (.A(n_8_0_6853), .B1(n_8_0_5150), .B2(n_8_0_5144), 
      .ZN(n_153));
   NOR4_X1 i_8_0_5357 (.A1(n_8_0_5164), .A2(n_8_0_5145), .A3(n_8_0_5160), 
      .A4(n_8_0_5157), .ZN(n_8_0_5144));
   OAI211_X1 i_8_0_5358 (.A(n_8_0_5146), .B(n_8_0_5154), .C1(n_8_0_6595), 
      .C2(n_8_0_20), .ZN(n_8_0_5145));
   NOR4_X1 i_8_0_5359 (.A1(n_8_0_5162), .A2(n_8_0_5149), .A3(n_8_0_5148), 
      .A4(n_8_0_5168), .ZN(n_8_0_5146));
   NOR2_X1 i_8_0_5360 (.A1(n_8_0_5148), .A2(n_8_0_5149), .ZN(n_8_0_5147));
   OAI21_X1 i_8_0_5361 (.A(n_8_0_6575), .B1(n_8_0_6572), .B2(n_8_0_209), 
      .ZN(n_8_0_5148));
   AOI211_X1 i_8_0_5362 (.A(n_8_0_6656), .B(n_8_0_6161), .C1(n_8_0_6844), 
      .C2(n_8_0_209), .ZN(n_8_0_5149));
   NOR2_X1 i_8_0_5363 (.A1(n_8_0_5152), .A2(n_8_0_5151), .ZN(n_8_0_5150));
   AOI211_X1 i_8_0_5364 (.A(n_8_0_272), .B(n_8_0_5221), .C1(n_8_0_5929), 
      .C2(n_8_0_6171), .ZN(n_8_0_5151));
   AOI211_X1 i_8_0_5365 (.A(n_8_0_5224), .B(n_8_0_6556), .C1(n_8_0_7034), 
      .C2(n_8_0_6171), .ZN(n_8_0_5152));
   INV_X1 i_8_0_5366 (.A(n_8_0_5154), .ZN(n_8_0_5153));
   NAND3_X1 i_8_0_5367 (.A1(n_8_0_5455), .A2(n_8_0_5156), .A3(n_8_0_5155), 
      .ZN(n_8_0_5154));
   OAI211_X1 i_8_0_5368 (.A(n_8_0_7011), .B(n_8_0_6293), .C1(n_8_0_6755), 
      .C2(n_8_0_398), .ZN(n_8_0_5155));
   NAND2_X1 i_8_0_5369 (.A1(n_8_0_6590), .A2(n_8_0_398), .ZN(n_8_0_5156));
   OAI211_X1 i_8_0_5370 (.A(n_8_0_6511), .B(n_8_0_5158), .C1(n_8_0_6376), 
      .C2(n_8_0_335), .ZN(n_8_0_5157));
   NAND3_X1 i_8_0_5371 (.A1(n_8_0_5159), .A2(n_8_0_6686), .A3(n_8_0_6165), 
      .ZN(n_8_0_5158));
   NAND2_X1 i_8_0_5372 (.A1(n_8_0_6619), .A2(n_8_0_335), .ZN(n_8_0_5159));
   AOI22_X1 i_8_0_5373 (.A1(n_8_0_6247), .A2(n_8_0_5161), .B1(n_8_0_6812), 
      .B2(n_8_0_20), .ZN(n_8_0_5160));
   NAND3_X1 i_8_0_5374 (.A1(n_8_0_6175), .A2(\out_bs[0] [4]), .A3(\out_bs[0] [6]), 
      .ZN(n_8_0_5161));
   AOI221_X1 i_8_0_5375 (.A(n_8_0_5428), .B1(n_8_0_5426), .B2(n_8_0_6151), 
      .C1(n_8_0_5163), .C2(n_8_0_146), .ZN(n_8_0_5162));
   OAI21_X1 i_8_0_5376 (.A(n_8_0_6607), .B1(n_8_0_6150), .B2(\out_bs[2] [5]), 
      .ZN(n_8_0_5163));
   AOI21_X1 i_8_0_5377 (.A(n_8_0_5165), .B1(n_8_0_5166), .B2(n_8_0_6232), 
      .ZN(n_8_0_5164));
   NOR2_X1 i_8_0_5378 (.A1(n_8_0_6873), .A2(n_8_0_5167), .ZN(n_8_0_5165));
   NAND2_X1 i_8_0_5379 (.A1(n_8_0_6873), .A2(n_8_0_5167), .ZN(n_8_0_5166));
   OAI21_X1 i_8_0_5380 (.A(n_8_0_6727), .B1(n_8_0_6157), .B2(n_8_0_6716), 
      .ZN(n_8_0_5167));
   AOI21_X1 i_8_0_5381 (.A(n_8_0_5169), .B1(n_8_0_6526), .B2(n_8_0_83), .ZN(
      n_8_0_5168));
   OAI21_X1 i_8_0_5382 (.A(n_8_0_5394), .B1(n_8_0_5170), .B2(\out_bs[1] [5]), 
      .ZN(n_8_0_5169));
   OAI21_X1 i_8_0_5383 (.A(n_8_0_6147), .B1(n_8_0_6782), .B2(n_8_0_83), .ZN(
      n_8_0_5170));
   AOI21_X1 i_8_0_5391 (.A(n_8_0_6375), .B1(n_8_0_6210), .B2(n_8_0_6686), 
      .ZN(n_8_0_5177));
   OAI21_X1 i_8_0_5393 (.A(n_8_0_5180), .B1(n_8_0_6215), .B2(\out_bs[3] [5]), 
      .ZN(n_8_0_5179));
   AOI22_X1 i_8_0_5394 (.A1(n_8_0_6844), .A2(n_8_0_210), .B1(n_8_0_6656), 
      .B2(n_8_0_6658), .ZN(n_8_0_5180));
   INV_X1 i_8_0_5395 (.A(n_8_0_5182), .ZN(n_8_0_5181));
   NOR2_X1 i_8_0_5397 (.A1(n_8_0_5185), .A2(n_8_0_7012), .ZN(n_8_0_5183));
   OAI21_X1 i_8_0_5398 (.A(n_8_0_399), .B1(n_8_0_6590), .B2(n_8_0_5185), 
      .ZN(n_8_0_5184));
   NOR2_X1 i_8_0_5399 (.A1(\out_bs[6] [5]), .A2(n_8_0_6197), .ZN(n_8_0_5185));
   OAI21_X1 i_8_0_5401 (.A(n_8_0_6607), .B1(n_8_0_6181), .B2(\out_bs[2] [5]), 
      .ZN(n_8_0_5187));
   OAI21_X1 i_8_0_5403 (.A(n_8_0_6526), .B1(n_8_0_5395), .B2(n_8_0_84), .ZN(
      n_8_0_5189));
   OAI21_X1 i_8_0_5404 (.A(n_8_0_6206), .B1(n_8_0_6782), .B2(n_8_0_84), .ZN(
      n_8_0_5190));
   NOR2_X1 i_8_0_5405 (.A1(n_8_0_6185), .A2(\out_bs[0] [5]), .ZN(n_8_0_5191));
   AOI21_X1 i_8_0_5408 (.A(n_8_0_6728), .B1(n_8_0_6201), .B2(n_8_0_6717), 
      .ZN(n_8_0_5194));
   NOR2_X1 i_8_0_5410 (.A1(n_8_0_6191), .A2(n_8_0_5928), .ZN(n_8_0_5196));
   NOR2_X1 i_8_0_5411 (.A1(n_8_0_6191), .A2(n_8_0_6636), .ZN(n_8_0_5197));
   AOI21_X1 i_8_0_5412 (.A(n_8_0_6853), .B1(n_8_0_5206), .B2(n_8_0_5198), 
      .ZN(n_154));
   AOI211_X1 i_8_0_5413 (.A(n_8_0_5200), .B(n_8_0_5199), .C1(n_8_0_6233), 
      .C2(n_8_0_5217), .ZN(n_8_0_5198));
   NAND2_X1 i_8_0_5414 (.A1(n_8_0_5225), .A2(n_8_0_5209), .ZN(n_8_0_5199));
   NAND3_X1 i_8_0_5415 (.A1(n_8_0_5212), .A2(n_8_0_5201), .A3(n_8_0_5204), 
      .ZN(n_8_0_5200));
   NOR3_X1 i_8_0_5416 (.A1(n_8_0_5219), .A2(n_8_0_5216), .A3(n_8_0_5202), 
      .ZN(n_8_0_5201));
   OAI21_X1 i_8_0_5417 (.A(n_8_0_5203), .B1(n_8_0_6595), .B2(n_8_0_22), .ZN(
      n_8_0_5202));
   AOI21_X1 i_8_0_5418 (.A(n_8_0_6248), .B1(n_8_0_5218), .B2(\out_bs[0] [6]), 
      .ZN(n_8_0_5203));
   OAI211_X1 i_8_0_5419 (.A(n_8_0_5455), .B(n_8_0_5205), .C1(n_8_0_5451), 
      .C2(n_8_0_6225), .ZN(n_8_0_5204));
   OAI211_X1 i_8_0_5420 (.A(n_8_0_400), .B(n_8_0_6588), .C1(n_8_0_6590), 
      .C2(n_8_0_6226), .ZN(n_8_0_5205));
   NOR2_X1 i_8_0_5421 (.A1(n_8_0_5207), .A2(n_8_0_6512), .ZN(n_8_0_5206));
   OAI22_X1 i_8_0_5422 (.A1(n_8_0_337), .A2(n_8_0_5208), .B1(n_8_0_5470), 
      .B2(n_8_0_6301), .ZN(n_8_0_5207));
   AOI21_X1 i_8_0_5423 (.A(n_8_0_6375), .B1(n_8_0_6300), .B2(n_8_0_6686), 
      .ZN(n_8_0_5208));
   OAI211_X1 i_8_0_5424 (.A(n_8_0_5394), .B(n_8_0_5210), .C1(n_8_0_5262), 
      .C2(n_8_0_6271), .ZN(n_8_0_5209));
   OAI21_X1 i_8_0_5425 (.A(n_8_0_85), .B1(n_8_0_6526), .B2(n_8_0_5211), .ZN(
      n_8_0_5210));
   NOR2_X1 i_8_0_5426 (.A1(\out_bs[1] [5]), .A2(n_8_0_6271), .ZN(n_8_0_5211));
   INV_X1 i_8_0_5427 (.A(n_8_0_5213), .ZN(n_8_0_5212));
   OAI21_X1 i_8_0_5428 (.A(n_8_0_5214), .B1(n_8_0_6772), .B2(n_8_0_148), 
      .ZN(n_8_0_5213));
   OAI211_X1 i_8_0_5429 (.A(n_8_0_5215), .B(\out_bs[2] [6]), .C1(\out_bs[2] [5]), 
      .C2(n_8_0_6288), .ZN(n_8_0_5214));
   NAND2_X1 i_8_0_5430 (.A1(n_8_0_6772), .A2(n_8_0_148), .ZN(n_8_0_5215));
   AOI21_X1 i_8_0_5431 (.A(n_8_0_463), .B1(n_8_0_6727), .B2(n_8_0_6236), 
      .ZN(n_8_0_5216));
   NAND3_X1 i_8_0_5432 (.A1(n_8_0_6236), .A2(n_8_0_463), .A3(n_8_0_6727), 
      .ZN(n_8_0_5217));
   AOI21_X1 i_8_0_5433 (.A(n_8_0_6252), .B1(n_8_0_6812), .B2(n_8_0_22), .ZN(
      n_8_0_5218));
   OAI33_X1 i_8_0_5434 (.A1(n_8_0_274), .A2(n_8_0_5221), .A3(n_8_0_5220), 
      .B1(n_8_0_6556), .B2(n_8_0_5224), .B3(n_8_0_5222), .ZN(n_8_0_5219));
   NOR2_X1 i_8_0_5435 (.A1(n_8_0_6244), .A2(n_8_0_5928), .ZN(n_8_0_5220));
   AOI21_X1 i_8_0_5436 (.A(n_8_0_6794), .B1(n_8_0_5223), .B2(\out_bs[4] [6]), 
      .ZN(n_8_0_5221));
   NOR2_X1 i_8_0_5437 (.A1(n_8_0_6244), .A2(n_8_0_6636), .ZN(n_8_0_5222));
   NAND2_X1 i_8_0_5438 (.A1(n_8_0_7034), .A2(n_8_0_7033), .ZN(n_8_0_5223));
   NOR2_X1 i_8_0_5439 (.A1(\out_bs[4] [5]), .A2(\out_bs[4] [4]), .ZN(n_8_0_5224));
   AOI221_X1 i_8_0_5440 (.A(n_8_0_6576), .B1(n_8_0_6217), .B2(n_8_0_5226), 
      .C1(n_8_0_5227), .C2(n_8_0_6929), .ZN(n_8_0_5225));
   NOR2_X1 i_8_0_5441 (.A1(n_8_0_7045), .A2(n_8_0_6577), .ZN(n_8_0_5226));
   OAI21_X1 i_8_0_5442 (.A(n_8_0_6572), .B1(n_8_0_6218), .B2(n_8_0_6656), 
      .ZN(n_8_0_5227));
   AOI21_X1 i_8_0_5443 (.A(n_8_0_6853), .B1(n_8_0_5230), .B2(n_8_0_5228), 
      .ZN(n_155));
   NOR2_X1 i_8_0_5444 (.A1(n_8_0_5236), .A2(n_8_0_5229), .ZN(n_8_0_5228));
   NAND4_X1 i_8_0_5445 (.A1(n_8_0_5247), .A2(n_8_0_5242), .A3(n_8_0_5231), 
      .A4(n_8_0_5244), .ZN(n_8_0_5229));
   NOR3_X1 i_8_0_5446 (.A1(n_8_0_5234), .A2(n_8_0_5239), .A3(n_8_0_5250), 
      .ZN(n_8_0_5230));
   OAI21_X1 i_8_0_5447 (.A(n_8_0_5232), .B1(n_8_0_5233), .B2(\out_bs[0] [5]), 
      .ZN(n_8_0_5231));
   OAI21_X1 i_8_0_5448 (.A(n_8_0_6249), .B1(n_8_0_5274), .B2(n_8_0_23), .ZN(
      n_8_0_5232));
   OAI21_X1 i_8_0_5449 (.A(n_8_0_6261), .B1(n_8_0_6811), .B2(n_8_0_23), .ZN(
      n_8_0_5233));
   OAI221_X1 i_8_0_5450 (.A(n_8_0_6511), .B1(n_8_0_6298), .B2(n_8_0_5470), 
      .C1(n_8_0_5235), .C2(n_8_0_338), .ZN(n_8_0_5234));
   AOI21_X1 i_8_0_5451 (.A(n_8_0_6375), .B1(n_8_0_6299), .B2(n_8_0_6686), 
      .ZN(n_8_0_5235));
   OAI211_X1 i_8_0_5452 (.A(n_8_0_6575), .B(n_8_0_5237), .C1(n_8_0_6572), 
      .C2(n_8_0_212), .ZN(n_8_0_5236));
   NAND2_X1 i_8_0_5453 (.A1(n_8_0_6657), .A2(n_8_0_5238), .ZN(n_8_0_5237));
   AOI21_X1 i_8_0_5454 (.A(n_8_0_5698), .B1(n_8_0_6844), .B2(n_8_0_212), 
      .ZN(n_8_0_5238));
   INV_X1 i_8_0_5455 (.A(n_8_0_5240), .ZN(n_8_0_5239));
   OAI211_X1 i_8_0_5456 (.A(n_8_0_5455), .B(n_8_0_5241), .C1(n_8_0_5451), 
      .C2(n_8_0_6291), .ZN(n_8_0_5240));
   OAI211_X1 i_8_0_5457 (.A(n_8_0_401), .B(n_8_0_6588), .C1(n_8_0_6590), 
      .C2(n_8_0_6292), .ZN(n_8_0_5241));
   AOI21_X1 i_8_0_5458 (.A(n_8_0_5243), .B1(n_8_0_6773), .B2(n_8_0_6958), 
      .ZN(n_8_0_5242));
   AOI221_X1 i_8_0_5459 (.A(n_8_0_7060), .B1(n_8_0_7059), .B2(n_8_0_6286), 
      .C1(n_8_0_6772), .C2(n_8_0_149), .ZN(n_8_0_5243));
   OAI21_X1 i_8_0_5460 (.A(n_8_0_5245), .B1(n_8_0_5262), .B2(n_8_0_6268), 
      .ZN(n_8_0_5244));
   AOI21_X1 i_8_0_5461 (.A(n_8_0_5395), .B1(n_8_0_5246), .B2(n_8_0_86), .ZN(
      n_8_0_5245));
   OAI21_X1 i_8_0_5462 (.A(n_8_0_6527), .B1(n_8_0_6268), .B2(\out_bs[1] [5]), 
      .ZN(n_8_0_5246));
   OAI21_X1 i_8_0_5463 (.A(n_8_0_5249), .B1(n_8_0_5248), .B2(n_8_0_6728), 
      .ZN(n_8_0_5247));
   OAI22_X1 i_8_0_5464 (.A1(n_8_0_464), .A2(n_8_0_6730), .B1(n_8_0_6716), 
      .B2(n_8_0_6279), .ZN(n_8_0_5248));
   NAND2_X1 i_8_0_5465 (.A1(n_8_0_464), .A2(n_8_0_6730), .ZN(n_8_0_5249));
   AOI22_X1 i_8_0_5466 (.A1(n_8_0_275), .A2(n_8_0_5252), .B1(n_8_0_6795), 
      .B2(n_8_0_5251), .ZN(n_8_0_5250));
   OAI21_X1 i_8_0_5467 (.A(\out_bs[4] [6]), .B1(n_8_0_6275), .B2(\out_bs[4] [5]), 
      .ZN(n_8_0_5251));
   OAI21_X1 i_8_0_5468 (.A(n_8_0_6557), .B1(n_8_0_6275), .B2(\out_bs[4] [5]), 
      .ZN(n_8_0_5252));
   AOI21_X1 i_8_0_5469 (.A(n_8_0_6853), .B1(n_8_0_5255), .B2(n_8_0_5253), 
      .ZN(n_156));
   NOR3_X1 i_8_0_5470 (.A1(n_8_0_5256), .A2(n_8_0_5254), .A3(n_8_0_5261), 
      .ZN(n_8_0_5253));
   NAND2_X1 i_8_0_5471 (.A1(n_8_0_5270), .A2(n_8_0_5268), .ZN(n_8_0_5254));
   AOI211_X1 i_8_0_5472 (.A(n_8_0_5276), .B(n_8_0_5265), .C1(n_8_0_5273), 
      .C2(n_8_0_5275), .ZN(n_8_0_5255));
   NAND2_X1 i_8_0_5473 (.A1(n_8_0_5259), .A2(n_8_0_5257), .ZN(n_8_0_5256));
   OAI211_X1 i_8_0_5474 (.A(n_8_0_5427), .B(n_8_0_5258), .C1(n_8_0_5425), 
      .C2(n_8_0_6709), .ZN(n_8_0_5257));
   OAI211_X1 i_8_0_5475 (.A(n_8_0_150), .B(n_8_0_6604), .C1(n_8_0_6606), 
      .C2(n_8_0_6708), .ZN(n_8_0_5258));
   OAI21_X1 i_8_0_5476 (.A(n_8_0_5260), .B1(n_8_0_5481), .B2(n_8_0_6731), 
      .ZN(n_8_0_5259));
   OAI21_X1 i_8_0_5477 (.A(n_8_0_465), .B1(n_8_0_6232), .B2(n_8_0_5482), 
      .ZN(n_8_0_5260));
   AOI221_X1 i_8_0_5478 (.A(n_8_0_5395), .B1(n_8_0_5263), .B2(n_8_0_6695), 
      .C1(n_8_0_5264), .C2(n_8_0_87), .ZN(n_8_0_5261));
   NAND2_X1 i_8_0_5479 (.A1(n_8_0_6782), .A2(n_8_0_7071), .ZN(n_8_0_5262));
   NOR2_X1 i_8_0_5480 (.A1(n_8_0_6781), .A2(\out_bs[1] [5]), .ZN(n_8_0_5263));
   OAI21_X1 i_8_0_5481 (.A(n_8_0_6527), .B1(n_8_0_6696), .B2(\out_bs[1] [5]), 
      .ZN(n_8_0_5264));
   AOI211_X1 i_8_0_5482 (.A(n_8_0_5302), .B(n_8_0_5266), .C1(n_8_0_339), 
      .C2(n_8_0_6513), .ZN(n_8_0_5265));
   AOI21_X1 i_8_0_5483 (.A(n_8_0_5267), .B1(\out_bs[5] [3]), .B2(\out_bs[5] [4]), 
      .ZN(n_8_0_5266));
   OAI21_X1 i_8_0_5484 (.A(n_8_0_7023), .B1(n_8_0_6824), .B2(n_8_0_339), 
      .ZN(n_8_0_5267));
   AOI21_X1 i_8_0_5485 (.A(n_8_0_5269), .B1(n_8_0_6838), .B2(n_8_0_6928), 
      .ZN(n_8_0_5268));
   AOI221_X1 i_8_0_5486 (.A(n_8_0_7047), .B1(n_8_0_7046), .B2(n_8_0_6647), 
      .C1(n_8_0_6844), .C2(n_8_0_213), .ZN(n_8_0_5269));
   OAI21_X1 i_8_0_5487 (.A(n_8_0_5271), .B1(n_8_0_5272), .B2(\out_bs[6] [5]), 
      .ZN(n_8_0_5270));
   AOI21_X1 i_8_0_5488 (.A(n_8_0_5456), .B1(n_8_0_6590), .B2(n_8_0_402), 
      .ZN(n_8_0_5271));
   OAI21_X1 i_8_0_5489 (.A(n_8_0_6750), .B1(n_8_0_6755), .B2(n_8_0_402), 
      .ZN(n_8_0_5272));
   OAI21_X1 i_8_0_5490 (.A(n_8_0_6249), .B1(n_8_0_5274), .B2(n_8_0_24), .ZN(
      n_8_0_5273));
   NOR2_X1 i_8_0_5491 (.A1(n_8_0_6815), .A2(\out_bs[0] [6]), .ZN(n_8_0_5274));
   OAI211_X1 i_8_0_5492 (.A(n_8_0_7084), .B(n_8_0_6662), .C1(n_8_0_6811), 
      .C2(n_8_0_24), .ZN(n_8_0_5275));
   AOI211_X1 i_8_0_5493 (.A(n_8_0_5460), .B(n_8_0_5277), .C1(n_8_0_276), 
      .C2(n_8_0_6556), .ZN(n_8_0_5276));
   NOR2_X1 i_8_0_5494 (.A1(n_8_0_5278), .A2(\out_bs[4] [5]), .ZN(n_8_0_5277));
   OAI21_X1 i_8_0_5495 (.A(n_8_0_6632), .B1(n_8_0_6795), .B2(n_8_0_276), 
      .ZN(n_8_0_5278));
   NOR2_X1 i_8_0_5496 (.A1(n_8_0_5279), .A2(n_8_0_6853), .ZN(n_157));
   AOI211_X1 i_8_0_5497 (.A(n_8_0_5285), .B(n_8_0_5280), .C1(n_8_0_6233), 
      .C2(n_8_0_5286), .ZN(n_8_0_5279));
   OAI21_X1 i_8_0_5498 (.A(n_8_0_5281), .B1(n_8_0_5298), .B2(n_8_0_25), .ZN(
      n_8_0_5280));
   NOR4_X1 i_8_0_5499 (.A1(n_8_0_5303), .A2(n_8_0_5282), .A3(n_8_0_5288), 
      .A4(n_8_0_5283), .ZN(n_8_0_5281));
   OR3_X1 i_8_0_5500 (.A1(n_8_0_6248), .A2(n_8_0_5299), .A3(n_8_0_5293), 
      .ZN(n_8_0_5282));
   NAND3_X1 i_8_0_5501 (.A1(n_8_0_5295), .A2(n_8_0_5290), .A3(n_8_0_5284), 
      .ZN(n_8_0_5283));
   NAND2_X1 i_8_0_5502 (.A1(n_8_0_6343), .A2(n_8_0_6250), .ZN(n_8_0_5284));
   NOR2_X1 i_8_0_5503 (.A1(n_8_0_466), .A2(n_8_0_5287), .ZN(n_8_0_5285));
   NAND2_X1 i_8_0_5504 (.A1(n_8_0_466), .A2(n_8_0_5287), .ZN(n_8_0_5286));
   OAI21_X1 i_8_0_5505 (.A(n_8_0_5481), .B1(n_8_0_6363), .B2(n_8_0_6728), 
      .ZN(n_8_0_5287));
   AOI221_X1 i_8_0_5506 (.A(n_8_0_5428), .B1(n_8_0_5426), .B2(n_8_0_6333), 
      .C1(n_8_0_5289), .C2(n_8_0_151), .ZN(n_8_0_5288));
   OAI21_X1 i_8_0_5507 (.A(n_8_0_6607), .B1(n_8_0_6334), .B2(\out_bs[2] [5]), 
      .ZN(n_8_0_5289));
   OAI21_X1 i_8_0_5508 (.A(n_8_0_5291), .B1(n_8_0_5292), .B2(n_8_0_6340), 
      .ZN(n_8_0_5290));
   OAI21_X1 i_8_0_5509 (.A(n_8_0_6526), .B1(n_8_0_5395), .B2(n_8_0_88), .ZN(
      n_8_0_5291));
   OAI21_X1 i_8_0_5510 (.A(n_8_0_7071), .B1(n_8_0_88), .B2(n_8_0_6782), .ZN(
      n_8_0_5292));
   AOI221_X1 i_8_0_5511 (.A(n_8_0_5456), .B1(n_8_0_5452), .B2(n_8_0_6366), 
      .C1(n_8_0_5294), .C2(n_8_0_403), .ZN(n_8_0_5293));
   OAI21_X1 i_8_0_5512 (.A(n_8_0_6591), .B1(n_8_0_6367), .B2(\out_bs[6] [5]), 
      .ZN(n_8_0_5294));
   OAI211_X1 i_8_0_5513 (.A(n_8_0_5459), .B(n_8_0_5296), .C1(n_8_0_5458), 
      .C2(n_8_0_6349), .ZN(n_8_0_5295));
   OAI21_X1 i_8_0_5514 (.A(n_8_0_277), .B1(n_8_0_6556), .B2(n_8_0_5297), 
      .ZN(n_8_0_5296));
   NOR2_X1 i_8_0_5515 (.A1(\out_bs[4] [5]), .A2(n_8_0_6349), .ZN(n_8_0_5297));
   AOI21_X1 i_8_0_5516 (.A(n_8_0_6594), .B1(n_8_0_6438), .B2(n_8_0_6344), 
      .ZN(n_8_0_5298));
   AOI211_X1 i_8_0_5517 (.A(n_8_0_5302), .B(n_8_0_5300), .C1(n_8_0_340), 
      .C2(n_8_0_6513), .ZN(n_8_0_5299));
   NOR2_X1 i_8_0_5518 (.A1(n_8_0_5301), .A2(\out_bs[5] [5]), .ZN(n_8_0_5300));
   OAI21_X1 i_8_0_5519 (.A(n_8_0_6372), .B1(n_8_0_6824), .B2(n_8_0_340), 
      .ZN(n_8_0_5301));
   NOR2_X1 i_8_0_5520 (.A1(n_8_0_6827), .A2(\out_bs[5] [6]), .ZN(n_8_0_5302));
   OAI21_X1 i_8_0_5521 (.A(n_8_0_5304), .B1(n_8_0_6837), .B2(n_8_0_214), 
      .ZN(n_8_0_5303));
   OAI211_X1 i_8_0_5522 (.A(n_8_0_5305), .B(\out_bs[3] [6]), .C1(\out_bs[3] [5]), 
      .C2(n_8_0_6356), .ZN(n_8_0_5304));
   NAND2_X1 i_8_0_5523 (.A1(n_8_0_6844), .A2(n_8_0_214), .ZN(n_8_0_5305));
   AOI21_X1 i_8_0_5524 (.A(n_8_0_6853), .B1(n_8_0_5306), .B2(n_8_0_5328), 
      .ZN(n_158));
   NOR4_X1 i_8_0_5525 (.A1(n_8_0_5318), .A2(n_8_0_5307), .A3(n_8_0_5316), 
      .A4(n_8_0_5323), .ZN(n_8_0_5306));
   OAI211_X1 i_8_0_5526 (.A(n_8_0_5308), .B(n_8_0_5309), .C1(n_8_0_5317), 
      .C2(n_8_0_6812), .ZN(n_8_0_5307));
   NOR4_X1 i_8_0_5527 (.A1(n_8_0_5321), .A2(n_8_0_6248), .A3(n_8_0_5326), 
      .A4(n_8_0_5312), .ZN(n_8_0_5308));
   OAI21_X1 i_8_0_5528 (.A(n_8_0_5310), .B1(n_8_0_5311), .B2(n_8_0_6233), 
      .ZN(n_8_0_5309));
   OAI211_X1 i_8_0_5529 (.A(n_8_0_467), .B(n_8_0_6727), .C1(n_8_0_6543), 
      .C2(n_8_0_6405), .ZN(n_8_0_5310));
   AOI211_X1 i_8_0_5530 (.A(n_8_0_467), .B(n_8_0_5482), .C1(n_8_0_6405), 
      .C2(n_8_0_6727), .ZN(n_8_0_5311));
   INV_X1 i_8_0_5531 (.A(n_8_0_5313), .ZN(n_8_0_5312));
   AOI21_X1 i_8_0_5532 (.A(n_8_0_5314), .B1(n_8_0_6773), .B2(n_8_0_6957), 
      .ZN(n_8_0_5313));
   AOI21_X1 i_8_0_5533 (.A(n_8_0_5315), .B1(n_8_0_6772), .B2(n_8_0_152), 
      .ZN(n_8_0_5314));
   AOI21_X1 i_8_0_5534 (.A(n_8_0_6712), .B1(n_8_0_6398), .B2(\out_bs[2] [6]), 
      .ZN(n_8_0_5315));
   AOI21_X1 i_8_0_5535 (.A(n_8_0_26), .B1(n_8_0_6595), .B2(n_8_0_5317), .ZN(
      n_8_0_5316));
   NAND2_X1 i_8_0_5536 (.A1(n_8_0_6438), .A2(n_8_0_6420), .ZN(n_8_0_5317));
   AOI21_X1 i_8_0_5537 (.A(n_8_0_5319), .B1(n_8_0_5320), .B2(n_8_0_404), 
      .ZN(n_8_0_5318));
   OAI21_X1 i_8_0_5538 (.A(n_8_0_5455), .B1(n_8_0_5451), .B2(n_8_0_6385), 
      .ZN(n_8_0_5319));
   OAI21_X1 i_8_0_5539 (.A(n_8_0_6591), .B1(n_8_0_6385), .B2(\out_bs[6] [5]), 
      .ZN(n_8_0_5320));
   OAI221_X1 i_8_0_5540 (.A(n_8_0_6511), .B1(n_8_0_6408), .B2(n_8_0_5470), 
      .C1(n_8_0_5322), .C2(n_8_0_341), .ZN(n_8_0_5321));
   AOI21_X1 i_8_0_5541 (.A(n_8_0_6375), .B1(n_8_0_6409), .B2(n_8_0_6686), 
      .ZN(n_8_0_5322));
   OAI21_X1 i_8_0_5542 (.A(n_8_0_5324), .B1(n_8_0_6837), .B2(n_8_0_215), 
      .ZN(n_8_0_5323));
   OAI211_X1 i_8_0_5543 (.A(n_8_0_5325), .B(\out_bs[3] [6]), .C1(\out_bs[3] [5]), 
      .C2(n_8_0_6412), .ZN(n_8_0_5324));
   NAND2_X1 i_8_0_5544 (.A1(n_8_0_6844), .A2(n_8_0_215), .ZN(n_8_0_5325));
   OAI211_X1 i_8_0_5545 (.A(n_8_0_6525), .B(n_8_0_5327), .C1(n_8_0_6265), 
      .C2(n_8_0_89), .ZN(n_8_0_5326));
   OAI211_X1 i_8_0_5546 (.A(\out_bs[1] [6]), .B(n_8_0_6393), .C1(n_8_0_6783), 
      .C2(n_8_0_6976), .ZN(n_8_0_5327));
   OAI211_X1 i_8_0_5547 (.A(n_8_0_5459), .B(n_8_0_5329), .C1(n_8_0_5458), 
      .C2(n_8_0_6380), .ZN(n_8_0_5328));
   OAI21_X1 i_8_0_5548 (.A(n_8_0_278), .B1(n_8_0_6556), .B2(n_8_0_5330), 
      .ZN(n_8_0_5329));
   NOR2_X1 i_8_0_5549 (.A1(\out_bs[4] [5]), .A2(n_8_0_6380), .ZN(n_8_0_5330));
   NOR2_X1 i_8_0_5550 (.A1(n_8_0_5331), .A2(n_8_0_6853), .ZN(n_159));
   NOR3_X1 i_8_0_5551 (.A1(n_8_0_5353), .A2(n_8_0_5332), .A3(n_8_0_5351), 
      .ZN(n_8_0_5331));
   NAND3_X1 i_8_0_5552 (.A1(n_8_0_5333), .A2(n_8_0_5348), .A3(n_8_0_5345), 
      .ZN(n_8_0_5332));
   NOR4_X1 i_8_0_5553 (.A1(n_8_0_5339), .A2(n_8_0_5334), .A3(n_8_0_5338), 
      .A4(n_8_0_5341), .ZN(n_8_0_5333));
   OAI211_X1 i_8_0_5554 (.A(n_8_0_6247), .B(n_8_0_5335), .C1(n_8_0_27), .C2(
      n_8_0_6595), .ZN(n_8_0_5334));
   OAI211_X1 i_8_0_5555 (.A(n_8_0_5427), .B(n_8_0_5336), .C1(n_8_0_5425), 
      .C2(n_8_0_6451), .ZN(n_8_0_5335));
   OAI21_X1 i_8_0_5556 (.A(n_8_0_153), .B1(n_8_0_6606), .B2(n_8_0_5337), 
      .ZN(n_8_0_5336));
   NOR2_X1 i_8_0_5557 (.A1(\out_bs[2] [5]), .A2(n_8_0_6451), .ZN(n_8_0_5337));
   AOI211_X1 i_8_0_5558 (.A(n_8_0_6442), .B(n_8_0_6437), .C1(n_8_0_6812), 
      .C2(n_8_0_27), .ZN(n_8_0_5338));
   OAI211_X1 i_8_0_5559 (.A(n_8_0_6525), .B(n_8_0_5340), .C1(n_8_0_6265), 
      .C2(n_8_0_90), .ZN(n_8_0_5339));
   OAI211_X1 i_8_0_5560 (.A(\out_bs[1] [6]), .B(n_8_0_6446), .C1(n_8_0_6783), 
      .C2(n_8_0_6975), .ZN(n_8_0_5340));
   AOI21_X1 i_8_0_5561 (.A(n_8_0_5343), .B1(n_8_0_5342), .B2(n_8_0_6232), 
      .ZN(n_8_0_5341));
   OR2_X1 i_8_0_5562 (.A1(n_8_0_468), .A2(n_8_0_5344), .ZN(n_8_0_5342));
   AND2_X1 i_8_0_5563 (.A1(n_8_0_468), .A2(n_8_0_5344), .ZN(n_8_0_5343));
   OAI21_X1 i_8_0_5564 (.A(n_8_0_5481), .B1(n_8_0_6475), .B2(n_8_0_6728), 
      .ZN(n_8_0_5344));
   AOI21_X1 i_8_0_5565 (.A(n_8_0_5346), .B1(n_8_0_6838), .B2(n_8_0_6927), 
      .ZN(n_8_0_5345));
   AOI21_X1 i_8_0_5566 (.A(n_8_0_5347), .B1(n_8_0_6844), .B2(n_8_0_216), 
      .ZN(n_8_0_5346));
   AOI21_X1 i_8_0_5567 (.A(n_8_0_6659), .B1(n_8_0_6657), .B2(n_8_0_6427), 
      .ZN(n_8_0_5347));
   OAI21_X1 i_8_0_5568 (.A(n_8_0_5350), .B1(n_8_0_5349), .B2(\out_bs[4] [5]), 
      .ZN(n_8_0_5348));
   OAI21_X1 i_8_0_5569 (.A(n_8_0_6433), .B1(n_8_0_6795), .B2(n_8_0_279), 
      .ZN(n_8_0_5349));
   OAI21_X1 i_8_0_5570 (.A(n_8_0_6556), .B1(n_8_0_5460), .B2(n_8_0_279), 
      .ZN(n_8_0_5350));
   AOI221_X1 i_8_0_5571 (.A(n_8_0_5456), .B1(n_8_0_5452), .B2(n_8_0_6478), 
      .C1(n_8_0_5352), .C2(n_8_0_405), .ZN(n_8_0_5351));
   OAI21_X1 i_8_0_5572 (.A(n_8_0_6591), .B1(n_8_0_6479), .B2(\out_bs[6] [5]), 
      .ZN(n_8_0_5352));
   OAI211_X1 i_8_0_5573 (.A(n_8_0_6511), .B(n_8_0_5354), .C1(n_8_0_6376), 
      .C2(n_8_0_342), .ZN(n_8_0_5353));
   NAND3_X1 i_8_0_5574 (.A1(n_8_0_5355), .A2(n_8_0_6460), .A3(n_8_0_6686), 
      .ZN(n_8_0_5354));
   NAND2_X1 i_8_0_5575 (.A1(n_8_0_6619), .A2(n_8_0_342), .ZN(n_8_0_5355));
   AOI21_X1 i_8_0_5581 (.A(n_8_0_6248), .B1(n_8_0_6438), .B2(\out_bs[0] [2]), 
      .ZN(n_8_0_5360));
   OAI21_X1 i_8_0_5584 (.A(n_8_0_154), .B1(n_8_0_6606), .B2(n_8_0_5364), 
      .ZN(n_8_0_5363));
   NOR2_X1 i_8_0_5585 (.A1(\out_bs[2] [5]), .A2(n_8_0_6707), .ZN(n_8_0_5364));
   NAND4_X1 i_8_0_5587 (.A1(n_8_0_5367), .A2(n_8_0_6696), .A3(\out_bs[1] [2]), 
      .A4(\out_bs[1] [6]), .ZN(n_8_0_5366));
   NAND2_X1 i_8_0_5588 (.A1(n_8_0_6784), .A2(n_8_0_91), .ZN(n_8_0_5367));
   OAI21_X1 i_8_0_5589 (.A(n_8_0_5369), .B1(n_8_0_5370), .B2(\out_bs[6] [5]), 
      .ZN(n_8_0_5368));
   AOI21_X1 i_8_0_5590 (.A(n_8_0_5456), .B1(n_8_0_6590), .B2(n_8_0_406), 
      .ZN(n_8_0_5369));
   OAI21_X1 i_8_0_5591 (.A(n_8_0_6748), .B1(n_8_0_6755), .B2(n_8_0_406), 
      .ZN(n_8_0_5370));
   OAI21_X1 i_8_0_5593 (.A(n_8_0_5459), .B1(n_8_0_5458), .B2(n_8_0_6631), 
      .ZN(n_8_0_5372));
   OAI21_X1 i_8_0_5594 (.A(n_8_0_6557), .B1(n_8_0_6631), .B2(\out_bs[4] [5]), 
      .ZN(n_8_0_5373));
   OAI211_X1 i_8_0_5596 (.A(n_8_0_5376), .B(\out_bs[3] [6]), .C1(\out_bs[3] [5]), 
      .C2(n_8_0_5468), .ZN(n_8_0_5375));
   NAND2_X1 i_8_0_5597 (.A1(n_8_0_6844), .A2(n_8_0_217), .ZN(n_8_0_5376));
   NAND3_X1 i_8_0_5599 (.A1(n_8_0_5379), .A2(n_8_0_6679), .A3(n_8_0_6686), 
      .ZN(n_8_0_5378));
   NAND2_X1 i_8_0_5600 (.A1(n_8_0_6824), .A2(n_8_0_343), .ZN(n_8_0_5379));
   NOR3_X1 i_8_0_5604 (.A1(n_8_0_6248), .A2(n_8_0_5387), .A3(n_8_0_5383), 
      .ZN(n_8_0_5382));
   INV_X1 i_8_0_5605 (.A(n_8_0_5384), .ZN(n_8_0_5383));
   OAI211_X1 i_8_0_5606 (.A(n_8_0_5455), .B(n_8_0_5385), .C1(n_8_0_5451), 
      .C2(n_8_0_6549), .ZN(n_8_0_5384));
   OAI21_X1 i_8_0_5607 (.A(n_8_0_407), .B1(n_8_0_6590), .B2(n_8_0_5386), 
      .ZN(n_8_0_5385));
   NOR2_X1 i_8_0_5608 (.A1(\out_bs[6] [5]), .A2(n_8_0_6549), .ZN(n_8_0_5386));
   AOI211_X1 i_8_0_5609 (.A(n_8_0_6523), .B(n_8_0_6437), .C1(n_8_0_6812), 
      .C2(n_8_0_29), .ZN(n_8_0_5387));
   NAND3_X1 i_8_0_5611 (.A1(\out_bs[3] [6]), .A2(n_8_0_6648), .A3(n_8_0_5390), 
      .ZN(n_8_0_5389));
   AOI21_X1 i_8_0_5612 (.A(n_8_0_6566), .B1(n_8_0_6844), .B2(n_8_0_218), 
      .ZN(n_8_0_5390));
   AOI21_X1 i_8_0_5615 (.A(\out_bs[1] [5]), .B1(n_8_0_6974), .B2(n_8_0_6781), 
      .ZN(n_8_0_5393));
   NAND2_X1 i_8_0_5616 (.A1(n_8_0_5397), .A2(n_8_0_7072), .ZN(n_8_0_5394));
   NOR2_X1 i_8_0_5617 (.A1(n_8_0_5396), .A2(\out_bs[1] [6]), .ZN(n_8_0_5395));
   NAND2_X1 i_8_0_5618 (.A1(n_8_0_6786), .A2(n_8_0_7078), .ZN(n_8_0_5396));
   NOR2_X1 i_8_0_5619 (.A1(n_8_0_6785), .A2(\out_as[1] [6]), .ZN(n_8_0_5397));
   AOI22_X1 i_8_0_5621 (.A1(n_8_0_6956), .A2(n_8_0_6773), .B1(n_8_0_5400), 
      .B2(\out_bs[2] [6]), .ZN(n_8_0_5399));
   OAI21_X1 i_8_0_5622 (.A(n_8_0_7059), .B1(n_8_0_6537), .B2(n_8_0_6708), 
      .ZN(n_8_0_5400));
   AOI21_X1 i_8_0_5628 (.A(n_8_0_6375), .B1(n_8_0_6516), .B2(n_8_0_6686), 
      .ZN(n_8_0_5406));
   OAI21_X1 i_8_0_5630 (.A(n_8_0_6557), .B1(n_8_0_6558), .B2(\out_bs[4] [5]), 
      .ZN(n_8_0_5408));
   NOR2_X1 i_8_0_5631 (.A1(\out_bs[4] [5]), .A2(n_8_0_6558), .ZN(n_8_0_5409));
   AOI221_X1 i_8_0_5638 (.A(n_8_0_7047), .B1(n_8_0_7046), .B2(n_8_0_6579), 
      .C1(n_8_0_6844), .C2(n_8_0_219), .ZN(n_8_0_5415));
   OAI21_X1 i_8_0_5640 (.A(n_8_0_5418), .B1(n_8_0_5472), .B2(n_8_0_6375), 
      .ZN(n_8_0_5417));
   OAI21_X1 i_8_0_5641 (.A(n_8_0_345), .B1(n_8_0_6675), .B2(n_8_0_5470), 
      .ZN(n_8_0_5418));
   INV_X1 i_8_0_5642 (.A(n_8_0_5420), .ZN(n_8_0_5419));
   AOI21_X1 i_8_0_5644 (.A(n_8_0_408), .B1(n_8_0_5452), .B2(n_8_0_6741), 
      .ZN(n_8_0_5421));
   AOI21_X1 i_8_0_5645 (.A(n_8_0_6590), .B1(n_8_0_6741), .B2(n_8_0_7011), 
      .ZN(n_8_0_5422));
   OAI21_X1 i_8_0_5647 (.A(n_8_0_6607), .B1(n_8_0_6611), .B2(\out_bs[2] [5]), 
      .ZN(n_8_0_5424));
   NAND2_X1 i_8_0_5648 (.A1(n_8_0_7059), .A2(n_8_0_6772), .ZN(n_8_0_5425));
   NOR2_X1 i_8_0_5649 (.A1(\out_bs[2] [5]), .A2(n_8_0_6773), .ZN(n_8_0_5426));
   NAND2_X1 i_8_0_5650 (.A1(n_8_0_6774), .A2(n_8_0_7060), .ZN(n_8_0_5427));
   NOR2_X1 i_8_0_5651 (.A1(n_8_0_6775), .A2(\out_bs[2] [6]), .ZN(n_8_0_5428));
   INV_X1 i_8_0_5652 (.A(n_8_0_5430), .ZN(n_8_0_5429));
   NAND3_X1 i_8_0_5654 (.A1(\out_bs[1] [6]), .A2(n_8_0_6700), .A3(n_8_0_5432), 
      .ZN(n_8_0_5431));
   AOI21_X1 i_8_0_5655 (.A(n_8_0_6695), .B1(n_8_0_6784), .B2(n_8_0_93), .ZN(
      n_8_0_5432));
   INV_X1 i_8_0_5656 (.A(n_8_0_5434), .ZN(n_8_0_5433));
   AOI211_X1 i_8_0_5657 (.A(n_8_0_471), .B(n_8_0_5482), .C1(n_8_0_6724), 
      .C2(n_8_0_6727), .ZN(n_8_0_5434));
   INV_X1 i_8_0_5658 (.A(n_8_0_5436), .ZN(n_8_0_5435));
   NAND2_X1 i_8_0_5662 (.A1(n_8_0_6557), .A2(n_8_0_5441), .ZN(n_8_0_5439));
   AOI21_X1 i_8_0_5663 (.A(n_8_0_6794), .B1(n_8_0_5441), .B2(\out_bs[4] [6]), 
      .ZN(n_8_0_5440));
   OAI21_X1 i_8_0_5664 (.A(n_8_0_7034), .B1(n_8_0_6642), .B2(n_8_0_6632), 
      .ZN(n_8_0_5441));
   AOI21_X1 i_8_0_5665 (.A(\out_bs[4] [5]), .B1(n_8_0_6643), .B2(n_8_0_6633), 
      .ZN(n_8_0_5442));
   NOR2_X1 i_8_0_5666 (.A1(n_8_0_5443), .A2(n_8_0_6853), .ZN(n_160));
   NOR4_X1 i_8_0_5667 (.A1(n_8_0_5473), .A2(n_8_0_5469), .A3(n_8_0_5463), 
      .A4(n_8_0_5444), .ZN(n_8_0_5443));
   NAND4_X1 i_8_0_5668 (.A1(n_8_0_5457), .A2(n_8_0_5449), .A3(n_8_0_5446), 
      .A4(n_8_0_5445), .ZN(n_8_0_5444));
   AOI21_X1 i_8_0_5669 (.A(n_8_0_5479), .B1(n_8_0_6233), .B2(n_8_0_5478), 
      .ZN(n_8_0_5445));
   NOR3_X1 i_8_0_5670 (.A1(n_8_0_5476), .A2(n_8_0_5447), .A3(n_8_0_5483), 
      .ZN(n_8_0_5446));
   OAI21_X1 i_8_0_5671 (.A(n_8_0_6247), .B1(n_8_0_5484), .B2(n_8_0_6812), 
      .ZN(n_8_0_5447));
   INV_X1 i_8_0_5672 (.A(n_8_0_5449), .ZN(n_8_0_5448));
   OAI21_X1 i_8_0_5673 (.A(n_8_0_5450), .B1(n_8_0_5451), .B2(n_8_0_5454), 
      .ZN(n_8_0_5449));
   AOI21_X1 i_8_0_5674 (.A(n_8_0_5456), .B1(n_8_0_5453), .B2(n_8_0_409), 
      .ZN(n_8_0_5450));
   NAND2_X1 i_8_0_5675 (.A1(n_8_0_6755), .A2(n_8_0_7011), .ZN(n_8_0_5451));
   NOR2_X1 i_8_0_5676 (.A1(n_8_0_6754), .A2(\out_bs[6] [5]), .ZN(n_8_0_5452));
   OAI21_X1 i_8_0_5677 (.A(n_8_0_6591), .B1(n_8_0_5454), .B2(\out_bs[6] [5]), 
      .ZN(n_8_0_5453));
   NOR2_X1 i_8_0_5678 (.A1(n_8_0_6748), .A2(n_8_0_6745), .ZN(n_8_0_5454));
   NAND2_X1 i_8_0_5679 (.A1(n_8_0_6761), .A2(n_8_0_7012), .ZN(n_8_0_5455));
   NOR2_X1 i_8_0_5680 (.A1(n_8_0_6760), .A2(\out_bs[6] [6]), .ZN(n_8_0_5456));
   OAI211_X1 i_8_0_5681 (.A(n_8_0_5461), .B(n_8_0_5459), .C1(n_8_0_5458), 
      .C2(n_8_0_6628), .ZN(n_8_0_5457));
   NAND2_X1 i_8_0_5682 (.A1(n_8_0_6795), .A2(n_8_0_7034), .ZN(n_8_0_5458));
   NAND2_X1 i_8_0_5683 (.A1(n_8_0_6801), .A2(n_8_0_7035), .ZN(n_8_0_5459));
   NOR2_X1 i_8_0_5684 (.A1(n_8_0_6800), .A2(\out_bs[4] [6]), .ZN(n_8_0_5460));
   OAI21_X1 i_8_0_5685 (.A(n_8_0_283), .B1(n_8_0_6556), .B2(n_8_0_5462), 
      .ZN(n_8_0_5461));
   NOR2_X1 i_8_0_5686 (.A1(\out_bs[4] [5]), .A2(n_8_0_6628), .ZN(n_8_0_5462));
   OAI21_X1 i_8_0_5687 (.A(n_8_0_5464), .B1(n_8_0_6837), .B2(n_8_0_220), 
      .ZN(n_8_0_5463));
   OAI21_X1 i_8_0_5688 (.A(n_8_0_5465), .B1(n_8_0_6843), .B2(n_8_0_6925), 
      .ZN(n_8_0_5464));
   OAI21_X1 i_8_0_5689 (.A(n_8_0_6658), .B1(n_8_0_5466), .B2(n_8_0_7047), 
      .ZN(n_8_0_5465));
   NAND2_X1 i_8_0_5690 (.A1(n_8_0_6650), .A2(n_8_0_6648), .ZN(n_8_0_5466));
   NAND2_X1 i_8_0_5691 (.A1(\out_bs[3] [2]), .A2(n_8_0_6648), .ZN(n_8_0_5467));
   NOR2_X1 i_8_0_5692 (.A1(n_8_0_7043), .A2(n_8_0_6647), .ZN(n_8_0_5468));
   OAI221_X1 i_8_0_5693 (.A(n_8_0_6511), .B1(n_8_0_5470), .B2(n_8_0_6673), 
      .C1(n_8_0_5471), .C2(n_8_0_346), .ZN(n_8_0_5469));
   NAND2_X1 i_8_0_5694 (.A1(\out_bs[5] [4]), .A2(n_8_0_6514), .ZN(n_8_0_5470));
   AOI21_X1 i_8_0_5695 (.A(n_8_0_6375), .B1(n_8_0_6674), .B2(n_8_0_6686), 
      .ZN(n_8_0_5471));
   AND2_X1 i_8_0_5696 (.A1(n_8_0_6686), .A2(n_8_0_6676), .ZN(n_8_0_5472));
   OAI21_X1 i_8_0_5697 (.A(n_8_0_5474), .B1(n_8_0_6772), .B2(n_8_0_157), 
      .ZN(n_8_0_5473));
   OAI211_X1 i_8_0_5698 (.A(n_8_0_5475), .B(\out_bs[2] [6]), .C1(\out_bs[2] [5]), 
      .C2(n_8_0_6704), .ZN(n_8_0_5474));
   NAND2_X1 i_8_0_5699 (.A1(n_8_0_6772), .A2(n_8_0_157), .ZN(n_8_0_5475));
   OAI211_X1 i_8_0_5700 (.A(n_8_0_6525), .B(n_8_0_5477), .C1(n_8_0_6265), 
      .C2(n_8_0_94), .ZN(n_8_0_5476));
   OAI211_X1 i_8_0_5701 (.A(\out_bs[1] [6]), .B(n_8_0_6688), .C1(n_8_0_6783), 
      .C2(n_8_0_6973), .ZN(n_8_0_5477));
   OAI211_X1 i_8_0_5702 (.A(n_8_0_472), .B(n_8_0_6727), .C1(n_8_0_6722), 
      .C2(n_8_0_6543), .ZN(n_8_0_5478));
   AOI211_X1 i_8_0_5703 (.A(n_8_0_472), .B(n_8_0_5482), .C1(n_8_0_6722), 
      .C2(n_8_0_6727), .ZN(n_8_0_5479));
   NAND2_X1 i_8_0_5705 (.A1(n_8_0_6727), .A2(n_8_0_6543), .ZN(n_8_0_5481));
   AOI21_X1 i_8_0_5706 (.A(n_8_0_6728), .B1(n_8_0_6717), .B2(\out_bs[7] [3]), 
      .ZN(n_8_0_5482));
   AOI21_X1 i_8_0_5707 (.A(n_8_0_31), .B1(n_8_0_6595), .B2(n_8_0_5484), .ZN(
      n_8_0_5483));
   NAND2_X1 i_8_0_5708 (.A1(n_8_0_6666), .A2(n_8_0_6438), .ZN(n_8_0_5484));
   AOI21_X1 i_8_0_5709 (.A(n_8_0_6853), .B1(n_8_0_5487), .B2(n_8_0_5485), 
      .ZN(n_161));
   NOR4_X1 i_8_0_5710 (.A1(n_8_0_5486), .A2(n_8_0_5490), .A3(n_8_0_5492), 
      .A4(n_8_0_5494), .ZN(n_8_0_5485));
   OR2_X1 i_8_0_5711 (.A1(n_8_0_5489), .A2(n_8_0_5496), .ZN(n_8_0_5486));
   NOR4_X1 i_8_0_5712 (.A1(n_8_0_6248), .A2(n_8_0_5491), .A3(n_8_0_5488), 
      .A4(n_8_0_5495), .ZN(n_8_0_5487));
   OAI22_X1 i_8_0_5713 (.A1(n_8_0_6727), .A2(n_8_0_6232), .B1(n_8_0_6595), 
      .B2(n_8_0_32), .ZN(n_8_0_5488));
   OAI21_X1 i_8_0_5714 (.A(n_8_0_6554), .B1(n_8_0_5929), .B2(n_8_0_284), 
      .ZN(n_8_0_5489));
   AOI22_X1 i_8_0_5715 (.A1(n_8_0_6755), .A2(n_8_0_6752), .B1(n_8_0_6588), 
      .B2(n_8_0_410), .ZN(n_8_0_5490));
   OAI21_X1 i_8_0_5716 (.A(n_8_0_6511), .B1(n_8_0_6376), .B2(n_8_0_347), 
      .ZN(n_8_0_5491));
   OAI21_X1 i_8_0_5717 (.A(n_8_0_6604), .B1(n_8_0_5493), .B2(n_8_0_158), 
      .ZN(n_8_0_5492));
   NOR2_X1 i_8_0_5718 (.A1(n_8_0_6773), .A2(n_8_0_6712), .ZN(n_8_0_5493));
   AOI21_X1 i_8_0_5719 (.A(n_8_0_473), .B1(n_8_0_6727), .B2(n_8_0_6232), 
      .ZN(n_8_0_5494));
   AOI21_X1 i_8_0_5720 (.A(n_8_0_6265), .B1(n_8_0_6525), .B2(n_8_0_95), .ZN(
      n_8_0_5495));
   AOI21_X1 i_8_0_5721 (.A(n_8_0_6572), .B1(n_8_0_6575), .B2(n_8_0_221), 
      .ZN(n_8_0_5496));
   NOR2_X1 i_8_0_5722 (.A1(n_8_0_5497), .A2(n_8_0_6853), .ZN(n_162));
   NOR4_X1 i_8_0_5723 (.A1(n_8_0_5507), .A2(n_8_0_5503), .A3(n_8_0_5498), 
      .A4(n_8_0_5527), .ZN(n_8_0_5497));
   OAI21_X1 i_8_0_5724 (.A(n_8_0_5499), .B1(n_8_0_6837), .B2(n_8_0_222), 
      .ZN(n_8_0_5498));
   NAND3_X1 i_8_0_5725 (.A1(n_8_0_5502), .A2(n_8_0_5500), .A3(n_8_0_6659), 
      .ZN(n_8_0_5499));
   NAND2_X1 i_8_0_5726 (.A1(n_8_0_5564), .A2(n_8_0_7041), .ZN(n_8_0_5500));
   NOR2_X1 i_8_0_5727 (.A1(n_8_0_6357), .A2(n_8_0_6007), .ZN(n_8_0_5501));
   NAND2_X1 i_8_0_5728 (.A1(n_8_0_222), .A2(n_8_0_6842), .ZN(n_8_0_5502));
   AOI221_X1 i_8_0_5729 (.A(n_8_0_6595), .B1(n_8_0_5506), .B2(n_8_0_6811), 
      .C1(n_8_0_5504), .C2(n_8_0_33), .ZN(n_8_0_5503));
   NAND2_X1 i_8_0_5730 (.A1(n_8_0_6248), .A2(n_8_0_5505), .ZN(n_8_0_5504));
   NAND2_X1 i_8_0_5731 (.A1(n_8_0_6345), .A2(n_8_0_5944), .ZN(n_8_0_5505));
   NOR2_X1 i_8_0_5732 (.A1(n_8_0_5554), .A2(\out_bs[0] [0]), .ZN(n_8_0_5506));
   NAND4_X1 i_8_0_5733 (.A1(n_8_0_5516), .A2(n_8_0_5508), .A3(n_8_0_5523), 
      .A4(n_8_0_5520), .ZN(n_8_0_5507));
   AOI211_X1 i_8_0_5734 (.A(n_8_0_5512), .B(n_8_0_5509), .C1(n_8_0_5510), 
      .C2(n_8_0_6233), .ZN(n_8_0_5508));
   NOR2_X1 i_8_0_5735 (.A1(n_8_0_5511), .A2(n_8_0_474), .ZN(n_8_0_5509));
   NAND2_X1 i_8_0_5736 (.A1(n_8_0_5511), .A2(n_8_0_474), .ZN(n_8_0_5510));
   OAI21_X1 i_8_0_5737 (.A(n_8_0_6728), .B1(n_8_0_6363), .B2(n_8_0_5975), 
      .ZN(n_8_0_5511));
   INV_X1 i_8_0_5738 (.A(n_8_0_5513), .ZN(n_8_0_5512));
   OAI21_X1 i_8_0_5739 (.A(n_8_0_5514), .B1(n_8_0_6773), .B2(n_8_0_6955), 
      .ZN(n_8_0_5513));
   OAI22_X1 i_8_0_5740 (.A1(n_8_0_159), .A2(n_8_0_6772), .B1(n_8_0_6711), 
      .B2(n_8_0_5515), .ZN(n_8_0_5514));
   NOR2_X1 i_8_0_5741 (.A1(n_8_0_6335), .A2(n_8_0_5814), .ZN(n_8_0_5515));
   AOI21_X1 i_8_0_5742 (.A(n_8_0_5517), .B1(n_8_0_6825), .B2(n_8_0_6902), 
      .ZN(n_8_0_5516));
   AOI211_X1 i_8_0_5743 (.A(n_8_0_6685), .B(n_8_0_5518), .C1(n_8_0_6824), 
      .C2(n_8_0_348), .ZN(n_8_0_5517));
   INV_X1 i_8_0_5744 (.A(n_8_0_5519), .ZN(n_8_0_5518));
   NAND3_X1 i_8_0_5745 (.A1(n_8_0_6518), .A2(n_8_0_6166), .A3(n_8_0_7022), 
      .ZN(n_8_0_5519));
   AOI22_X1 i_8_0_5746 (.A1(n_8_0_5521), .A2(n_8_0_5522), .B1(n_8_0_6754), 
      .B2(n_8_0_6890), .ZN(n_8_0_5520));
   AOI21_X1 i_8_0_5747 (.A(n_8_0_6752), .B1(n_8_0_6758), .B2(n_8_0_411), 
      .ZN(n_8_0_5521));
   NAND2_X1 i_8_0_5748 (.A1(n_8_0_5543), .A2(n_8_0_7006), .ZN(n_8_0_5522));
   OAI211_X1 i_8_0_5749 (.A(n_8_0_6264), .B(n_8_0_5524), .C1(n_8_0_5525), 
      .C2(n_8_0_6781), .ZN(n_8_0_5523));
   OAI21_X1 i_8_0_5750 (.A(n_8_0_96), .B1(n_8_0_6525), .B2(n_8_0_5526), .ZN(
      n_8_0_5524));
   NAND2_X1 i_8_0_5751 (.A1(n_8_0_6342), .A2(n_8_0_5984), .ZN(n_8_0_5525));
   NOR2_X1 i_8_0_5752 (.A1(n_8_0_5547), .A2(\out_bs[1] [0]), .ZN(n_8_0_5526));
   AOI22_X1 i_8_0_5753 (.A1(n_8_0_285), .A2(n_8_0_5529), .B1(n_8_0_6795), 
      .B2(n_8_0_5528), .ZN(n_8_0_5527));
   OAI21_X1 i_8_0_5754 (.A(n_8_0_6636), .B1(n_8_0_6352), .B2(n_8_0_5744), 
      .ZN(n_8_0_5528));
   OAI21_X1 i_8_0_5755 (.A(n_8_0_6555), .B1(n_8_0_6031), .B2(\out_bs[4] [4]), 
      .ZN(n_8_0_5529));
   AOI21_X1 i_8_0_5756 (.A(n_8_0_6853), .B1(n_8_0_5533), .B2(n_8_0_5530), 
      .ZN(n_163));
   NOR4_X1 i_8_0_5757 (.A1(n_8_0_5538), .A2(n_8_0_5534), .A3(n_8_0_5532), 
      .A4(n_8_0_5531), .ZN(n_8_0_5530));
   OAI211_X1 i_8_0_5758 (.A(n_8_0_5561), .B(n_8_0_5545), .C1(n_8_0_34), .C2(
      n_8_0_6811), .ZN(n_8_0_5531));
   AOI211_X1 i_8_0_5759 (.A(n_8_0_6670), .B(n_8_0_5553), .C1(n_8_0_6812), 
      .C2(n_8_0_34), .ZN(n_8_0_5532));
   NOR4_X1 i_8_0_5760 (.A1(n_8_0_5556), .A2(n_8_0_5555), .A3(n_8_0_5549), 
      .A4(n_8_0_5541), .ZN(n_8_0_5533));
   AOI221_X1 i_8_0_5761 (.A(n_8_0_5929), .B1(n_8_0_5535), .B2(n_8_0_5536), 
      .C1(n_8_0_286), .C2(n_8_0_6554), .ZN(n_8_0_5534));
   OR2_X1 i_8_0_5762 (.A1(n_8_0_286), .A2(n_8_0_6795), .ZN(n_8_0_5535));
   NOR2_X1 i_8_0_5763 (.A1(n_8_0_6382), .A2(n_8_0_5744), .ZN(n_8_0_5536));
   INV_X1 i_8_0_5764 (.A(n_8_0_5538), .ZN(n_8_0_5537));
   AOI211_X1 i_8_0_5765 (.A(n_8_0_6376), .B(n_8_0_5539), .C1(n_8_0_5540), 
      .C2(n_8_0_349), .ZN(n_8_0_5538));
   NOR3_X1 i_8_0_5766 (.A1(\out_bs[5] [4]), .A2(n_8_0_6825), .A3(n_8_0_6097), 
      .ZN(n_8_0_5539));
   OAI21_X1 i_8_0_5767 (.A(n_8_0_6512), .B1(n_8_0_6097), .B2(\out_bs[5] [4]), 
      .ZN(n_8_0_5540));
   OAI21_X1 i_8_0_5768 (.A(n_8_0_5542), .B1(n_8_0_6755), .B2(n_8_0_412), 
      .ZN(n_8_0_5541));
   OAI211_X1 i_8_0_5769 (.A(n_8_0_6753), .B(n_8_0_5544), .C1(n_8_0_6759), 
      .C2(n_8_0_6889), .ZN(n_8_0_5542));
   INV_X1 i_8_0_5770 (.A(n_8_0_5544), .ZN(n_8_0_5543));
   NAND2_X1 i_8_0_5771 (.A1(n_8_0_6387), .A2(n_8_0_5894), .ZN(n_8_0_5544));
   OAI211_X1 i_8_0_5772 (.A(n_8_0_6264), .B(n_8_0_5546), .C1(n_8_0_5547), 
      .C2(n_8_0_6781), .ZN(n_8_0_5545));
   OAI21_X1 i_8_0_5773 (.A(n_8_0_97), .B1(n_8_0_6525), .B2(n_8_0_5548), .ZN(
      n_8_0_5546));
   NAND2_X1 i_8_0_5774 (.A1(n_8_0_6395), .A2(n_8_0_5984), .ZN(n_8_0_5547));
   NOR2_X1 i_8_0_5775 (.A1(n_8_0_6394), .A2(n_8_0_5983), .ZN(n_8_0_5548));
   AOI21_X1 i_8_0_5776 (.A(n_8_0_5550), .B1(n_8_0_6772), .B2(n_8_0_160), 
      .ZN(n_8_0_5549));
   INV_X1 i_8_0_5777 (.A(n_8_0_5551), .ZN(n_8_0_5550));
   OAI22_X1 i_8_0_5778 (.A1(n_8_0_160), .A2(n_8_0_6772), .B1(n_8_0_6711), 
      .B2(n_8_0_5552), .ZN(n_8_0_5551));
   NOR2_X1 i_8_0_5779 (.A1(n_8_0_6399), .A2(n_8_0_5814), .ZN(n_8_0_5552));
   INV_X1 i_8_0_5780 (.A(n_8_0_5554), .ZN(n_8_0_5553));
   NAND2_X1 i_8_0_5781 (.A1(n_8_0_6421), .A2(n_8_0_5944), .ZN(n_8_0_5554));
   NOR2_X1 i_8_0_5782 (.A1(n_8_0_5559), .A2(n_8_0_475), .ZN(n_8_0_5555));
   INV_X1 i_8_0_5783 (.A(n_8_0_5557), .ZN(n_8_0_5556));
   NAND2_X1 i_8_0_5784 (.A1(n_8_0_6233), .A2(n_8_0_5558), .ZN(n_8_0_5557));
   NAND2_X1 i_8_0_5785 (.A1(n_8_0_5559), .A2(n_8_0_475), .ZN(n_8_0_5558));
   NAND2_X1 i_8_0_5786 (.A1(n_8_0_5560), .A2(n_8_0_6728), .ZN(n_8_0_5559));
   NAND2_X1 i_8_0_5787 (.A1(n_8_0_6405), .A2(n_8_0_5976), .ZN(n_8_0_5560));
   OAI21_X1 i_8_0_5788 (.A(n_8_0_5563), .B1(n_8_0_5562), .B2(n_8_0_6838), 
      .ZN(n_8_0_5561));
   NOR2_X1 i_8_0_5789 (.A1(n_8_0_5564), .A2(n_8_0_6658), .ZN(n_8_0_5562));
   OAI21_X1 i_8_0_5790 (.A(n_8_0_223), .B1(n_8_0_6575), .B2(n_8_0_5564), 
      .ZN(n_8_0_5563));
   NOR2_X1 i_8_0_5791 (.A1(n_8_0_6413), .A2(n_8_0_6007), .ZN(n_8_0_5564));
   AOI21_X1 i_8_0_5792 (.A(n_8_0_6853), .B1(n_8_0_5567), .B2(n_8_0_5565), 
      .ZN(n_164));
   NOR3_X1 i_8_0_5793 (.A1(n_8_0_5566), .A2(n_8_0_5582), .A3(n_8_0_5584), 
      .ZN(n_8_0_5565));
   NAND3_X1 i_8_0_5794 (.A1(n_8_0_5578), .A2(n_8_0_5575), .A3(n_8_0_5570), 
      .ZN(n_8_0_5566));
   AOI211_X1 i_8_0_5795 (.A(n_8_0_5591), .B(n_8_0_5568), .C1(n_8_0_6233), 
      .C2(n_8_0_5592), .ZN(n_8_0_5567));
   OAI211_X1 i_8_0_5796 (.A(n_8_0_5587), .B(n_8_0_5569), .C1(n_8_0_35), .C2(
      n_8_0_6811), .ZN(n_8_0_5568));
   OAI211_X1 i_8_0_5797 (.A(n_8_0_6671), .B(n_8_0_5595), .C1(n_8_0_6813), 
      .C2(n_8_0_6985), .ZN(n_8_0_5569));
   NAND2_X1 i_8_0_5798 (.A1(n_8_0_5571), .A2(n_8_0_5572), .ZN(n_8_0_5570));
   OAI21_X1 i_8_0_5799 (.A(n_8_0_6795), .B1(n_8_0_6635), .B2(n_8_0_5573), 
      .ZN(n_8_0_5571));
   OAI21_X1 i_8_0_5800 (.A(n_8_0_287), .B1(n_8_0_6554), .B2(n_8_0_5573), 
      .ZN(n_8_0_5572));
   NOR2_X1 i_8_0_5801 (.A1(n_8_0_6435), .A2(n_8_0_5744), .ZN(n_8_0_5573));
   INV_X1 i_8_0_5802 (.A(n_8_0_5575), .ZN(n_8_0_5574));
   OAI21_X1 i_8_0_5803 (.A(n_8_0_5576), .B1(n_8_0_5577), .B2(n_8_0_6461), 
      .ZN(n_8_0_5575));
   OAI21_X1 i_8_0_5804 (.A(n_8_0_6511), .B1(n_8_0_6376), .B2(n_8_0_350), 
      .ZN(n_8_0_5576));
   OAI21_X1 i_8_0_5805 (.A(n_8_0_5748), .B1(n_8_0_6824), .B2(n_8_0_350), 
      .ZN(n_8_0_5577));
   OAI21_X1 i_8_0_5806 (.A(n_8_0_5580), .B1(n_8_0_5579), .B2(n_8_0_6838), 
      .ZN(n_8_0_5578));
   NOR2_X1 i_8_0_5807 (.A1(n_8_0_5581), .A2(n_8_0_6658), .ZN(n_8_0_5579));
   OAI21_X1 i_8_0_5808 (.A(n_8_0_224), .B1(n_8_0_6575), .B2(n_8_0_5581), 
      .ZN(n_8_0_5580));
   NOR2_X1 i_8_0_5809 (.A1(n_8_0_6428), .A2(n_8_0_6007), .ZN(n_8_0_5581));
   OAI22_X1 i_8_0_5810 (.A1(n_8_0_6752), .A2(n_8_0_5583), .B1(n_8_0_413), 
      .B2(n_8_0_6755), .ZN(n_8_0_5582));
   OAI22_X1 i_8_0_5811 (.A1(n_8_0_6759), .A2(n_8_0_6888), .B1(n_8_0_5893), 
      .B2(n_8_0_6480), .ZN(n_8_0_5583));
   OAI21_X1 i_8_0_5812 (.A(n_8_0_5585), .B1(n_8_0_6782), .B2(n_8_0_98), .ZN(
      n_8_0_5584));
   OAI211_X1 i_8_0_5813 (.A(n_8_0_6694), .B(n_8_0_5586), .C1(n_8_0_6783), 
      .C2(n_8_0_6972), .ZN(n_8_0_5585));
   NAND2_X1 i_8_0_5814 (.A1(n_8_0_6448), .A2(n_8_0_5984), .ZN(n_8_0_5586));
   AOI21_X1 i_8_0_5815 (.A(n_8_0_5590), .B1(n_8_0_5588), .B2(n_8_0_5589), 
      .ZN(n_8_0_5587));
   AOI21_X1 i_8_0_5816 (.A(n_8_0_6711), .B1(n_8_0_6772), .B2(n_8_0_161), 
      .ZN(n_8_0_5588));
   NAND2_X1 i_8_0_5817 (.A1(n_8_0_6453), .A2(n_8_0_5815), .ZN(n_8_0_5589));
   NOR2_X1 i_8_0_5818 (.A1(n_8_0_6772), .A2(n_8_0_161), .ZN(n_8_0_5590));
   NOR2_X1 i_8_0_5819 (.A1(n_8_0_5593), .A2(n_8_0_476), .ZN(n_8_0_5591));
   NAND2_X1 i_8_0_5820 (.A1(n_8_0_5593), .A2(n_8_0_476), .ZN(n_8_0_5592));
   NAND2_X1 i_8_0_5821 (.A1(n_8_0_5594), .A2(n_8_0_6728), .ZN(n_8_0_5593));
   NAND2_X1 i_8_0_5823 (.A1(n_8_0_6442), .A2(n_8_0_5944), .ZN(n_8_0_5595));
   NOR2_X1 i_8_0_5824 (.A1(n_8_0_5596), .A2(n_8_0_6853), .ZN(n_165));
   NOR4_X1 i_8_0_5825 (.A1(n_8_0_5603), .A2(n_8_0_5600), .A3(n_8_0_5597), 
      .A4(n_8_0_5608), .ZN(n_8_0_5596));
   OAI21_X1 i_8_0_5826 (.A(n_8_0_5598), .B1(n_8_0_6837), .B2(n_8_0_225), 
      .ZN(n_8_0_5597));
   OAI211_X1 i_8_0_5827 (.A(n_8_0_5599), .B(n_8_0_6659), .C1(\out_bs[3] [2]), 
      .C2(n_8_0_6007), .ZN(n_8_0_5598));
   NAND2_X1 i_8_0_5828 (.A1(n_8_0_225), .A2(n_8_0_6842), .ZN(n_8_0_5599));
   AOI21_X1 i_8_0_5829 (.A(n_8_0_5601), .B1(n_8_0_6511), .B2(n_8_0_351), 
      .ZN(n_8_0_5600));
   OAI21_X1 i_8_0_5830 (.A(n_8_0_6375), .B1(n_8_0_5602), .B2(\out_bs[5] [4]), 
      .ZN(n_8_0_5601));
   OAI21_X1 i_8_0_5831 (.A(n_8_0_6166), .B1(n_8_0_6824), .B2(n_8_0_351), 
      .ZN(n_8_0_5602));
   AOI221_X1 i_8_0_5832 (.A(n_8_0_5929), .B1(n_8_0_5607), .B2(n_8_0_6795), 
      .C1(n_8_0_5604), .C2(n_8_0_288), .ZN(n_8_0_5603));
   NAND2_X1 i_8_0_5833 (.A1(n_8_0_6557), .A2(n_8_0_5606), .ZN(n_8_0_5604));
   INV_X1 i_8_0_5834 (.A(n_8_0_5606), .ZN(n_8_0_5605));
   NOR2_X1 i_8_0_5835 (.A1(n_8_0_5607), .A2(n_8_0_7034), .ZN(n_8_0_5606));
   NOR2_X1 i_8_0_5836 (.A1(n_8_0_5744), .A2(\out_bs[4] [2]), .ZN(n_8_0_5607));
   NAND4_X1 i_8_0_5837 (.A1(n_8_0_5623), .A2(n_8_0_5613), .A3(n_8_0_5609), 
      .A4(n_8_0_5616), .ZN(n_8_0_5608));
   OAI21_X1 i_8_0_5838 (.A(n_8_0_5610), .B1(n_8_0_5611), .B2(n_8_0_6233), 
      .ZN(n_8_0_5609));
   NAND2_X1 i_8_0_5839 (.A1(n_8_0_5612), .A2(n_8_0_477), .ZN(n_8_0_5610));
   NOR2_X1 i_8_0_5840 (.A1(n_8_0_5612), .A2(n_8_0_477), .ZN(n_8_0_5611));
   OAI21_X1 i_8_0_5841 (.A(n_8_0_6728), .B1(n_8_0_5975), .B2(\out_bs[7] [2]), 
      .ZN(n_8_0_5612));
   OAI21_X1 i_8_0_5842 (.A(n_8_0_5614), .B1(n_8_0_6773), .B2(n_8_0_6954), 
      .ZN(n_8_0_5613));
   OAI22_X1 i_8_0_5843 (.A1(n_8_0_162), .A2(n_8_0_6772), .B1(n_8_0_6711), 
      .B2(n_8_0_5615), .ZN(n_8_0_5614));
   NOR2_X1 i_8_0_5844 (.A1(n_8_0_5814), .A2(\out_bs[2] [2]), .ZN(n_8_0_5615));
   NOR3_X1 i_8_0_5845 (.A1(n_8_0_5619), .A2(n_8_0_5618), .A3(n_8_0_5617), 
      .ZN(n_8_0_5616));
   NOR2_X1 i_8_0_5846 (.A1(n_8_0_36), .A2(n_8_0_6811), .ZN(n_8_0_5617));
   AOI221_X1 i_8_0_5847 (.A(n_8_0_6670), .B1(n_8_0_5944), .B2(n_8_0_7081), 
      .C1(n_8_0_6812), .C2(n_8_0_36), .ZN(n_8_0_5618));
   OAI21_X1 i_8_0_5848 (.A(n_8_0_5620), .B1(n_8_0_6782), .B2(n_8_0_99), .ZN(
      n_8_0_5619));
   INV_X1 i_8_0_5849 (.A(n_8_0_5621), .ZN(n_8_0_5620));
   AOI211_X1 i_8_0_5850 (.A(n_8_0_6693), .B(n_8_0_5622), .C1(n_8_0_6784), 
      .C2(n_8_0_99), .ZN(n_8_0_5621));
   NOR2_X1 i_8_0_5851 (.A1(n_8_0_5983), .A2(\out_bs[1] [2]), .ZN(n_8_0_5622));
   OAI21_X1 i_8_0_5852 (.A(n_8_0_5625), .B1(n_8_0_5624), .B2(n_8_0_6754), 
      .ZN(n_8_0_5623));
   NOR2_X1 i_8_0_5853 (.A1(n_8_0_5626), .A2(n_8_0_6752), .ZN(n_8_0_5624));
   OAI21_X1 i_8_0_5854 (.A(n_8_0_414), .B1(n_8_0_6588), .B2(n_8_0_5626), 
      .ZN(n_8_0_5625));
   NOR2_X1 i_8_0_5855 (.A1(n_8_0_5893), .A2(\out_bs[6] [2]), .ZN(n_8_0_5626));
   AOI21_X1 i_8_0_5856 (.A(n_8_0_6853), .B1(n_8_0_5627), .B2(n_8_0_5632), 
      .ZN(n_166));
   NOR2_X1 i_8_0_5857 (.A1(n_8_0_5634), .A2(n_8_0_5628), .ZN(n_8_0_5627));
   OAI21_X1 i_8_0_5858 (.A(n_8_0_5629), .B1(n_8_0_6837), .B2(n_8_0_226), 
      .ZN(n_8_0_5628));
   OAI21_X1 i_8_0_5859 (.A(n_8_0_5630), .B1(n_8_0_6007), .B2(n_8_0_6565), 
      .ZN(n_8_0_5629));
   AOI21_X1 i_8_0_5860 (.A(n_8_0_6658), .B1(n_8_0_6842), .B2(n_8_0_226), 
      .ZN(n_8_0_5630));
   INV_X1 i_8_0_5861 (.A(n_8_0_5632), .ZN(n_8_0_5631));
   OAI211_X1 i_8_0_5862 (.A(n_8_0_5928), .B(n_8_0_5633), .C1(n_8_0_6915), 
      .C2(n_8_0_6555), .ZN(n_8_0_5632));
   OAI211_X1 i_8_0_5863 (.A(n_8_0_7033), .B(n_8_0_6192), .C1(n_8_0_6795), 
      .C2(n_8_0_289), .ZN(n_8_0_5633));
   NAND4_X1 i_8_0_5864 (.A1(n_8_0_5654), .A2(n_8_0_5639), .A3(n_8_0_5636), 
      .A4(n_8_0_5635), .ZN(n_8_0_5634));
   NOR3_X1 i_8_0_5865 (.A1(n_8_0_5657), .A2(n_8_0_5651), .A3(n_8_0_5648), 
      .ZN(n_8_0_5635));
   AOI21_X1 i_8_0_5866 (.A(n_8_0_5637), .B1(n_8_0_5638), .B2(n_8_0_6671), 
      .ZN(n_8_0_5636));
   OAI21_X1 i_8_0_5867 (.A(n_8_0_5643), .B1(n_8_0_6811), .B2(n_8_0_37), .ZN(
      n_8_0_5637));
   AOI21_X1 i_8_0_5868 (.A(n_8_0_5653), .B1(n_8_0_6812), .B2(n_8_0_37), .ZN(
      n_8_0_5638));
   AOI21_X1 i_8_0_5869 (.A(n_8_0_5640), .B1(n_8_0_5642), .B2(n_8_0_6605), 
      .ZN(n_8_0_5639));
   AOI21_X1 i_8_0_5870 (.A(n_8_0_163), .B1(n_8_0_6772), .B2(n_8_0_5641), 
      .ZN(n_8_0_5640));
   NAND2_X1 i_8_0_5871 (.A1(n_8_0_5642), .A2(n_8_0_6712), .ZN(n_8_0_5641));
   NAND2_X1 i_8_0_5872 (.A1(n_8_0_6537), .A2(n_8_0_5815), .ZN(n_8_0_5642));
   INV_X1 i_8_0_5873 (.A(n_8_0_5644), .ZN(n_8_0_5643));
   AOI21_X1 i_8_0_5874 (.A(n_8_0_5645), .B1(n_8_0_5646), .B2(n_8_0_100), 
      .ZN(n_8_0_5644));
   AOI21_X1 i_8_0_5875 (.A(n_8_0_6781), .B1(n_8_0_6694), .B2(n_8_0_5647), 
      .ZN(n_8_0_5645));
   NAND3_X1 i_8_0_5876 (.A1(n_8_0_6783), .A2(n_8_0_6694), .A3(n_8_0_5647), 
      .ZN(n_8_0_5646));
   NAND2_X1 i_8_0_5877 (.A1(n_8_0_6532), .A2(n_8_0_5984), .ZN(n_8_0_5647));
   INV_X1 i_8_0_5878 (.A(n_8_0_5649), .ZN(n_8_0_5648));
   NAND2_X1 i_8_0_5879 (.A1(n_8_0_6233), .A2(n_8_0_5650), .ZN(n_8_0_5649));
   OAI21_X1 i_8_0_5880 (.A(n_8_0_478), .B1(n_8_0_5652), .B2(n_8_0_6727), 
      .ZN(n_8_0_5650));
   NOR3_X1 i_8_0_5881 (.A1(n_8_0_478), .A2(n_8_0_5652), .A3(n_8_0_6727), 
      .ZN(n_8_0_5651));
   NOR2_X1 i_8_0_5883 (.A1(n_8_0_6522), .A2(n_8_0_5943), .ZN(n_8_0_5653));
   NAND2_X1 i_8_0_5884 (.A1(n_8_0_5656), .A2(n_8_0_5655), .ZN(n_8_0_5654));
   OAI221_X1 i_8_0_5885 (.A(n_8_0_6683), .B1(n_8_0_6211), .B2(n_8_0_6685), 
      .C1(n_8_0_6824), .C2(n_8_0_352), .ZN(n_8_0_5655));
   NAND2_X1 i_8_0_5886 (.A1(n_8_0_6619), .A2(n_8_0_352), .ZN(n_8_0_5656));
   OAI22_X1 i_8_0_5887 (.A1(n_8_0_6752), .A2(n_8_0_5658), .B1(n_8_0_415), 
      .B2(n_8_0_6755), .ZN(n_8_0_5657));
   OAI22_X1 i_8_0_5888 (.A1(n_8_0_6759), .A2(n_8_0_6886), .B1(n_8_0_5893), 
      .B2(n_8_0_6550), .ZN(n_8_0_5658));
   AOI21_X1 i_8_0_5889 (.A(n_8_0_6853), .B1(n_8_0_5659), .B2(n_8_0_5684), 
      .ZN(n_167));
   NOR4_X1 i_8_0_5890 (.A1(n_8_0_5660), .A2(n_8_0_5678), .A3(n_8_0_5683), 
      .A4(n_8_0_5688), .ZN(n_8_0_5659));
   NAND4_X1 i_8_0_5891 (.A1(n_8_0_5675), .A2(n_8_0_5662), .A3(n_8_0_5661), 
      .A4(n_8_0_5670), .ZN(n_8_0_5660));
   AOI21_X1 i_8_0_5892 (.A(n_8_0_5666), .B1(n_8_0_6810), .B2(n_8_0_6984), 
      .ZN(n_8_0_5661));
   OAI21_X1 i_8_0_5893 (.A(n_8_0_5663), .B1(n_8_0_6773), .B2(n_8_0_6952), 
      .ZN(n_8_0_5662));
   OAI22_X1 i_8_0_5894 (.A1(n_8_0_164), .A2(n_8_0_6772), .B1(n_8_0_6711), 
      .B2(n_8_0_5665), .ZN(n_8_0_5663));
   NAND2_X1 i_8_0_5895 (.A1(n_8_0_5815), .A2(n_8_0_6612), .ZN(n_8_0_5664));
   NOR2_X1 i_8_0_5896 (.A1(n_8_0_6613), .A2(n_8_0_5814), .ZN(n_8_0_5665));
   OAI22_X1 i_8_0_5897 (.A1(n_8_0_101), .A2(n_8_0_5667), .B1(n_8_0_5669), 
      .B2(n_8_0_6525), .ZN(n_8_0_5666));
   AOI21_X1 i_8_0_5898 (.A(n_8_0_6781), .B1(n_8_0_6694), .B2(n_8_0_5668), 
      .ZN(n_8_0_5667));
   NAND2_X1 i_8_0_5899 (.A1(n_8_0_5984), .A2(n_8_0_6699), .ZN(n_8_0_5668));
   NOR2_X1 i_8_0_5900 (.A1(n_8_0_6700), .A2(n_8_0_5983), .ZN(n_8_0_5669));
   OAI21_X1 i_8_0_5901 (.A(n_8_0_5671), .B1(n_8_0_5672), .B2(n_8_0_6233), 
      .ZN(n_8_0_5670));
   NAND2_X1 i_8_0_5902 (.A1(n_8_0_5673), .A2(n_8_0_479), .ZN(n_8_0_5671));
   NOR2_X1 i_8_0_5903 (.A1(n_8_0_5673), .A2(n_8_0_479), .ZN(n_8_0_5672));
   NAND2_X1 i_8_0_5904 (.A1(n_8_0_5674), .A2(n_8_0_6728), .ZN(n_8_0_5673));
   AOI22_X1 i_8_0_5906 (.A1(n_8_0_5676), .A2(n_8_0_5677), .B1(n_8_0_6754), 
      .B2(n_8_0_6885), .ZN(n_8_0_5675));
   AOI21_X1 i_8_0_5907 (.A(n_8_0_6752), .B1(n_8_0_6758), .B2(n_8_0_416), 
      .ZN(n_8_0_5676));
   NAND2_X1 i_8_0_5908 (.A1(n_8_0_5894), .A2(n_8_0_6743), .ZN(n_8_0_5677));
   INV_X1 i_8_0_5909 (.A(n_8_0_5679), .ZN(n_8_0_5678));
   NAND3_X1 i_8_0_5910 (.A1(n_8_0_6375), .A2(n_8_0_5681), .A3(n_8_0_5680), 
      .ZN(n_8_0_5679));
   OAI21_X1 i_8_0_5911 (.A(n_8_0_353), .B1(n_8_0_6511), .B2(n_8_0_5682), 
      .ZN(n_8_0_5680));
   NAND2_X1 i_8_0_5912 (.A1(n_8_0_6824), .A2(n_8_0_5682), .ZN(n_8_0_5681));
   NOR2_X1 i_8_0_5913 (.A1(n_8_0_6300), .A2(\out_bs[5] [4]), .ZN(n_8_0_5682));
   AOI221_X1 i_8_0_5914 (.A(n_8_0_6595), .B1(n_8_0_6247), .B2(n_8_0_38), 
      .C1(n_8_0_5944), .C2(n_8_0_6667), .ZN(n_8_0_5683));
   OAI211_X1 i_8_0_5915 (.A(n_8_0_6571), .B(n_8_0_5685), .C1(n_8_0_5687), 
      .C2(n_8_0_6838), .ZN(n_8_0_5684));
   OAI21_X1 i_8_0_5916 (.A(n_8_0_227), .B1(n_8_0_6575), .B2(n_8_0_5686), 
      .ZN(n_8_0_5685));
   INV_X1 i_8_0_5917 (.A(n_8_0_5687), .ZN(n_8_0_5686));
   NAND2_X1 i_8_0_5918 (.A1(n_8_0_6008), .A2(n_8_0_6652), .ZN(n_8_0_5687));
   OAI22_X1 i_8_0_5919 (.A1(n_8_0_290), .A2(n_8_0_5689), .B1(n_8_0_5691), 
      .B2(n_8_0_6554), .ZN(n_8_0_5688));
   AOI21_X1 i_8_0_5920 (.A(n_8_0_6794), .B1(n_8_0_6636), .B2(n_8_0_5690), 
      .ZN(n_8_0_5689));
   NAND2_X1 i_8_0_5921 (.A1(n_8_0_5745), .A2(n_8_0_6642), .ZN(n_8_0_5690));
   NOR2_X1 i_8_0_5922 (.A1(n_8_0_6643), .A2(n_8_0_5744), .ZN(n_8_0_5691));
   AOI21_X1 i_8_0_5923 (.A(n_8_0_6853), .B1(n_8_0_5692), .B2(n_8_0_5725), 
      .ZN(n_168));
   NOR4_X1 i_8_0_5924 (.A1(n_8_0_5699), .A2(n_8_0_5693), .A3(n_8_0_5718), 
      .A4(n_8_0_5703), .ZN(n_8_0_5692));
   AOI21_X1 i_8_0_5925 (.A(n_8_0_5694), .B1(n_8_0_5695), .B2(n_8_0_228), 
      .ZN(n_8_0_5693));
   AOI21_X1 i_8_0_5926 (.A(n_8_0_6838), .B1(n_8_0_6659), .B2(n_8_0_5697), 
      .ZN(n_8_0_5694));
   NAND2_X1 i_8_0_5927 (.A1(n_8_0_6576), .A2(n_8_0_5697), .ZN(n_8_0_5695));
   INV_X1 i_8_0_5928 (.A(n_8_0_5697), .ZN(n_8_0_5696));
   NAND2_X1 i_8_0_5929 (.A1(n_8_0_6649), .A2(n_8_0_6008), .ZN(n_8_0_5697));
   NOR2_X1 i_8_0_5930 (.A1(\out_bs[3] [3]), .A2(n_8_0_6650), .ZN(n_8_0_5698));
   AOI21_X1 i_8_0_5931 (.A(n_8_0_5700), .B1(n_8_0_6824), .B2(n_8_0_354), 
      .ZN(n_8_0_5699));
   INV_X1 i_8_0_5932 (.A(n_8_0_5701), .ZN(n_8_0_5700));
   OAI22_X1 i_8_0_5933 (.A1(n_8_0_354), .A2(n_8_0_6824), .B1(n_8_0_6685), 
      .B2(n_8_0_5702), .ZN(n_8_0_5701));
   NOR2_X1 i_8_0_5934 (.A1(\out_bs[5] [4]), .A2(n_8_0_6299), .ZN(n_8_0_5702));
   NAND4_X1 i_8_0_5935 (.A1(n_8_0_5717), .A2(n_8_0_5704), .A3(n_8_0_5712), 
      .A4(n_8_0_5708), .ZN(n_8_0_5703));
   OAI21_X1 i_8_0_5936 (.A(n_8_0_5705), .B1(n_8_0_6773), .B2(n_8_0_6951), 
      .ZN(n_8_0_5704));
   OAI22_X1 i_8_0_5937 (.A1(n_8_0_165), .A2(n_8_0_6772), .B1(n_8_0_6711), 
      .B2(n_8_0_5707), .ZN(n_8_0_5705));
   OAI21_X1 i_8_0_5938 (.A(n_8_0_5815), .B1(n_8_0_6612), .B2(n_8_0_7054), 
      .ZN(n_8_0_5706));
   AOI21_X1 i_8_0_5939 (.A(n_8_0_5814), .B1(n_8_0_6613), .B2(\out_bs[2] [0]), 
      .ZN(n_8_0_5707));
   OAI21_X1 i_8_0_5940 (.A(n_8_0_5709), .B1(n_8_0_5710), .B2(n_8_0_5711), 
      .ZN(n_8_0_5708));
   AOI21_X1 i_8_0_5941 (.A(n_8_0_6265), .B1(n_8_0_6525), .B2(n_8_0_102), 
      .ZN(n_8_0_5709));
   NOR2_X1 i_8_0_5942 (.A1(n_8_0_102), .A2(n_8_0_6782), .ZN(n_8_0_5710));
   NAND2_X1 i_8_0_5943 (.A1(n_8_0_6697), .A2(n_8_0_5984), .ZN(n_8_0_5711));
   OAI21_X1 i_8_0_5944 (.A(n_8_0_5713), .B1(n_8_0_5714), .B2(n_8_0_6233), 
      .ZN(n_8_0_5712));
   NAND2_X1 i_8_0_5945 (.A1(n_8_0_5715), .A2(n_8_0_480), .ZN(n_8_0_5713));
   NOR2_X1 i_8_0_5946 (.A1(n_8_0_5715), .A2(n_8_0_480), .ZN(n_8_0_5714));
   NAND2_X1 i_8_0_5947 (.A1(n_8_0_5716), .A2(n_8_0_6728), .ZN(n_8_0_5715));
   NAND2_X1 i_8_0_5948 (.A1(n_8_0_6722), .A2(n_8_0_5976), .ZN(n_8_0_5716));
   NAND2_X1 i_8_0_5949 (.A1(n_8_0_6248), .A2(n_8_0_5724), .ZN(n_8_0_5717));
   OAI21_X1 i_8_0_5950 (.A(n_8_0_5720), .B1(n_8_0_5723), .B2(n_8_0_39), .ZN(
      n_8_0_5718));
   INV_X1 i_8_0_5951 (.A(n_8_0_5720), .ZN(n_8_0_5719));
   AOI22_X1 i_8_0_5952 (.A1(n_8_0_5721), .A2(n_8_0_5722), .B1(n_8_0_6754), 
      .B2(n_8_0_6884), .ZN(n_8_0_5720));
   AOI21_X1 i_8_0_5953 (.A(n_8_0_6752), .B1(n_8_0_6758), .B2(n_8_0_417), 
      .ZN(n_8_0_5721));
   OAI21_X1 i_8_0_5954 (.A(n_8_0_5894), .B1(n_8_0_6743), .B2(n_8_0_7006), 
      .ZN(n_8_0_5722));
   AOI21_X1 i_8_0_5955 (.A(n_8_0_6810), .B1(n_8_0_6671), .B2(n_8_0_5724), 
      .ZN(n_8_0_5723));
   OAI211_X1 i_8_0_5957 (.A(n_8_0_5928), .B(n_8_0_5726), .C1(n_8_0_5728), 
      .C2(n_8_0_6794), .ZN(n_8_0_5725));
   OAI21_X1 i_8_0_5958 (.A(n_8_0_291), .B1(n_8_0_6554), .B2(n_8_0_5727), 
      .ZN(n_8_0_5726));
   INV_X1 i_8_0_5959 (.A(n_8_0_5728), .ZN(n_8_0_5727));
   NAND2_X1 i_8_0_5960 (.A1(n_8_0_6629), .A2(n_8_0_5745), .ZN(n_8_0_5728));
   AOI21_X1 i_8_0_5961 (.A(n_8_0_6853), .B1(n_8_0_5741), .B2(n_8_0_5729), 
      .ZN(n_169));
   NOR4_X1 i_8_0_5962 (.A1(n_8_0_5738), .A2(n_8_0_5730), .A3(n_8_0_5737), 
      .A4(n_8_0_5735), .ZN(n_8_0_5729));
   OAI211_X1 i_8_0_5963 (.A(n_8_0_5733), .B(n_8_0_5731), .C1(n_8_0_6247), 
      .C2(n_8_0_5944), .ZN(n_8_0_5730));
   OAI211_X1 i_8_0_5964 (.A(n_8_0_6264), .B(n_8_0_5732), .C1(n_8_0_5983), 
      .C2(n_8_0_6781), .ZN(n_8_0_5731));
   OAI21_X1 i_8_0_5965 (.A(n_8_0_103), .B1(n_8_0_6525), .B2(n_8_0_5984), 
      .ZN(n_8_0_5732));
   OAI21_X1 i_8_0_5966 (.A(n_8_0_5734), .B1(n_8_0_6773), .B2(n_8_0_6950), 
      .ZN(n_8_0_5733));
   OAI22_X1 i_8_0_5967 (.A1(n_8_0_166), .A2(n_8_0_6772), .B1(n_8_0_6711), 
      .B2(n_8_0_5815), .ZN(n_8_0_5734));
   OAI22_X1 i_8_0_5968 (.A1(n_8_0_481), .A2(n_8_0_5736), .B1(n_8_0_5976), 
      .B2(n_8_0_6464), .ZN(n_8_0_5735));
   AOI21_X1 i_8_0_5969 (.A(n_8_0_6729), .B1(n_8_0_6728), .B2(n_8_0_5975), 
      .ZN(n_8_0_5736));
   AOI211_X1 i_8_0_5970 (.A(n_8_0_40), .B(n_8_0_6595), .C1(n_8_0_5944), .C2(
      n_8_0_6811), .ZN(n_8_0_5737));
   AOI21_X1 i_8_0_5971 (.A(n_8_0_5739), .B1(n_8_0_5740), .B2(n_8_0_229), 
      .ZN(n_8_0_5738));
   AOI21_X1 i_8_0_5972 (.A(n_8_0_6838), .B1(n_8_0_6659), .B2(n_8_0_6007), 
      .ZN(n_8_0_5739));
   NAND2_X1 i_8_0_5973 (.A1(n_8_0_6576), .A2(n_8_0_6007), .ZN(n_8_0_5740));
   NOR3_X1 i_8_0_5974 (.A1(n_8_0_5749), .A2(n_8_0_5746), .A3(n_8_0_5742), 
      .ZN(n_8_0_5741));
   OAI22_X1 i_8_0_5975 (.A1(n_8_0_292), .A2(n_8_0_5743), .B1(n_8_0_5745), 
      .B2(n_8_0_6554), .ZN(n_8_0_5742));
   AOI21_X1 i_8_0_5976 (.A(n_8_0_6794), .B1(n_8_0_6636), .B2(n_8_0_5744), 
      .ZN(n_8_0_5743));
   NAND2_X1 i_8_0_5977 (.A1(n_8_0_7033), .A2(n_8_0_7032), .ZN(n_8_0_5744));
   NOR2_X1 i_8_0_5978 (.A1(\out_bs[4] [4]), .A2(\out_bs[4] [3]), .ZN(n_8_0_5745));
   AOI221_X1 i_8_0_5979 (.A(n_8_0_6376), .B1(n_8_0_5748), .B2(n_8_0_6824), 
      .C1(n_8_0_5747), .C2(n_8_0_355), .ZN(n_8_0_5746));
   OAI21_X1 i_8_0_5980 (.A(n_8_0_6512), .B1(\out_bs[5] [3]), .B2(\out_bs[5] [4]), 
      .ZN(n_8_0_5747));
   NOR2_X1 i_8_0_5981 (.A1(\out_bs[5] [4]), .A2(\out_bs[5] [3]), .ZN(n_8_0_5748));
   AOI21_X1 i_8_0_5982 (.A(n_8_0_5750), .B1(n_8_0_5751), .B2(n_8_0_418), 
      .ZN(n_8_0_5749));
   AOI21_X1 i_8_0_5983 (.A(n_8_0_6754), .B1(n_8_0_6753), .B2(n_8_0_5893), 
      .ZN(n_8_0_5750));
   NAND2_X1 i_8_0_5984 (.A1(n_8_0_6589), .A2(n_8_0_5893), .ZN(n_8_0_5751));
   NOR2_X1 i_8_0_5985 (.A1(n_8_0_5752), .A2(n_8_0_6853), .ZN(n_170));
   NOR3_X1 i_8_0_5986 (.A1(n_8_0_5776), .A2(n_8_0_5754), .A3(n_8_0_5753), 
      .ZN(n_8_0_5752));
   OAI21_X1 i_8_0_5987 (.A(n_8_0_5772), .B1(n_8_0_5770), .B2(n_8_0_5769), 
      .ZN(n_8_0_5753));
   NAND3_X1 i_8_0_5988 (.A1(n_8_0_5765), .A2(n_8_0_5759), .A3(n_8_0_5755), 
      .ZN(n_8_0_5754));
   NAND2_X1 i_8_0_5989 (.A1(n_8_0_5756), .A2(n_8_0_5757), .ZN(n_8_0_5755));
   OAI21_X1 i_8_0_5990 (.A(n_8_0_6782), .B1(n_8_0_6693), .B2(n_8_0_5758), 
      .ZN(n_8_0_5756));
   OAI21_X1 i_8_0_5991 (.A(n_8_0_104), .B1(n_8_0_6525), .B2(n_8_0_5758), 
      .ZN(n_8_0_5757));
   NOR2_X1 i_8_0_5992 (.A1(\out_bs[1] [4]), .A2(n_8_0_6341), .ZN(n_8_0_5758));
   OAI21_X1 i_8_0_5993 (.A(n_8_0_5760), .B1(n_8_0_5762), .B2(n_8_0_6233), 
      .ZN(n_8_0_5759));
   OAI21_X1 i_8_0_5994 (.A(n_8_0_482), .B1(n_8_0_6232), .B2(n_8_0_5761), 
      .ZN(n_8_0_5760));
   INV_X1 i_8_0_5995 (.A(n_8_0_5762), .ZN(n_8_0_5761));
   NOR2_X1 i_8_0_5996 (.A1(n_8_0_5764), .A2(n_8_0_6727), .ZN(n_8_0_5762));
   INV_X1 i_8_0_5997 (.A(n_8_0_5764), .ZN(n_8_0_5763));
   NOR2_X1 i_8_0_5998 (.A1(\out_bs[7] [4]), .A2(n_8_0_6362), .ZN(n_8_0_5764));
   AOI22_X1 i_8_0_5999 (.A1(n_8_0_6753), .A2(n_8_0_5766), .B1(n_8_0_6883), 
      .B2(n_8_0_6754), .ZN(n_8_0_5765));
   AOI21_X1 i_8_0_6000 (.A(n_8_0_5768), .B1(n_8_0_6758), .B2(n_8_0_419), 
      .ZN(n_8_0_5766));
   OR2_X1 i_8_0_6001 (.A1(\out_bs[6] [4]), .A2(n_8_0_6368), .ZN(n_8_0_5767));
   NOR2_X1 i_8_0_6002 (.A1(\out_bs[6] [4]), .A2(n_8_0_6368), .ZN(n_8_0_5768));
   AOI21_X1 i_8_0_6003 (.A(n_8_0_6810), .B1(n_8_0_6671), .B2(n_8_0_5771), 
      .ZN(n_8_0_5769));
   AOI21_X1 i_8_0_6004 (.A(n_8_0_6983), .B1(n_8_0_6248), .B2(n_8_0_5771), 
      .ZN(n_8_0_5770));
   AOI21_X1 i_8_0_6005 (.A(n_8_0_5944), .B1(n_8_0_6345), .B2(n_8_0_7083), 
      .ZN(n_8_0_5771));
   NAND2_X1 i_8_0_6006 (.A1(n_8_0_5774), .A2(n_8_0_5773), .ZN(n_8_0_5772));
   OAI21_X1 i_8_0_6007 (.A(n_8_0_6824), .B1(n_8_0_6685), .B2(n_8_0_5775), 
      .ZN(n_8_0_5773));
   OAI21_X1 i_8_0_6008 (.A(n_8_0_356), .B1(n_8_0_6511), .B2(n_8_0_5775), 
      .ZN(n_8_0_5774));
   NOR2_X1 i_8_0_6009 (.A1(n_8_0_6374), .A2(\out_bs[5] [4]), .ZN(n_8_0_5775));
   NAND3_X1 i_8_0_6010 (.A1(n_8_0_5784), .A2(n_8_0_5780), .A3(n_8_0_5777), 
      .ZN(n_8_0_5776));
   OAI21_X1 i_8_0_6011 (.A(n_8_0_5778), .B1(n_8_0_6773), .B2(n_8_0_6949), 
      .ZN(n_8_0_5777));
   OAI22_X1 i_8_0_6012 (.A1(n_8_0_167), .A2(n_8_0_6772), .B1(n_8_0_6711), 
      .B2(n_8_0_5779), .ZN(n_8_0_5778));
   AOI21_X1 i_8_0_6013 (.A(\out_bs[2] [4]), .B1(n_8_0_6335), .B2(\out_bs[2] [3]), 
      .ZN(n_8_0_5779));
   OAI211_X1 i_8_0_6014 (.A(n_8_0_5928), .B(n_8_0_5781), .C1(n_8_0_5782), 
      .C2(n_8_0_6794), .ZN(n_8_0_5780));
   OAI21_X1 i_8_0_6015 (.A(n_8_0_293), .B1(n_8_0_6554), .B2(n_8_0_5783), 
      .ZN(n_8_0_5781));
   NAND2_X1 i_8_0_6016 (.A1(n_8_0_7033), .A2(n_8_0_6350), .ZN(n_8_0_5782));
   NOR2_X1 i_8_0_6017 (.A1(\out_bs[4] [4]), .A2(n_8_0_6351), .ZN(n_8_0_5783));
   OAI21_X1 i_8_0_6018 (.A(n_8_0_5786), .B1(n_8_0_5785), .B2(n_8_0_6838), 
      .ZN(n_8_0_5784));
   NOR2_X1 i_8_0_6019 (.A1(n_8_0_5788), .A2(n_8_0_6658), .ZN(n_8_0_5785));
   OAI21_X1 i_8_0_6020 (.A(n_8_0_230), .B1(n_8_0_6575), .B2(n_8_0_5788), 
      .ZN(n_8_0_5786));
   INV_X1 i_8_0_6021 (.A(n_8_0_5788), .ZN(n_8_0_5787));
   AOI21_X1 i_8_0_6022 (.A(\out_bs[3] [4]), .B1(n_8_0_6357), .B2(\out_bs[3] [3]), 
      .ZN(n_8_0_5788));
   AOI21_X1 i_8_0_6023 (.A(n_8_0_6853), .B1(n_8_0_5790), .B2(n_8_0_5789), 
      .ZN(n_171));
   NOR4_X1 i_8_0_6024 (.A1(n_8_0_5820), .A2(n_8_0_5794), .A3(n_8_0_5806), 
      .A4(n_8_0_5800), .ZN(n_8_0_5789));
   NOR4_X1 i_8_0_6025 (.A1(n_8_0_5816), .A2(n_8_0_5811), .A3(n_8_0_5797), 
      .A4(n_8_0_5791), .ZN(n_8_0_5790));
   OAI21_X1 i_8_0_6026 (.A(n_8_0_5792), .B1(n_8_0_6837), .B2(n_8_0_231), 
      .ZN(n_8_0_5791));
   OAI211_X1 i_8_0_6027 (.A(n_8_0_6659), .B(n_8_0_5793), .C1(n_8_0_6843), 
      .C2(n_8_0_6924), .ZN(n_8_0_5792));
   OAI21_X1 i_8_0_6028 (.A(n_8_0_7045), .B1(n_8_0_6414), .B2(n_8_0_7044), 
      .ZN(n_8_0_5793));
   AOI221_X1 i_8_0_6029 (.A(n_8_0_6376), .B1(n_8_0_6511), .B2(n_8_0_357), 
      .C1(n_8_0_7022), .C2(n_8_0_5795), .ZN(n_8_0_5794));
   INV_X1 i_8_0_6030 (.A(n_8_0_5796), .ZN(n_8_0_5795));
   OAI21_X1 i_8_0_6031 (.A(n_8_0_6408), .B1(n_8_0_6824), .B2(n_8_0_357), 
      .ZN(n_8_0_5796));
   OAI21_X1 i_8_0_6032 (.A(n_8_0_5798), .B1(n_8_0_6795), .B2(n_8_0_294), 
      .ZN(n_8_0_5797));
   OAI211_X1 i_8_0_6033 (.A(n_8_0_6636), .B(n_8_0_5799), .C1(n_8_0_6796), 
      .C2(n_8_0_6914), .ZN(n_8_0_5798));
   OR2_X1 i_8_0_6034 (.A1(\out_bs[4] [4]), .A2(n_8_0_6381), .ZN(n_8_0_5799));
   AOI21_X1 i_8_0_6035 (.A(n_8_0_5801), .B1(n_8_0_5802), .B2(n_8_0_42), .ZN(
      n_8_0_5800));
   AOI21_X1 i_8_0_6036 (.A(n_8_0_6810), .B1(n_8_0_6671), .B2(n_8_0_5805), 
      .ZN(n_8_0_5801));
   NAND2_X1 i_8_0_6037 (.A1(n_8_0_6248), .A2(n_8_0_5805), .ZN(n_8_0_5802));
   NAND2_X1 i_8_0_6038 (.A1(n_8_0_5943), .A2(\out_bs[0] [6]), .ZN(n_8_0_5803));
   INV_X1 i_8_0_6039 (.A(n_8_0_5805), .ZN(n_8_0_5804));
   OAI21_X1 i_8_0_6040 (.A(n_8_0_7083), .B1(n_8_0_6421), .B2(n_8_0_7082), 
      .ZN(n_8_0_5805));
   AOI21_X1 i_8_0_6041 (.A(n_8_0_5807), .B1(n_8_0_5808), .B2(n_8_0_6232), 
      .ZN(n_8_0_5806));
   AND2_X1 i_8_0_6042 (.A1(n_8_0_483), .A2(n_8_0_5809), .ZN(n_8_0_5807));
   OR2_X1 i_8_0_6043 (.A1(n_8_0_483), .A2(n_8_0_5809), .ZN(n_8_0_5808));
   OAI21_X1 i_8_0_6044 (.A(n_8_0_6728), .B1(n_8_0_6404), .B2(\out_bs[7] [4]), 
      .ZN(n_8_0_5809));
   INV_X1 i_8_0_6045 (.A(n_8_0_5811), .ZN(n_8_0_5810));
   AOI21_X1 i_8_0_6046 (.A(n_8_0_5812), .B1(n_8_0_6772), .B2(n_8_0_168), 
      .ZN(n_8_0_5811));
   AOI22_X1 i_8_0_6047 (.A1(n_8_0_6948), .A2(n_8_0_6773), .B1(n_8_0_6712), 
      .B2(n_8_0_5813), .ZN(n_8_0_5812));
   OAI21_X1 i_8_0_6048 (.A(n_8_0_7058), .B1(n_8_0_6400), .B2(n_8_0_7057), 
      .ZN(n_8_0_5813));
   NAND2_X1 i_8_0_6049 (.A1(n_8_0_7058), .A2(n_8_0_7057), .ZN(n_8_0_5814));
   NOR2_X1 i_8_0_6050 (.A1(\out_bs[2] [4]), .A2(\out_bs[2] [3]), .ZN(n_8_0_5815));
   OAI22_X1 i_8_0_6051 (.A1(n_8_0_105), .A2(n_8_0_6782), .B1(n_8_0_6693), 
      .B2(n_8_0_5817), .ZN(n_8_0_5816));
   INV_X1 i_8_0_6052 (.A(n_8_0_5818), .ZN(n_8_0_5817));
   AOI21_X1 i_8_0_6053 (.A(n_8_0_5819), .B1(n_8_0_6784), .B2(n_8_0_105), 
      .ZN(n_8_0_5818));
   AOI21_X1 i_8_0_6054 (.A(\out_bs[1] [4]), .B1(n_8_0_6394), .B2(\out_bs[1] [3]), 
      .ZN(n_8_0_5819));
   OAI21_X1 i_8_0_6055 (.A(n_8_0_5821), .B1(n_8_0_6755), .B2(n_8_0_420), 
      .ZN(n_8_0_5820));
   INV_X1 i_8_0_6056 (.A(n_8_0_5822), .ZN(n_8_0_5821));
   AOI211_X1 i_8_0_6057 (.A(n_8_0_6752), .B(n_8_0_5823), .C1(n_8_0_6758), 
      .C2(n_8_0_420), .ZN(n_8_0_5822));
   AOI21_X1 i_8_0_6058 (.A(\out_bs[6] [4]), .B1(n_8_0_6386), .B2(\out_bs[6] [3]), 
      .ZN(n_8_0_5823));
   AOI21_X1 i_8_0_6059 (.A(n_8_0_6853), .B1(n_8_0_5824), .B2(n_8_0_5855), 
      .ZN(n_172));
   NOR4_X1 i_8_0_6060 (.A1(n_8_0_5837), .A2(n_8_0_5832), .A3(n_8_0_5829), 
      .A4(n_8_0_5825), .ZN(n_8_0_5824));
   OAI21_X1 i_8_0_6061 (.A(n_8_0_5826), .B1(n_8_0_6755), .B2(n_8_0_421), 
      .ZN(n_8_0_5825));
   OAI211_X1 i_8_0_6062 (.A(n_8_0_6753), .B(n_8_0_5827), .C1(n_8_0_6759), 
      .C2(n_8_0_6882), .ZN(n_8_0_5826));
   INV_X1 i_8_0_6063 (.A(n_8_0_5828), .ZN(n_8_0_5827));
   AOI21_X1 i_8_0_6064 (.A(\out_bs[6] [4]), .B1(n_8_0_6480), .B2(\out_bs[6] [3]), 
      .ZN(n_8_0_5828));
   OAI22_X1 i_8_0_6065 (.A1(n_8_0_6685), .A2(n_8_0_5830), .B1(n_8_0_358), 
      .B2(n_8_0_6824), .ZN(n_8_0_5829));
   OAI21_X1 i_8_0_6066 (.A(n_8_0_5831), .B1(n_8_0_6460), .B2(\out_bs[5] [4]), 
      .ZN(n_8_0_5830));
   NAND2_X1 i_8_0_6067 (.A1(n_8_0_6824), .A2(n_8_0_358), .ZN(n_8_0_5831));
   AOI21_X1 i_8_0_6068 (.A(n_8_0_5833), .B1(n_8_0_5834), .B2(n_8_0_295), 
      .ZN(n_8_0_5832));
   AOI21_X1 i_8_0_6069 (.A(n_8_0_6794), .B1(n_8_0_6636), .B2(n_8_0_5835), 
      .ZN(n_8_0_5833));
   NAND2_X1 i_8_0_6070 (.A1(n_8_0_6555), .A2(n_8_0_5835), .ZN(n_8_0_5834));
   OR2_X1 i_8_0_6071 (.A1(\out_bs[4] [4]), .A2(n_8_0_6434), .ZN(n_8_0_5835));
   NOR2_X1 i_8_0_6072 (.A1(\out_bs[4] [4]), .A2(n_8_0_6434), .ZN(n_8_0_5836));
   NAND3_X1 i_8_0_6073 (.A1(n_8_0_5838), .A2(n_8_0_5847), .A3(n_8_0_5851), 
      .ZN(n_8_0_5837));
   AOI211_X1 i_8_0_6074 (.A(n_8_0_5843), .B(n_8_0_5840), .C1(n_8_0_5839), 
      .C2(n_8_0_6233), .ZN(n_8_0_5838));
   NAND2_X1 i_8_0_6075 (.A1(n_8_0_5841), .A2(n_8_0_484), .ZN(n_8_0_5839));
   NOR2_X1 i_8_0_6076 (.A1(n_8_0_5841), .A2(n_8_0_484), .ZN(n_8_0_5840));
   NAND2_X1 i_8_0_6077 (.A1(n_8_0_5842), .A2(n_8_0_6728), .ZN(n_8_0_5841));
   AOI21_X1 i_8_0_6079 (.A(n_8_0_5844), .B1(n_8_0_6772), .B2(n_8_0_169), 
      .ZN(n_8_0_5843));
   INV_X1 i_8_0_6080 (.A(n_8_0_5845), .ZN(n_8_0_5844));
   OAI22_X1 i_8_0_6081 (.A1(n_8_0_169), .A2(n_8_0_6772), .B1(n_8_0_6711), 
      .B2(n_8_0_5846), .ZN(n_8_0_5845));
   AND2_X1 i_8_0_6082 (.A1(n_8_0_7058), .A2(n_8_0_6452), .ZN(n_8_0_5846));
   OAI211_X1 i_8_0_6083 (.A(n_8_0_6264), .B(n_8_0_5848), .C1(n_8_0_5850), 
      .C2(n_8_0_6781), .ZN(n_8_0_5847));
   OAI21_X1 i_8_0_6084 (.A(n_8_0_106), .B1(n_8_0_6525), .B2(n_8_0_5849), 
      .ZN(n_8_0_5848));
   AOI21_X1 i_8_0_6085 (.A(\out_bs[1] [4]), .B1(n_8_0_6447), .B2(\out_bs[1] [3]), 
      .ZN(n_8_0_5849));
   AOI21_X1 i_8_0_6086 (.A(n_8_0_5984), .B1(n_8_0_5982), .B2(n_8_0_6690), 
      .ZN(n_8_0_5850));
   NAND2_X1 i_8_0_6087 (.A1(n_8_0_5853), .A2(n_8_0_5852), .ZN(n_8_0_5851));
   OAI21_X1 i_8_0_6088 (.A(n_8_0_43), .B1(n_8_0_6247), .B2(n_8_0_5854), .ZN(
      n_8_0_5852));
   OAI21_X1 i_8_0_6089 (.A(n_8_0_6811), .B1(n_8_0_6670), .B2(n_8_0_5854), 
      .ZN(n_8_0_5853));
   AOI21_X1 i_8_0_6090 (.A(\out_bs[0] [4]), .B1(n_8_0_6441), .B2(\out_bs[0] [3]), 
      .ZN(n_8_0_5854));
   OAI21_X1 i_8_0_6091 (.A(n_8_0_5857), .B1(n_8_0_5856), .B2(n_8_0_6838), 
      .ZN(n_8_0_5855));
   NOR2_X1 i_8_0_6092 (.A1(n_8_0_5859), .A2(n_8_0_6658), .ZN(n_8_0_5856));
   OAI21_X1 i_8_0_6093 (.A(n_8_0_232), .B1(n_8_0_6575), .B2(n_8_0_5859), 
      .ZN(n_8_0_5857));
   OAI21_X1 i_8_0_6094 (.A(n_8_0_7045), .B1(n_8_0_6429), .B2(n_8_0_7044), 
      .ZN(n_8_0_5858));
   NOR2_X1 i_8_0_6095 (.A1(\out_bs[3] [4]), .A2(n_8_0_6427), .ZN(n_8_0_5859));
   AOI21_X1 i_8_0_6096 (.A(n_8_0_6853), .B1(n_8_0_5860), .B2(n_8_0_5879), 
      .ZN(n_173));
   NOR3_X1 i_8_0_6097 (.A1(n_8_0_5866), .A2(n_8_0_5862), .A3(n_8_0_5861), 
      .ZN(n_8_0_5860));
   NAND4_X1 i_8_0_6098 (.A1(n_8_0_5874), .A2(n_8_0_5872), .A3(n_8_0_5869), 
      .A4(n_8_0_5882), .ZN(n_8_0_5861));
   AOI221_X1 i_8_0_6099 (.A(n_8_0_6572), .B1(n_8_0_5863), .B2(n_8_0_233), 
      .C1(n_8_0_5865), .C2(n_8_0_6837), .ZN(n_8_0_5862));
   NAND2_X1 i_8_0_6100 (.A1(n_8_0_6576), .A2(n_8_0_5864), .ZN(n_8_0_5863));
   OAI21_X1 i_8_0_6101 (.A(n_8_0_7045), .B1(n_8_0_7044), .B2(n_8_0_7043), 
      .ZN(n_8_0_5864));
   AOI21_X1 i_8_0_6102 (.A(\out_bs[3] [4]), .B1(\out_bs[3] [3]), .B2(
      \out_bs[3] [2]), .ZN(n_8_0_5865));
   AOI211_X1 i_8_0_6103 (.A(n_8_0_6376), .B(n_8_0_5867), .C1(n_8_0_359), 
      .C2(n_8_0_6511), .ZN(n_8_0_5866));
   NOR2_X1 i_8_0_6104 (.A1(n_8_0_5868), .A2(\out_bs[5] [4]), .ZN(n_8_0_5867));
   OAI21_X1 i_8_0_6105 (.A(n_8_0_6678), .B1(n_8_0_6824), .B2(n_8_0_359), 
      .ZN(n_8_0_5868));
   OAI21_X1 i_8_0_6106 (.A(n_8_0_5870), .B1(n_8_0_6796), .B2(n_8_0_6913), 
      .ZN(n_8_0_5869));
   OAI22_X1 i_8_0_6107 (.A1(n_8_0_296), .A2(n_8_0_6795), .B1(n_8_0_6635), 
      .B2(n_8_0_5871), .ZN(n_8_0_5870));
   AOI21_X1 i_8_0_6108 (.A(\out_bs[4] [4]), .B1(\out_bs[4] [3]), .B2(
      \out_bs[4] [2]), .ZN(n_8_0_5871));
   OAI21_X1 i_8_0_6109 (.A(n_8_0_5873), .B1(n_8_0_6759), .B2(n_8_0_6881), 
      .ZN(n_8_0_5872));
   OAI22_X1 i_8_0_6110 (.A1(n_8_0_422), .A2(n_8_0_6755), .B1(n_8_0_6752), 
      .B2(n_8_0_5970), .ZN(n_8_0_5873));
   AOI211_X1 i_8_0_6111 (.A(n_8_0_5877), .B(n_8_0_5875), .C1(n_8_0_6233), 
      .C2(n_8_0_5878), .ZN(n_8_0_5874));
   OAI22_X1 i_8_0_6112 (.A1(n_8_0_107), .A2(n_8_0_5876), .B1(n_8_0_5980), 
      .B2(n_8_0_6525), .ZN(n_8_0_5875));
   AOI21_X1 i_8_0_6113 (.A(n_8_0_6781), .B1(n_8_0_6694), .B2(n_8_0_5981), 
      .ZN(n_8_0_5876));
   NOR3_X1 i_8_0_6114 (.A1(n_8_0_485), .A2(n_8_0_5954), .A3(n_8_0_6727), 
      .ZN(n_8_0_5877));
   OAI21_X1 i_8_0_6115 (.A(n_8_0_485), .B1(n_8_0_5954), .B2(n_8_0_6727), 
      .ZN(n_8_0_5878));
   NAND2_X1 i_8_0_6116 (.A1(n_8_0_5881), .A2(n_8_0_5880), .ZN(n_8_0_5879));
   OAI21_X1 i_8_0_6117 (.A(n_8_0_6772), .B1(n_8_0_6711), .B2(n_8_0_5991), 
      .ZN(n_8_0_5880));
   OAI21_X1 i_8_0_6118 (.A(n_8_0_170), .B1(n_8_0_6604), .B2(n_8_0_5991), 
      .ZN(n_8_0_5881));
   OAI211_X1 i_8_0_6119 (.A(n_8_0_6594), .B(n_8_0_5883), .C1(n_8_0_5942), 
      .C2(n_8_0_6810), .ZN(n_8_0_5882));
   OAI21_X1 i_8_0_6120 (.A(n_8_0_44), .B1(n_8_0_6247), .B2(n_8_0_5941), .ZN(
      n_8_0_5883));
   AOI21_X1 i_8_0_6121 (.A(n_8_0_6853), .B1(n_8_0_5886), .B2(n_8_0_5884), 
      .ZN(n_174));
   NOR4_X1 i_8_0_6122 (.A1(n_8_0_5919), .A2(n_8_0_5915), .A3(n_8_0_5887), 
      .A4(n_8_0_5885), .ZN(n_8_0_5884));
   OAI21_X1 i_8_0_6123 (.A(n_8_0_5898), .B1(n_8_0_5908), .B2(n_8_0_6247), 
      .ZN(n_8_0_5885));
   NOR4_X1 i_8_0_6124 (.A1(n_8_0_5903), .A2(n_8_0_5895), .A3(n_8_0_5888), 
      .A4(n_8_0_5909), .ZN(n_8_0_5886));
   AOI211_X1 i_8_0_6125 (.A(n_8_0_45), .B(n_8_0_6595), .C1(n_8_0_5908), .C2(
      n_8_0_6811), .ZN(n_8_0_5887));
   AND2_X1 i_8_0_6126 (.A1(n_8_0_5890), .A2(n_8_0_5889), .ZN(n_8_0_5888));
   OAI21_X1 i_8_0_6127 (.A(n_8_0_6755), .B1(n_8_0_6752), .B2(n_8_0_5892), 
      .ZN(n_8_0_5889));
   OAI21_X1 i_8_0_6128 (.A(n_8_0_423), .B1(n_8_0_6588), .B2(n_8_0_5892), 
      .ZN(n_8_0_5890));
   INV_X1 i_8_0_6129 (.A(n_8_0_5892), .ZN(n_8_0_5891));
   AOI21_X1 i_8_0_6130 (.A(\out_bs[6] [4]), .B1(n_8_0_6550), .B2(\out_bs[6] [3]), 
      .ZN(n_8_0_5892));
   NAND2_X1 i_8_0_6131 (.A1(n_8_0_7010), .A2(n_8_0_7009), .ZN(n_8_0_5893));
   NOR2_X1 i_8_0_6132 (.A1(\out_bs[6] [4]), .A2(\out_bs[6] [3]), .ZN(n_8_0_5894));
   OAI21_X1 i_8_0_6133 (.A(n_8_0_5896), .B1(n_8_0_6795), .B2(n_8_0_297), 
      .ZN(n_8_0_5895));
   OAI211_X1 i_8_0_6134 (.A(n_8_0_6636), .B(n_8_0_5897), .C1(n_8_0_6796), 
      .C2(n_8_0_6912), .ZN(n_8_0_5896));
   OR2_X1 i_8_0_6135 (.A1(\out_bs[4] [4]), .A2(n_8_0_6559), .ZN(n_8_0_5897));
   AOI21_X1 i_8_0_6136 (.A(n_8_0_5899), .B1(n_8_0_5900), .B2(n_8_0_6264), 
      .ZN(n_8_0_5898));
   NOR2_X1 i_8_0_6137 (.A1(n_8_0_6525), .A2(n_8_0_5901), .ZN(n_8_0_5899));
   AOI21_X1 i_8_0_6138 (.A(n_8_0_108), .B1(n_8_0_6782), .B2(n_8_0_5901), 
      .ZN(n_8_0_5900));
   AOI21_X1 i_8_0_6139 (.A(\out_bs[1] [4]), .B1(n_8_0_6531), .B2(\out_bs[1] [3]), 
      .ZN(n_8_0_5901));
   AOI21_X1 i_8_0_6140 (.A(n_8_0_5984), .B1(n_8_0_6532), .B2(n_8_0_7070), 
      .ZN(n_8_0_5902));
   AOI21_X1 i_8_0_6141 (.A(n_8_0_5904), .B1(n_8_0_6772), .B2(n_8_0_171), 
      .ZN(n_8_0_5903));
   AOI22_X1 i_8_0_6142 (.A1(n_8_0_6773), .A2(n_8_0_6947), .B1(n_8_0_5905), 
      .B2(n_8_0_6712), .ZN(n_8_0_5904));
   NOR2_X1 i_8_0_6143 (.A1(n_8_0_5991), .A2(n_8_0_5906), .ZN(n_8_0_5905));
   NOR3_X1 i_8_0_6144 (.A1(\out_bs[2] [4]), .A2(\out_bs[2] [1]), .A3(
      \out_bs[2] [0]), .ZN(n_8_0_5906));
   INV_X1 i_8_0_6145 (.A(n_8_0_5908), .ZN(n_8_0_5907));
   AOI21_X1 i_8_0_6146 (.A(\out_bs[0] [4]), .B1(n_8_0_6522), .B2(\out_bs[0] [3]), 
      .ZN(n_8_0_5908));
   OAI21_X1 i_8_0_6147 (.A(n_8_0_5910), .B1(n_8_0_5913), .B2(n_8_0_486), 
      .ZN(n_8_0_5909));
   NAND2_X1 i_8_0_6148 (.A1(n_8_0_6233), .A2(n_8_0_5911), .ZN(n_8_0_5910));
   NAND2_X1 i_8_0_6149 (.A1(n_8_0_5913), .A2(n_8_0_486), .ZN(n_8_0_5911));
   NOR2_X1 i_8_0_6150 (.A1(n_8_0_5913), .A2(n_8_0_486), .ZN(n_8_0_5912));
   NAND2_X1 i_8_0_6151 (.A1(n_8_0_5914), .A2(n_8_0_6728), .ZN(n_8_0_5913));
   OAI21_X1 i_8_0_6153 (.A(n_8_0_5916), .B1(n_8_0_6837), .B2(n_8_0_234), 
      .ZN(n_8_0_5915));
   OAI211_X1 i_8_0_6154 (.A(n_8_0_6659), .B(n_8_0_5917), .C1(n_8_0_6843), 
      .C2(n_8_0_6923), .ZN(n_8_0_5916));
   NOR2_X1 i_8_0_6155 (.A1(n_8_0_6008), .A2(n_8_0_5918), .ZN(n_8_0_5917));
   NOR2_X1 i_8_0_6156 (.A1(n_8_0_6565), .A2(\out_bs[3] [4]), .ZN(n_8_0_5918));
   AOI211_X1 i_8_0_6157 (.A(n_8_0_6376), .B(n_8_0_5920), .C1(n_8_0_360), 
      .C2(n_8_0_6511), .ZN(n_8_0_5919));
   NOR2_X1 i_8_0_6158 (.A1(n_8_0_5921), .A2(\out_bs[5] [4]), .ZN(n_8_0_5920));
   OAI21_X1 i_8_0_6159 (.A(n_8_0_6515), .B1(n_8_0_6824), .B2(n_8_0_360), 
      .ZN(n_8_0_5921));
   AOI21_X1 i_8_0_6160 (.A(n_8_0_6853), .B1(n_8_0_5923), .B2(n_8_0_5922), 
      .ZN(n_175));
   NOR4_X1 i_8_0_6161 (.A1(n_8_0_5945), .A2(n_8_0_5937), .A3(n_8_0_5933), 
      .A4(n_8_0_5925), .ZN(n_8_0_5922));
   AOI211_X1 i_8_0_6162 (.A(n_8_0_5949), .B(n_8_0_5924), .C1(n_8_0_6731), 
      .C2(n_8_0_5950), .ZN(n_8_0_5923));
   NAND3_X1 i_8_0_6163 (.A1(n_8_0_5955), .A2(n_8_0_5930), .A3(n_8_0_5958), 
      .ZN(n_8_0_5924));
   AOI221_X1 i_8_0_6164 (.A(n_8_0_5929), .B1(n_8_0_5927), .B2(n_8_0_6795), 
      .C1(n_8_0_5926), .C2(n_8_0_298), .ZN(n_8_0_5925));
   OAI21_X1 i_8_0_6165 (.A(n_8_0_6555), .B1(n_8_0_6640), .B2(\out_bs[4] [4]), 
      .ZN(n_8_0_5926));
   NOR2_X1 i_8_0_6166 (.A1(\out_bs[4] [4]), .A2(n_8_0_6640), .ZN(n_8_0_5927));
   NAND2_X1 i_8_0_6167 (.A1(n_8_0_6795), .A2(n_8_0_6635), .ZN(n_8_0_5928));
   NOR2_X1 i_8_0_6168 (.A1(n_8_0_6794), .A2(n_8_0_6636), .ZN(n_8_0_5929));
   AOI22_X1 i_8_0_6169 (.A1(n_8_0_6838), .A2(n_8_0_6922), .B1(n_8_0_5931), 
      .B2(n_8_0_6659), .ZN(n_8_0_5930));
   AOI21_X1 i_8_0_6170 (.A(n_8_0_5932), .B1(n_8_0_6844), .B2(n_8_0_235), 
      .ZN(n_8_0_5931));
   AOI21_X1 i_8_0_6171 (.A(\out_bs[3] [4]), .B1(\out_bs[3] [3]), .B2(n_8_0_6653), 
      .ZN(n_8_0_5932));
   OAI21_X1 i_8_0_6172 (.A(n_8_0_5934), .B1(n_8_0_6755), .B2(n_8_0_424), 
      .ZN(n_8_0_5933));
   OAI211_X1 i_8_0_6173 (.A(n_8_0_6753), .B(n_8_0_5935), .C1(n_8_0_6759), 
      .C2(n_8_0_6880), .ZN(n_8_0_5934));
   OAI21_X1 i_8_0_6174 (.A(n_8_0_7010), .B1(n_8_0_7009), .B2(n_8_0_6743), 
      .ZN(n_8_0_5935));
   AOI21_X1 i_8_0_6175 (.A(\out_bs[6] [4]), .B1(\out_bs[6] [3]), .B2(n_8_0_6744), 
      .ZN(n_8_0_5936));
   AOI21_X1 i_8_0_6176 (.A(n_8_0_5938), .B1(n_8_0_5939), .B2(n_8_0_46), .ZN(
      n_8_0_5937));
   AOI21_X1 i_8_0_6177 (.A(n_8_0_6810), .B1(n_8_0_6671), .B2(n_8_0_5940), 
      .ZN(n_8_0_5938));
   NAND2_X1 i_8_0_6178 (.A1(n_8_0_6248), .A2(n_8_0_5940), .ZN(n_8_0_5939));
   OAI21_X1 i_8_0_6179 (.A(n_8_0_7083), .B1(n_8_0_7082), .B2(n_8_0_6667), 
      .ZN(n_8_0_5940));
   AOI21_X1 i_8_0_6180 (.A(\out_bs[0] [4]), .B1(\out_bs[0] [3]), .B2(
      \out_bs[0] [2]), .ZN(n_8_0_5941));
   OAI21_X1 i_8_0_6181 (.A(n_8_0_7083), .B1(n_8_0_7082), .B2(n_8_0_7081), 
      .ZN(n_8_0_5942));
   NAND2_X1 i_8_0_6182 (.A1(n_8_0_7083), .A2(n_8_0_7082), .ZN(n_8_0_5943));
   NOR2_X1 i_8_0_6183 (.A1(\out_bs[0] [4]), .A2(\out_bs[0] [3]), .ZN(n_8_0_5944));
   AOI21_X1 i_8_0_6184 (.A(n_8_0_5946), .B1(n_8_0_6772), .B2(n_8_0_172), 
      .ZN(n_8_0_5945));
   AOI22_X1 i_8_0_6185 (.A1(n_8_0_6773), .A2(n_8_0_6946), .B1(n_8_0_5948), 
      .B2(n_8_0_6712), .ZN(n_8_0_5946));
   AOI21_X1 i_8_0_6186 (.A(\out_bs[2] [4]), .B1(\out_bs[2] [3]), .B2(n_8_0_6613), 
      .ZN(n_8_0_5947));
   OAI21_X1 i_8_0_6187 (.A(n_8_0_7058), .B1(n_8_0_7057), .B2(n_8_0_6612), 
      .ZN(n_8_0_5948));
   NOR2_X1 i_8_0_6188 (.A1(n_8_0_5951), .A2(n_8_0_487), .ZN(n_8_0_5949));
   NAND2_X1 i_8_0_6189 (.A1(n_8_0_5951), .A2(n_8_0_487), .ZN(n_8_0_5950));
   NAND2_X1 i_8_0_6190 (.A1(n_8_0_6728), .A2(n_8_0_5952), .ZN(n_8_0_5951));
   INV_X1 i_8_0_6192 (.A(n_8_0_5954), .ZN(n_8_0_5953));
   AOI21_X1 i_8_0_6194 (.A(n_8_0_5956), .B1(n_8_0_6825), .B2(n_8_0_6900), 
      .ZN(n_8_0_5955));
   AOI211_X1 i_8_0_6195 (.A(n_8_0_6685), .B(n_8_0_5957), .C1(n_8_0_6824), 
      .C2(n_8_0_361), .ZN(n_8_0_5956));
   NOR2_X1 i_8_0_6196 (.A1(\out_bs[5] [4]), .A2(n_8_0_6676), .ZN(n_8_0_5957));
   NAND2_X1 i_8_0_6197 (.A1(n_8_0_5959), .A2(n_8_0_5960), .ZN(n_8_0_5958));
   OAI21_X1 i_8_0_6198 (.A(n_8_0_6782), .B1(n_8_0_6693), .B2(n_8_0_5961), 
      .ZN(n_8_0_5959));
   OAI21_X1 i_8_0_6199 (.A(n_8_0_109), .B1(n_8_0_6525), .B2(n_8_0_5961), 
      .ZN(n_8_0_5960));
   OAI21_X1 i_8_0_6200 (.A(n_8_0_5983), .B1(n_8_0_6700), .B2(\out_bs[1] [4]), 
      .ZN(n_8_0_5961));
   OAI21_X1 i_8_0_6205 (.A(n_8_0_6511), .B1(n_8_0_6376), .B2(n_8_0_362), 
      .ZN(n_8_0_5965));
   OAI21_X1 i_8_0_6206 (.A(n_8_0_6673), .B1(n_8_0_6824), .B2(n_8_0_362), 
      .ZN(n_8_0_5966));
   AOI21_X1 i_8_0_6209 (.A(n_8_0_5970), .B1(n_8_0_6745), .B2(n_8_0_7010), 
      .ZN(n_8_0_5969));
   AOI21_X1 i_8_0_6210 (.A(\out_bs[6] [4]), .B1(\out_bs[6] [3]), .B2(
      \out_bs[6] [2]), .ZN(n_8_0_5970));
   AOI22_X1 i_8_0_6217 (.A1(n_8_0_5979), .A2(n_8_0_5978), .B1(n_8_0_6970), 
      .B2(n_8_0_6781), .ZN(n_8_0_5977));
   AOI21_X1 i_8_0_6218 (.A(n_8_0_6693), .B1(n_8_0_6784), .B2(n_8_0_110), 
      .ZN(n_8_0_5978));
   AOI21_X1 i_8_0_6219 (.A(n_8_0_5980), .B1(n_8_0_6690), .B2(n_8_0_7070), 
      .ZN(n_8_0_5979));
   AOI21_X1 i_8_0_6220 (.A(\out_bs[1] [4]), .B1(\out_bs[1] [3]), .B2(
      \out_bs[1] [2]), .ZN(n_8_0_5980));
   NOR2_X1 i_8_0_6221 (.A1(n_8_0_5984), .A2(n_8_0_5982), .ZN(n_8_0_5981));
   NOR2_X1 i_8_0_6222 (.A1(\out_bs[1] [4]), .A2(\out_bs[1] [2]), .ZN(n_8_0_5982));
   NAND2_X1 i_8_0_6223 (.A1(n_8_0_7070), .A2(n_8_0_7069), .ZN(n_8_0_5983));
   NOR2_X1 i_8_0_6224 (.A1(\out_bs[1] [4]), .A2(\out_bs[1] [3]), .ZN(n_8_0_5984));
   INV_X1 i_8_0_6226 (.A(n_8_0_5987), .ZN(n_8_0_5986));
   OAI22_X1 i_8_0_6227 (.A1(n_8_0_6772), .A2(n_8_0_173), .B1(n_8_0_5988), 
      .B2(n_8_0_6711), .ZN(n_8_0_5987));
   OAI21_X1 i_8_0_6228 (.A(n_8_0_5990), .B1(n_8_0_6710), .B2(\out_bs[2] [4]), 
      .ZN(n_8_0_5988));
   NOR2_X1 i_8_0_6229 (.A1(n_8_0_5992), .A2(n_8_0_5991), .ZN(n_8_0_5989));
   INV_X1 i_8_0_6230 (.A(n_8_0_5991), .ZN(n_8_0_5990));
   AOI21_X1 i_8_0_6231 (.A(\out_bs[2] [4]), .B1(\out_bs[2] [3]), .B2(
      \out_bs[2] [2]), .ZN(n_8_0_5991));
   NOR2_X1 i_8_0_6232 (.A1(\out_bs[2] [4]), .A2(n_8_0_6710), .ZN(n_8_0_5992));
   INV_X1 i_8_0_6234 (.A(n_8_0_5995), .ZN(n_8_0_5994));
   AOI211_X1 i_8_0_6235 (.A(n_8_0_5996), .B(n_8_0_6635), .C1(n_8_0_6795), 
      .C2(n_8_0_299), .ZN(n_8_0_5995));
   AOI21_X1 i_8_0_6236 (.A(\out_bs[4] [4]), .B1(\out_bs[4] [0]), .B2(n_8_0_6640), 
      .ZN(n_8_0_5996));
   OAI211_X1 i_8_0_6237 (.A(n_8_0_6594), .B(n_8_0_5998), .C1(n_8_0_5999), 
      .C2(n_8_0_6810), .ZN(n_8_0_5997));
   OAI21_X1 i_8_0_6238 (.A(n_8_0_47), .B1(n_8_0_6247), .B2(n_8_0_6000), .ZN(
      n_8_0_5998));
   OAI21_X1 i_8_0_6239 (.A(n_8_0_7083), .B1(n_8_0_7082), .B2(n_8_0_6665), 
      .ZN(n_8_0_5999));
   NOR2_X1 i_8_0_6240 (.A1(\out_bs[0] [4]), .A2(n_8_0_6664), .ZN(n_8_0_6000));
   INV_X1 i_8_0_6241 (.A(n_8_0_6002), .ZN(n_8_0_6001));
   OAI21_X1 i_8_0_6242 (.A(n_8_0_6004), .B1(n_8_0_6003), .B2(n_8_0_6838), 
      .ZN(n_8_0_6002));
   NOR2_X1 i_8_0_6243 (.A1(n_8_0_6006), .A2(n_8_0_6658), .ZN(n_8_0_6003));
   OAI21_X1 i_8_0_6244 (.A(n_8_0_236), .B1(n_8_0_6575), .B2(n_8_0_6006), 
      .ZN(n_8_0_6004));
   AOI21_X1 i_8_0_6245 (.A(n_8_0_6008), .B1(n_8_0_6649), .B2(n_8_0_7045), 
      .ZN(n_8_0_6005));
   OAI21_X1 i_8_0_6246 (.A(n_8_0_6007), .B1(n_8_0_6650), .B2(\out_bs[3] [4]), 
      .ZN(n_8_0_6006));
   NAND2_X1 i_8_0_6247 (.A1(n_8_0_7045), .A2(n_8_0_7044), .ZN(n_8_0_6007));
   NOR2_X1 i_8_0_6248 (.A1(\out_bs[3] [4]), .A2(\out_bs[3] [3]), .ZN(n_8_0_6008));
   AOI21_X1 i_8_0_6249 (.A(n_8_0_6853), .B1(n_8_0_6010), .B2(n_8_0_6009), 
      .ZN(n_176));
   NOR3_X1 i_8_0_6250 (.A1(n_8_0_6014), .A2(n_8_0_6013), .A3(n_8_0_6012), 
      .ZN(n_8_0_6009));
   NOR3_X1 i_8_0_6251 (.A1(n_8_0_6016), .A2(n_8_0_6015), .A3(n_8_0_6011), 
      .ZN(n_8_0_6010));
   AOI22_X1 i_8_0_6252 (.A1(n_8_0_6587), .A2(n_8_0_426), .B1(n_8_0_6747), 
      .B2(n_8_0_6755), .ZN(n_8_0_6011));
   OAI21_X1 i_8_0_6253 (.A(n_8_0_6305), .B1(n_8_0_6219), .B2(n_8_0_237), 
      .ZN(n_8_0_6012));
   AOI22_X1 i_8_0_6254 (.A1(n_8_0_6509), .A2(n_8_0_363), .B1(n_8_0_6824), 
      .B2(n_8_0_6683), .ZN(n_8_0_6013));
   AOI22_X1 i_8_0_6255 (.A1(n_8_0_300), .A2(n_8_0_6189), .B1(n_8_0_6795), 
      .B2(n_8_0_6634), .ZN(n_8_0_6014));
   AOI21_X1 i_8_0_6256 (.A(n_8_0_48), .B1(n_8_0_6811), .B2(n_8_0_6669), .ZN(
      n_8_0_6015));
   NAND3_X1 i_8_0_6257 (.A1(n_8_0_6018), .A2(n_8_0_6017), .A3(n_8_0_6022), 
      .ZN(n_8_0_6016));
   AOI221_X1 i_8_0_6258 (.A(n_8_0_6021), .B1(n_8_0_6248), .B2(\out_bs[0] [4]), 
      .C1(n_8_0_6731), .C2(n_8_0_6020), .ZN(n_8_0_6017));
   AOI21_X1 i_8_0_6259 (.A(n_8_0_6019), .B1(n_8_0_6605), .B2(\out_bs[2] [4]), 
      .ZN(n_8_0_6018));
   AOI21_X1 i_8_0_6260 (.A(n_8_0_174), .B1(n_8_0_6772), .B2(n_8_0_6702), 
      .ZN(n_8_0_6019));
   NAND2_X1 i_8_0_6261 (.A1(n_8_0_6715), .A2(n_8_0_489), .ZN(n_8_0_6020));
   NOR2_X1 i_8_0_6262 (.A1(n_8_0_6715), .A2(n_8_0_489), .ZN(n_8_0_6021));
   OAI21_X1 i_8_0_6263 (.A(n_8_0_6023), .B1(n_8_0_6781), .B2(n_8_0_6969), 
      .ZN(n_8_0_6022));
   OAI22_X1 i_8_0_6264 (.A1(n_8_0_111), .A2(n_8_0_6782), .B1(n_8_0_6693), 
      .B2(n_8_0_7070), .ZN(n_8_0_6023));
   AOI21_X1 i_8_0_6265 (.A(n_8_0_6853), .B1(n_8_0_6027), .B2(n_8_0_6024), 
      .ZN(n_177));
   NOR2_X1 i_8_0_6266 (.A1(n_8_0_6037), .A2(n_8_0_6025), .ZN(n_8_0_6024));
   OAI211_X1 i_8_0_6267 (.A(n_8_0_6026), .B(n_8_0_6047), .C1(n_8_0_6051), 
      .C2(n_8_0_49), .ZN(n_8_0_6025));
   AOI21_X1 i_8_0_6268 (.A(n_8_0_6055), .B1(n_8_0_6053), .B2(n_8_0_6248), 
      .ZN(n_8_0_6026));
   NOR4_X1 i_8_0_6269 (.A1(n_8_0_6043), .A2(n_8_0_6032), .A3(n_8_0_6028), 
      .A4(n_8_0_6061), .ZN(n_8_0_6027));
   INV_X1 i_8_0_6270 (.A(n_8_0_6029), .ZN(n_8_0_6028));
   AOI22_X1 i_8_0_6271 (.A1(n_8_0_6910), .A2(n_8_0_6794), .B1(n_8_0_6031), 
      .B2(n_8_0_6030), .ZN(n_8_0_6029));
   AOI21_X1 i_8_0_6272 (.A(n_8_0_6634), .B1(n_8_0_6797), .B2(n_8_0_301), 
      .ZN(n_8_0_6030));
   OR2_X1 i_8_0_6273 (.A1(n_8_0_6092), .A2(\out_bs[4] [0]), .ZN(n_8_0_6031));
   OAI21_X1 i_8_0_6274 (.A(n_8_0_6033), .B1(n_8_0_6755), .B2(n_8_0_427), 
      .ZN(n_8_0_6032));
   INV_X1 i_8_0_6275 (.A(n_8_0_6034), .ZN(n_8_0_6033));
   AOI211_X1 i_8_0_6276 (.A(n_8_0_6747), .B(n_8_0_6036), .C1(n_8_0_6758), 
      .C2(n_8_0_427), .ZN(n_8_0_6034));
   NOR2_X1 i_8_0_6277 (.A1(n_8_0_6036), .A2(n_8_0_7010), .ZN(n_8_0_6035));
   NOR2_X1 i_8_0_6278 (.A1(n_8_0_6088), .A2(\out_bs[6] [0]), .ZN(n_8_0_6036));
   AOI21_X1 i_8_0_6279 (.A(n_8_0_6038), .B1(n_8_0_6039), .B2(n_8_0_6232), 
      .ZN(n_8_0_6037));
   AND2_X1 i_8_0_6280 (.A1(n_8_0_6040), .A2(n_8_0_490), .ZN(n_8_0_6038));
   OR2_X1 i_8_0_6281 (.A1(n_8_0_6040), .A2(n_8_0_490), .ZN(n_8_0_6039));
   NAND3_X1 i_8_0_6282 (.A1(n_8_0_6042), .A2(n_8_0_6728), .A3(\out_bs[7] [4]), 
      .ZN(n_8_0_6040));
   AOI21_X1 i_8_0_6285 (.A(n_8_0_6044), .B1(n_8_0_6772), .B2(n_8_0_175), 
      .ZN(n_8_0_6043));
   INV_X1 i_8_0_6286 (.A(n_8_0_6045), .ZN(n_8_0_6044));
   OAI22_X1 i_8_0_6287 (.A1(n_8_0_175), .A2(n_8_0_6772), .B1(n_8_0_6711), 
      .B2(n_8_0_6046), .ZN(n_8_0_6045));
   AOI21_X1 i_8_0_6288 (.A(n_8_0_6709), .B1(n_8_0_6335), .B2(\out_bs[2] [4]), 
      .ZN(n_8_0_6046));
   OAI21_X1 i_8_0_6289 (.A(n_8_0_6048), .B1(n_8_0_6783), .B2(n_8_0_6968), 
      .ZN(n_8_0_6047));
   OAI22_X1 i_8_0_6290 (.A1(n_8_0_112), .A2(n_8_0_6782), .B1(n_8_0_6693), 
      .B2(n_8_0_6049), .ZN(n_8_0_6048));
   NAND2_X1 i_8_0_6291 (.A1(n_8_0_6050), .A2(\out_bs[1] [4]), .ZN(n_8_0_6049));
   NAND2_X1 i_8_0_6292 (.A1(n_8_0_6395), .A2(n_8_0_6269), .ZN(n_8_0_6050));
   AOI21_X1 i_8_0_6293 (.A(n_8_0_6810), .B1(n_8_0_6671), .B2(n_8_0_6053), 
      .ZN(n_8_0_6051));
   NAND2_X1 i_8_0_6294 (.A1(n_8_0_6053), .A2(\out_bs[0] [6]), .ZN(n_8_0_6052));
   AOI21_X1 i_8_0_6295 (.A(n_8_0_7083), .B1(n_8_0_6345), .B2(n_8_0_7082), 
      .ZN(n_8_0_6053));
   AOI21_X1 i_8_0_6297 (.A(n_8_0_6056), .B1(n_8_0_6058), .B2(n_8_0_364), 
      .ZN(n_8_0_6055));
   AOI21_X1 i_8_0_6298 (.A(n_8_0_6825), .B1(n_8_0_6684), .B2(n_8_0_6059), 
      .ZN(n_8_0_6056));
   NAND2_X1 i_8_0_6299 (.A1(n_8_0_6059), .A2(\out_bs[5] [4]), .ZN(n_8_0_6057));
   NAND2_X1 i_8_0_6300 (.A1(n_8_0_6510), .A2(n_8_0_6059), .ZN(n_8_0_6058));
   NAND2_X1 i_8_0_6301 (.A1(n_8_0_6518), .A2(n_8_0_6166), .ZN(n_8_0_6059));
   INV_X1 i_8_0_6302 (.A(n_8_0_6061), .ZN(n_8_0_6060));
   OAI211_X1 i_8_0_6303 (.A(n_8_0_6574), .B(n_8_0_6062), .C1(n_8_0_6564), 
      .C2(n_8_0_238), .ZN(n_8_0_6061));
   NAND3_X1 i_8_0_6304 (.A1(n_8_0_6063), .A2(n_8_0_6655), .A3(n_8_0_6357), 
      .ZN(n_8_0_6062));
   NAND2_X1 i_8_0_6305 (.A1(n_8_0_238), .A2(n_8_0_6842), .ZN(n_8_0_6063));
   AND2_X1 i_8_0_6306 (.A1(n_8_0_6064), .A2(n_8_0_6854), .ZN(n_178));
   NAND3_X1 i_8_0_6307 (.A1(n_8_0_6099), .A2(n_8_0_6076), .A3(n_8_0_6065), 
      .ZN(n_8_0_6064));
   NOR4_X1 i_8_0_6308 (.A1(n_8_0_6094), .A2(n_8_0_6071), .A3(n_8_0_6066), 
      .A4(n_8_0_6067), .ZN(n_8_0_6065));
   OAI211_X1 i_8_0_6309 (.A(n_8_0_6083), .B(n_8_0_6089), .C1(n_8_0_50), .C2(
      n_8_0_6081), .ZN(n_8_0_6066));
   OAI21_X1 i_8_0_6310 (.A(n_8_0_6068), .B1(n_8_0_6772), .B2(n_8_0_176), 
      .ZN(n_8_0_6067));
   NAND3_X1 i_8_0_6311 (.A1(n_8_0_6070), .A2(n_8_0_6069), .A3(n_8_0_6712), 
      .ZN(n_8_0_6068));
   AOI21_X1 i_8_0_6312 (.A(n_8_0_7058), .B1(n_8_0_6400), .B2(n_8_0_7057), 
      .ZN(n_8_0_6069));
   NAND2_X1 i_8_0_6313 (.A1(n_8_0_6772), .A2(n_8_0_176), .ZN(n_8_0_6070));
   INV_X1 i_8_0_6314 (.A(n_8_0_6072), .ZN(n_8_0_6071));
   AOI22_X1 i_8_0_6315 (.A1(n_8_0_6073), .A2(n_8_0_6074), .B1(n_8_0_6781), 
      .B2(n_8_0_6967), .ZN(n_8_0_6072));
   AOI21_X1 i_8_0_6316 (.A(n_8_0_6693), .B1(n_8_0_6784), .B2(n_8_0_113), 
      .ZN(n_8_0_6073));
   INV_X1 i_8_0_6317 (.A(n_8_0_6075), .ZN(n_8_0_6074));
   OAI21_X1 i_8_0_6318 (.A(\out_bs[1] [4]), .B1(n_8_0_6394), .B2(\out_bs[1] [3]), 
      .ZN(n_8_0_6075));
   AOI221_X1 i_8_0_6319 (.A(n_8_0_6077), .B1(n_8_0_6248), .B2(n_8_0_6082), 
      .C1(n_8_0_6233), .C2(n_8_0_6078), .ZN(n_8_0_6076));
   NOR2_X1 i_8_0_6320 (.A1(n_8_0_6079), .A2(n_8_0_491), .ZN(n_8_0_6077));
   NAND2_X1 i_8_0_6321 (.A1(n_8_0_6079), .A2(n_8_0_491), .ZN(n_8_0_6078));
   NAND3_X1 i_8_0_6322 (.A1(n_8_0_6080), .A2(n_8_0_6728), .A3(\out_bs[7] [4]), 
      .ZN(n_8_0_6079));
   AOI21_X1 i_8_0_6324 (.A(n_8_0_6810), .B1(n_8_0_6671), .B2(n_8_0_6082), 
      .ZN(n_8_0_6081));
   AOI21_X1 i_8_0_6325 (.A(n_8_0_7083), .B1(n_8_0_6421), .B2(n_8_0_7082), 
      .ZN(n_8_0_6082));
   OAI21_X1 i_8_0_6326 (.A(n_8_0_6084), .B1(n_8_0_6085), .B2(n_8_0_6754), 
      .ZN(n_8_0_6083));
   OAI21_X1 i_8_0_6327 (.A(n_8_0_428), .B1(n_8_0_6588), .B2(n_8_0_6086), 
      .ZN(n_8_0_6084));
   NOR2_X1 i_8_0_6328 (.A1(n_8_0_6752), .A2(n_8_0_6086), .ZN(n_8_0_6085));
   NAND2_X1 i_8_0_6329 (.A1(n_8_0_6088), .A2(\out_bs[6] [4]), .ZN(n_8_0_6086));
   AOI21_X1 i_8_0_6330 (.A(n_8_0_7010), .B1(n_8_0_6387), .B2(n_8_0_7009), 
      .ZN(n_8_0_6087));
   NAND2_X1 i_8_0_6331 (.A1(n_8_0_6387), .A2(n_8_0_7009), .ZN(n_8_0_6088));
   NAND2_X1 i_8_0_6332 (.A1(n_8_0_6091), .A2(n_8_0_6090), .ZN(n_8_0_6089));
   OAI21_X1 i_8_0_6333 (.A(n_8_0_6795), .B1(n_8_0_6634), .B2(n_8_0_6093), 
      .ZN(n_8_0_6090));
   OAI21_X1 i_8_0_6334 (.A(n_8_0_302), .B1(n_8_0_6189), .B2(n_8_0_6093), 
      .ZN(n_8_0_6091));
   OR2_X1 i_8_0_6335 (.A1(n_8_0_6170), .A2(\out_bs[4] [1]), .ZN(n_8_0_6092));
   NOR2_X1 i_8_0_6336 (.A1(n_8_0_6170), .A2(\out_bs[4] [1]), .ZN(n_8_0_6093));
   AOI21_X1 i_8_0_6337 (.A(n_8_0_6095), .B1(n_8_0_6096), .B2(n_8_0_365), 
      .ZN(n_8_0_6094));
   AOI21_X1 i_8_0_6338 (.A(n_8_0_6825), .B1(n_8_0_6684), .B2(n_8_0_6097), 
      .ZN(n_8_0_6095));
   NAND2_X1 i_8_0_6339 (.A1(n_8_0_6510), .A2(n_8_0_6097), .ZN(n_8_0_6096));
   NAND2_X1 i_8_0_6340 (.A1(n_8_0_6166), .A2(n_8_0_7019), .ZN(n_8_0_6097));
   NOR2_X1 i_8_0_6341 (.A1(n_8_0_6165), .A2(\out_bs[5] [1]), .ZN(n_8_0_6098));
   AOI21_X1 i_8_0_6342 (.A(n_8_0_6100), .B1(n_8_0_6101), .B2(n_8_0_6413), 
      .ZN(n_8_0_6099));
   OAI21_X1 i_8_0_6343 (.A(n_8_0_6574), .B1(n_8_0_6564), .B2(n_8_0_239), 
      .ZN(n_8_0_6100));
   AOI21_X1 i_8_0_6344 (.A(n_8_0_6654), .B1(n_8_0_6842), .B2(n_8_0_239), 
      .ZN(n_8_0_6101));
   NAND3_X1 i_8_0_6350 (.A1(n_8_0_6107), .A2(n_8_0_6655), .A3(n_8_0_6108), 
      .ZN(n_8_0_6106));
   NAND2_X1 i_8_0_6351 (.A1(n_8_0_240), .A2(n_8_0_6842), .ZN(n_8_0_6107));
   NAND2_X1 i_8_0_6352 (.A1(n_8_0_6161), .A2(n_8_0_6651), .ZN(n_8_0_6108));
   NOR2_X1 i_8_0_6353 (.A1(n_8_0_6428), .A2(\out_bs[3] [3]), .ZN(n_8_0_6109));
   OAI21_X1 i_8_0_6355 (.A(n_8_0_6795), .B1(n_8_0_6634), .B2(n_8_0_6114), 
      .ZN(n_8_0_6111));
   OAI21_X1 i_8_0_6356 (.A(n_8_0_303), .B1(n_8_0_6189), .B2(n_8_0_6114), 
      .ZN(n_8_0_6112));
   NAND2_X1 i_8_0_6357 (.A1(n_8_0_6171), .A2(n_8_0_6639), .ZN(n_8_0_6113));
   NOR2_X1 i_8_0_6358 (.A1(n_8_0_6435), .A2(\out_bs[4] [3]), .ZN(n_8_0_6114));
   AOI21_X1 i_8_0_6364 (.A(n_8_0_6122), .B1(n_8_0_6121), .B2(n_8_0_6753), 
      .ZN(n_8_0_6120));
   AOI21_X1 i_8_0_6365 (.A(n_8_0_6123), .B1(n_8_0_6755), .B2(n_8_0_429), 
      .ZN(n_8_0_6121));
   NOR2_X1 i_8_0_6366 (.A1(n_8_0_429), .A2(n_8_0_6755), .ZN(n_8_0_6122));
   AOI21_X1 i_8_0_6367 (.A(n_8_0_6751), .B1(n_8_0_6480), .B2(\out_bs[6] [4]), 
      .ZN(n_8_0_6123));
   OAI22_X1 i_8_0_6369 (.A1(n_8_0_114), .A2(n_8_0_6782), .B1(n_8_0_6693), 
      .B2(n_8_0_6126), .ZN(n_8_0_6125));
   OAI21_X1 i_8_0_6370 (.A(\out_bs[1] [4]), .B1(n_8_0_6447), .B2(\out_bs[1] [3]), 
      .ZN(n_8_0_6126));
   OAI21_X1 i_8_0_6371 (.A(n_8_0_6147), .B1(n_8_0_6690), .B2(n_8_0_7070), 
      .ZN(n_8_0_6127));
   INV_X1 i_8_0_6372 (.A(n_8_0_6129), .ZN(n_8_0_6128));
   AOI22_X1 i_8_0_6374 (.A1(n_8_0_6945), .A2(n_8_0_6773), .B1(n_8_0_6712), 
      .B2(n_8_0_6131), .ZN(n_8_0_6130));
   NAND2_X1 i_8_0_6375 (.A1(n_8_0_6705), .A2(n_8_0_6151), .ZN(n_8_0_6131));
   INV_X1 i_8_0_6376 (.A(n_8_0_6133), .ZN(n_8_0_6132));
   OAI22_X1 i_8_0_6377 (.A1(n_8_0_366), .A2(n_8_0_6134), .B1(n_8_0_6135), 
      .B2(n_8_0_6509), .ZN(n_8_0_6133));
   AOI21_X1 i_8_0_6378 (.A(n_8_0_6825), .B1(n_8_0_6684), .B2(n_8_0_6136), 
      .ZN(n_8_0_6134));
   INV_X1 i_8_0_6379 (.A(n_8_0_6136), .ZN(n_8_0_6135));
   NAND2_X1 i_8_0_6380 (.A1(n_8_0_6166), .A2(n_8_0_6677), .ZN(n_8_0_6136));
   AOI21_X1 i_8_0_6382 (.A(n_8_0_51), .B1(n_8_0_6811), .B2(n_8_0_6139), .ZN(
      n_8_0_6138));
   INV_X1 i_8_0_6383 (.A(n_8_0_6140), .ZN(n_8_0_6139));
   AOI21_X1 i_8_0_6384 (.A(n_8_0_7083), .B1(n_8_0_6442), .B2(n_8_0_7082), 
      .ZN(n_8_0_6140));
   AND2_X1 i_8_0_6385 (.A1(n_8_0_6141), .A2(n_8_0_6854), .ZN(n_179));
   NAND4_X1 i_8_0_6386 (.A1(n_8_0_6142), .A2(n_8_0_6148), .A3(n_8_0_6155), 
      .A4(n_8_0_6143), .ZN(n_8_0_6141));
   NOR4_X1 i_8_0_6387 (.A1(n_8_0_6167), .A2(n_8_0_6163), .A3(n_8_0_6158), 
      .A4(n_8_0_6144), .ZN(n_8_0_6142));
   AOI21_X1 i_8_0_6388 (.A(n_8_0_6152), .B1(n_8_0_6172), .B2(n_8_0_6173), 
      .ZN(n_8_0_6143));
   OAI21_X1 i_8_0_6389 (.A(n_8_0_6145), .B1(n_8_0_6147), .B2(n_8_0_6525), 
      .ZN(n_8_0_6144));
   NAND2_X1 i_8_0_6390 (.A1(n_8_0_6146), .A2(n_8_0_6264), .ZN(n_8_0_6145));
   AOI21_X1 i_8_0_6391 (.A(n_8_0_115), .B1(n_8_0_6782), .B2(n_8_0_6147), 
      .ZN(n_8_0_6146));
   OAI21_X1 i_8_0_6392 (.A(\out_bs[1] [4]), .B1(\out_bs[1] [3]), .B2(
      \out_bs[1] [2]), .ZN(n_8_0_6147));
   OAI21_X1 i_8_0_6393 (.A(n_8_0_6149), .B1(n_8_0_6773), .B2(n_8_0_6944), 
      .ZN(n_8_0_6148));
   OAI22_X1 i_8_0_6394 (.A1(n_8_0_178), .A2(n_8_0_6772), .B1(n_8_0_6711), 
      .B2(n_8_0_6151), .ZN(n_8_0_6149));
   AOI21_X1 i_8_0_6395 (.A(n_8_0_7058), .B1(n_8_0_7057), .B2(n_8_0_7056), 
      .ZN(n_8_0_6150));
   OAI21_X1 i_8_0_6396 (.A(\out_bs[2] [4]), .B1(\out_bs[2] [3]), .B2(
      \out_bs[2] [2]), .ZN(n_8_0_6151));
   AOI21_X1 i_8_0_6397 (.A(n_8_0_6153), .B1(n_8_0_6755), .B2(n_8_0_430), 
      .ZN(n_8_0_6152));
   INV_X1 i_8_0_6398 (.A(n_8_0_6154), .ZN(n_8_0_6153));
   OAI22_X1 i_8_0_6399 (.A1(n_8_0_430), .A2(n_8_0_6755), .B1(n_8_0_6752), 
      .B2(n_8_0_6293), .ZN(n_8_0_6154));
   OAI21_X1 i_8_0_6400 (.A(n_8_0_6156), .B1(n_8_0_6729), .B2(n_8_0_6869), 
      .ZN(n_8_0_6155));
   OAI22_X1 i_8_0_6401 (.A1(n_8_0_493), .A2(n_8_0_6730), .B1(n_8_0_6715), 
      .B2(n_8_0_6157), .ZN(n_8_0_6156));
   OAI21_X1 i_8_0_6403 (.A(n_8_0_6159), .B1(n_8_0_6837), .B2(n_8_0_241), 
      .ZN(n_8_0_6158));
   NAND3_X1 i_8_0_6404 (.A1(n_8_0_6162), .A2(n_8_0_6160), .A3(n_8_0_6655), 
      .ZN(n_8_0_6159));
   NAND2_X1 i_8_0_6405 (.A1(n_8_0_7044), .A2(n_8_0_7043), .ZN(n_8_0_6160));
   NOR2_X1 i_8_0_6406 (.A1(\out_bs[3] [3]), .A2(\out_bs[3] [2]), .ZN(n_8_0_6161));
   NAND2_X1 i_8_0_6407 (.A1(n_8_0_241), .A2(n_8_0_6842), .ZN(n_8_0_6162));
   OAI22_X1 i_8_0_6408 (.A1(n_8_0_367), .A2(n_8_0_6164), .B1(n_8_0_6166), 
      .B2(n_8_0_6509), .ZN(n_8_0_6163));
   AOI21_X1 i_8_0_6409 (.A(n_8_0_6825), .B1(n_8_0_6684), .B2(n_8_0_6165), 
      .ZN(n_8_0_6164));
   NAND2_X1 i_8_0_6410 (.A1(n_8_0_7021), .A2(n_8_0_7020), .ZN(n_8_0_6165));
   NOR2_X1 i_8_0_6411 (.A1(\out_bs[5] [3]), .A2(\out_bs[5] [2]), .ZN(n_8_0_6166));
   AOI21_X1 i_8_0_6412 (.A(n_8_0_6168), .B1(n_8_0_6795), .B2(n_8_0_304), 
      .ZN(n_8_0_6167));
   INV_X1 i_8_0_6413 (.A(n_8_0_6169), .ZN(n_8_0_6168));
   OAI22_X1 i_8_0_6414 (.A1(n_8_0_304), .A2(n_8_0_6795), .B1(n_8_0_6634), 
      .B2(n_8_0_6171), .ZN(n_8_0_6169));
   NAND2_X1 i_8_0_6415 (.A1(n_8_0_7032), .A2(n_8_0_7031), .ZN(n_8_0_6170));
   NOR2_X1 i_8_0_6416 (.A1(\out_bs[4] [3]), .A2(\out_bs[4] [2]), .ZN(n_8_0_6171));
   OAI21_X1 i_8_0_6417 (.A(n_8_0_52), .B1(n_8_0_6247), .B2(n_8_0_6174), .ZN(
      n_8_0_6172));
   OAI21_X1 i_8_0_6418 (.A(n_8_0_6811), .B1(n_8_0_6670), .B2(n_8_0_6174), 
      .ZN(n_8_0_6173));
   NAND2_X1 i_8_0_6419 (.A1(n_8_0_6175), .A2(\out_bs[0] [4]), .ZN(n_8_0_6174));
   NAND2_X1 i_8_0_6420 (.A1(n_8_0_7082), .A2(n_8_0_7081), .ZN(n_8_0_6175));
   OAI22_X1 i_8_0_6426 (.A1(n_8_0_179), .A2(n_8_0_6772), .B1(n_8_0_6711), 
      .B2(n_8_0_6182), .ZN(n_8_0_6180));
   INV_X1 i_8_0_6427 (.A(n_8_0_6182), .ZN(n_8_0_6181));
   AOI21_X1 i_8_0_6428 (.A(n_8_0_6709), .B1(n_8_0_6536), .B2(\out_bs[2] [4]), 
      .ZN(n_8_0_6182));
   AOI21_X1 i_8_0_6429 (.A(n_8_0_53), .B1(n_8_0_6811), .B2(n_8_0_6184), .ZN(
      n_8_0_6183));
   NAND2_X1 i_8_0_6430 (.A1(n_8_0_6185), .A2(n_8_0_6671), .ZN(n_8_0_6184));
   AOI21_X1 i_8_0_6431 (.A(n_8_0_7083), .B1(n_8_0_6523), .B2(n_8_0_7082), 
      .ZN(n_8_0_6185));
   OAI21_X1 i_8_0_6433 (.A(n_8_0_6795), .B1(n_8_0_6634), .B2(n_8_0_6192), 
      .ZN(n_8_0_6187));
   OAI21_X1 i_8_0_6434 (.A(n_8_0_305), .B1(n_8_0_6554), .B2(n_8_0_6190), 
      .ZN(n_8_0_6188));
   NAND2_X1 i_8_0_6435 (.A1(n_8_0_6637), .A2(n_8_0_6557), .ZN(n_8_0_6189));
   NAND2_X1 i_8_0_6436 (.A1(n_8_0_6191), .A2(\out_bs[4] [4]), .ZN(n_8_0_6190));
   NAND2_X1 i_8_0_6437 (.A1(n_8_0_6245), .A2(n_8_0_6630), .ZN(n_8_0_6191));
   NOR2_X1 i_8_0_6438 (.A1(n_8_0_6560), .A2(\out_bs[4] [3]), .ZN(n_8_0_6192));
   INV_X1 i_8_0_6440 (.A(n_8_0_6195), .ZN(n_8_0_6194));
   AOI211_X1 i_8_0_6441 (.A(n_8_0_6752), .B(n_8_0_6196), .C1(n_8_0_6758), 
      .C2(n_8_0_431), .ZN(n_8_0_6195));
   OAI21_X1 i_8_0_6442 (.A(\out_bs[6] [4]), .B1(n_8_0_6550), .B2(\out_bs[6] [3]), 
      .ZN(n_8_0_6196));
   NOR2_X1 i_8_0_6443 (.A1(n_8_0_6198), .A2(n_8_0_7010), .ZN(n_8_0_6197));
   NOR2_X1 i_8_0_6444 (.A1(n_8_0_6550), .A2(\out_bs[6] [3]), .ZN(n_8_0_6198));
   OAI21_X1 i_8_0_6450 (.A(n_8_0_6782), .B1(n_8_0_6693), .B2(n_8_0_6206), 
      .ZN(n_8_0_6204));
   OAI21_X1 i_8_0_6451 (.A(n_8_0_116), .B1(n_8_0_6525), .B2(n_8_0_6206), 
      .ZN(n_8_0_6205));
   OAI21_X1 i_8_0_6452 (.A(\out_bs[1] [4]), .B1(n_8_0_6531), .B2(\out_bs[1] [3]), 
      .ZN(n_8_0_6206));
   NAND3_X1 i_8_0_6454 (.A1(n_8_0_6209), .A2(n_8_0_6684), .A3(n_8_0_6210), 
      .ZN(n_8_0_6208));
   NAND2_X1 i_8_0_6455 (.A1(n_8_0_6619), .A2(n_8_0_368), .ZN(n_8_0_6209));
   OAI21_X1 i_8_0_6456 (.A(n_8_0_7021), .B1(n_8_0_6518), .B2(n_8_0_7020), 
      .ZN(n_8_0_6210));
   NOR2_X1 i_8_0_6457 (.A1(\out_bs[5] [3]), .A2(n_8_0_6517), .ZN(n_8_0_6211));
   OAI21_X1 i_8_0_6459 (.A(n_8_0_6837), .B1(n_8_0_6654), .B2(n_8_0_6216), 
      .ZN(n_8_0_6213));
   OAI21_X1 i_8_0_6460 (.A(n_8_0_242), .B1(n_8_0_6305), .B2(n_8_0_6216), 
      .ZN(n_8_0_6214));
   NAND2_X1 i_8_0_6461 (.A1(n_8_0_6566), .A2(n_8_0_7044), .ZN(n_8_0_6215));
   NOR2_X1 i_8_0_6462 (.A1(n_8_0_6565), .A2(\out_bs[3] [3]), .ZN(n_8_0_6216));
   NAND2_X1 i_8_0_6463 (.A1(n_8_0_7044), .A2(n_8_0_6652), .ZN(n_8_0_6217));
   NOR2_X1 i_8_0_6464 (.A1(\out_bs[3] [3]), .A2(n_8_0_6653), .ZN(n_8_0_6218));
   NOR2_X1 i_8_0_6465 (.A1(n_8_0_6838), .A2(n_8_0_6655), .ZN(n_8_0_6219));
   NOR2_X1 i_8_0_6466 (.A1(n_8_0_6220), .A2(n_8_0_6853), .ZN(n_180));
   NOR4_X1 i_8_0_6467 (.A1(n_8_0_6246), .A2(n_8_0_6221), .A3(n_8_0_6241), 
      .A4(n_8_0_6254), .ZN(n_8_0_6220));
   NAND4_X1 i_8_0_6468 (.A1(n_8_0_6231), .A2(n_8_0_6222), .A3(n_8_0_6229), 
      .A4(n_8_0_6239), .ZN(n_8_0_6221));
   NOR2_X1 i_8_0_6469 (.A1(n_8_0_6227), .A2(n_8_0_6223), .ZN(n_8_0_6222));
   OAI22_X1 i_8_0_6470 (.A1(n_8_0_432), .A2(n_8_0_6224), .B1(n_8_0_6226), 
      .B2(n_8_0_6588), .ZN(n_8_0_6223));
   AOI21_X1 i_8_0_6471 (.A(n_8_0_6754), .B1(n_8_0_6753), .B2(n_8_0_6225), 
      .ZN(n_8_0_6224));
   OAI21_X1 i_8_0_6472 (.A(n_8_0_6750), .B1(n_8_0_6743), .B2(n_8_0_7010), 
      .ZN(n_8_0_6225));
   AOI21_X1 i_8_0_6473 (.A(n_8_0_6751), .B1(n_8_0_6744), .B2(\out_bs[6] [4]), 
      .ZN(n_8_0_6226));
   OAI22_X1 i_8_0_6474 (.A1(n_8_0_369), .A2(n_8_0_6228), .B1(n_8_0_6301), 
      .B2(n_8_0_6509), .ZN(n_8_0_6227));
   AOI21_X1 i_8_0_6475 (.A(n_8_0_6825), .B1(n_8_0_6684), .B2(n_8_0_6300), 
      .ZN(n_8_0_6228));
   OAI21_X1 i_8_0_6476 (.A(n_8_0_6230), .B1(n_8_0_6773), .B2(n_8_0_6942), 
      .ZN(n_8_0_6229));
   OAI22_X1 i_8_0_6477 (.A1(n_8_0_180), .A2(n_8_0_6772), .B1(n_8_0_6711), 
      .B2(n_8_0_6287), .ZN(n_8_0_6230));
   AOI21_X1 i_8_0_6478 (.A(n_8_0_6235), .B1(n_8_0_6233), .B2(n_8_0_6234), 
      .ZN(n_8_0_6231));
   OAI21_X1 i_8_0_6481 (.A(n_8_0_495), .B1(n_8_0_6236), .B2(n_8_0_6999), 
      .ZN(n_8_0_6234));
   NOR3_X1 i_8_0_6482 (.A1(n_8_0_6999), .A2(n_8_0_6236), .A3(n_8_0_495), 
      .ZN(n_8_0_6235));
   NAND2_X1 i_8_0_6483 (.A1(n_8_0_6237), .A2(n_8_0_6717), .ZN(n_8_0_6236));
   OAI21_X1 i_8_0_6486 (.A(n_8_0_6240), .B1(n_8_0_6783), .B2(n_8_0_6965), 
      .ZN(n_8_0_6239));
   OAI22_X1 i_8_0_6487 (.A1(n_8_0_117), .A2(n_8_0_6782), .B1(n_8_0_6693), 
      .B2(n_8_0_6270), .ZN(n_8_0_6240));
   OAI22_X1 i_8_0_6488 (.A1(n_8_0_306), .A2(n_8_0_6795), .B1(n_8_0_6245), 
      .B2(n_8_0_6242), .ZN(n_8_0_6241));
   INV_X1 i_8_0_6489 (.A(n_8_0_6243), .ZN(n_8_0_6242));
   AOI21_X1 i_8_0_6490 (.A(n_8_0_6634), .B1(n_8_0_6797), .B2(n_8_0_306), 
      .ZN(n_8_0_6243));
   NAND2_X1 i_8_0_6491 (.A1(n_8_0_7032), .A2(n_8_0_6642), .ZN(n_8_0_6244));
   NOR2_X1 i_8_0_6492 (.A1(\out_bs[4] [3]), .A2(n_8_0_6643), .ZN(n_8_0_6245));
   AOI211_X1 i_8_0_6493 (.A(n_8_0_6595), .B(n_8_0_6251), .C1(n_8_0_6247), 
      .C2(n_8_0_54), .ZN(n_8_0_6246));
   NOR2_X1 i_8_0_6495 (.A1(n_8_0_6812), .A2(n_8_0_6670), .ZN(n_8_0_6248));
   NOR2_X1 i_8_0_6497 (.A1(n_8_0_7085), .A2(n_8_0_6812), .ZN(n_8_0_6250));
   AOI21_X1 i_8_0_6498 (.A(n_8_0_6253), .B1(n_8_0_6810), .B2(n_8_0_6980), 
      .ZN(n_8_0_6251));
   INV_X1 i_8_0_6499 (.A(n_8_0_6253), .ZN(n_8_0_6252));
   OAI21_X1 i_8_0_6500 (.A(n_8_0_6662), .B1(n_8_0_6667), .B2(n_8_0_7083), 
      .ZN(n_8_0_6253));
   OAI211_X1 i_8_0_6501 (.A(n_8_0_6574), .B(n_8_0_6255), .C1(n_8_0_6564), 
      .C2(n_8_0_243), .ZN(n_8_0_6254));
   NAND3_X1 i_8_0_6502 (.A1(n_8_0_6256), .A2(n_8_0_6653), .A3(n_8_0_6655), 
      .ZN(n_8_0_6255));
   NAND2_X1 i_8_0_6503 (.A1(n_8_0_243), .A2(n_8_0_6842), .ZN(n_8_0_6256));
   AOI21_X1 i_8_0_6509 (.A(n_8_0_6663), .B1(n_8_0_6262), .B2(n_8_0_6668), 
      .ZN(n_8_0_6261));
   NOR2_X1 i_8_0_6510 (.A1(n_8_0_7083), .A2(n_8_0_7079), .ZN(n_8_0_6262));
   OAI211_X1 i_8_0_6511 (.A(n_8_0_6266), .B(n_8_0_6264), .C1(n_8_0_6781), 
      .C2(n_8_0_6268), .ZN(n_8_0_6263));
   NAND2_X1 i_8_0_6512 (.A1(n_8_0_6782), .A2(n_8_0_6693), .ZN(n_8_0_6264));
   NOR2_X1 i_8_0_6513 (.A1(n_8_0_6781), .A2(n_8_0_6694), .ZN(n_8_0_6265));
   NAND2_X1 i_8_0_6514 (.A1(n_8_0_6267), .A2(n_8_0_118), .ZN(n_8_0_6266));
   NAND3_X1 i_8_0_6515 (.A1(n_8_0_6783), .A2(n_8_0_6694), .A3(n_8_0_6268), 
      .ZN(n_8_0_6267));
   NOR2_X1 i_8_0_6516 (.A1(n_8_0_6270), .A2(n_8_0_6269), .ZN(n_8_0_6268));
   NOR2_X1 i_8_0_6517 (.A1(\out_bs[1] [3]), .A2(\out_bs[1] [0]), .ZN(n_8_0_6269));
   OAI21_X1 i_8_0_6518 (.A(\out_bs[1] [4]), .B1(\out_bs[1] [3]), .B2(n_8_0_6700), 
      .ZN(n_8_0_6270));
   OAI21_X1 i_8_0_6519 (.A(n_8_0_6695), .B1(n_8_0_6699), .B2(n_8_0_7070), 
      .ZN(n_8_0_6271));
   AOI21_X1 i_8_0_6521 (.A(n_8_0_6274), .B1(n_8_0_6797), .B2(n_8_0_307), 
      .ZN(n_8_0_6273));
   INV_X1 i_8_0_6522 (.A(n_8_0_6275), .ZN(n_8_0_6274));
   OAI21_X1 i_8_0_6523 (.A(n_8_0_6632), .B1(n_8_0_6629), .B2(n_8_0_7033), 
      .ZN(n_8_0_6275));
   OAI21_X1 i_8_0_6529 (.A(n_8_0_181), .B1(n_8_0_6604), .B2(n_8_0_6286), 
      .ZN(n_8_0_6281));
   NAND2_X1 i_8_0_6530 (.A1(\out_bs[2] [5]), .A2(n_8_0_6773), .ZN(n_8_0_6282));
   NOR2_X1 i_8_0_6531 (.A1(n_8_0_7059), .A2(n_8_0_6772), .ZN(n_8_0_6283));
   OAI21_X1 i_8_0_6532 (.A(n_8_0_6772), .B1(n_8_0_6711), .B2(n_8_0_6286), 
      .ZN(n_8_0_6284));
   INV_X1 i_8_0_6533 (.A(n_8_0_6286), .ZN(n_8_0_6285));
   OAI21_X1 i_8_0_6534 (.A(n_8_0_6288), .B1(n_8_0_6709), .B2(\out_bs[2] [0]), 
      .ZN(n_8_0_6286));
   INV_X1 i_8_0_6535 (.A(n_8_0_6288), .ZN(n_8_0_6287));
   OAI21_X1 i_8_0_6536 (.A(n_8_0_6708), .B1(n_8_0_6612), .B2(n_8_0_7058), 
      .ZN(n_8_0_6288));
   AOI21_X1 i_8_0_6538 (.A(n_8_0_6292), .B1(n_8_0_6758), .B2(n_8_0_433), 
      .ZN(n_8_0_6290));
   AOI21_X1 i_8_0_6539 (.A(n_8_0_6293), .B1(n_8_0_6745), .B2(n_8_0_6750), 
      .ZN(n_8_0_6291));
   OAI211_X1 i_8_0_6540 (.A(\out_bs[6] [4]), .B(n_8_0_6294), .C1(n_8_0_6746), 
      .C2(\out_bs[6] [3]), .ZN(n_8_0_6292));
   NAND2_X1 i_8_0_6541 (.A1(n_8_0_6294), .A2(\out_bs[6] [4]), .ZN(n_8_0_6293));
   NAND2_X1 i_8_0_6542 (.A1(n_8_0_7009), .A2(n_8_0_7008), .ZN(n_8_0_6294));
   INV_X1 i_8_0_6543 (.A(n_8_0_6296), .ZN(n_8_0_6295));
   AOI21_X1 i_8_0_6545 (.A(n_8_0_6825), .B1(n_8_0_6684), .B2(n_8_0_6299), 
      .ZN(n_8_0_6297));
   AOI21_X1 i_8_0_6546 (.A(\out_bs[5] [3]), .B1(\out_bs[5] [0]), .B2(n_8_0_6682), 
      .ZN(n_8_0_6298));
   OAI21_X1 i_8_0_6547 (.A(n_8_0_7021), .B1(n_8_0_7020), .B2(n_8_0_6677), 
      .ZN(n_8_0_6299));
   NAND2_X1 i_8_0_6548 (.A1(n_8_0_7021), .A2(n_8_0_6681), .ZN(n_8_0_6300));
   NOR2_X1 i_8_0_6549 (.A1(\out_bs[5] [3]), .A2(n_8_0_6682), .ZN(n_8_0_6301));
   OAI21_X1 i_8_0_6551 (.A(n_8_0_6564), .B1(n_8_0_6649), .B2(n_8_0_6654), 
      .ZN(n_8_0_6303));
   OAI21_X1 i_8_0_6552 (.A(n_8_0_244), .B1(n_8_0_6649), .B2(n_8_0_6305), 
      .ZN(n_8_0_6304));
   NAND2_X1 i_8_0_6553 (.A1(n_8_0_6841), .A2(n_8_0_6655), .ZN(n_8_0_6305));
   AOI21_X1 i_8_0_6554 (.A(n_8_0_6853), .B1(n_8_0_6323), .B2(n_8_0_6306), 
      .ZN(n_181));
   NOR4_X1 i_8_0_6555 (.A1(n_8_0_6314), .A2(n_8_0_6311), .A3(n_8_0_6310), 
      .A4(n_8_0_6307), .ZN(n_8_0_6306));
   AOI21_X1 i_8_0_6556 (.A(n_8_0_6432), .B1(n_8_0_6308), .B2(n_8_0_308), 
      .ZN(n_8_0_6307));
   NAND2_X1 i_8_0_6557 (.A1(n_8_0_6794), .A2(n_8_0_6624), .ZN(n_8_0_6308));
   INV_X1 i_8_0_6558 (.A(n_8_0_6310), .ZN(n_8_0_6309));
   AOI21_X1 i_8_0_6559 (.A(n_8_0_6584), .B1(n_8_0_6586), .B2(n_8_0_434), 
      .ZN(n_8_0_6310));
   OAI21_X1 i_8_0_6560 (.A(n_8_0_6312), .B1(n_8_0_6417), .B2(n_8_0_56), .ZN(
      n_8_0_6311));
   OAI21_X1 i_8_0_6561 (.A(n_8_0_6313), .B1(n_8_0_6825), .B2(n_8_0_6897), 
      .ZN(n_8_0_6312));
   OAI22_X1 i_8_0_6562 (.A1(n_8_0_6824), .A2(n_8_0_371), .B1(n_8_0_7021), 
      .B2(n_8_0_6683), .ZN(n_8_0_6313));
   NAND4_X1 i_8_0_6563 (.A1(n_8_0_6318), .A2(n_8_0_6599), .A3(n_8_0_6320), 
      .A4(n_8_0_6315), .ZN(n_8_0_6314));
   OAI21_X1 i_8_0_6564 (.A(n_8_0_6316), .B1(n_8_0_6317), .B2(n_8_0_6731), 
      .ZN(n_8_0_6315));
   NAND2_X1 i_8_0_6565 (.A1(n_8_0_6714), .A2(n_8_0_497), .ZN(n_8_0_6316));
   NOR2_X1 i_8_0_6566 (.A1(n_8_0_6714), .A2(n_8_0_497), .ZN(n_8_0_6317));
   OAI21_X1 i_8_0_6567 (.A(n_8_0_6319), .B1(n_8_0_6608), .B2(n_8_0_6773), 
      .ZN(n_8_0_6318));
   OAI21_X1 i_8_0_6568 (.A(n_8_0_182), .B1(n_8_0_6708), .B2(n_8_0_6604), 
      .ZN(n_8_0_6319));
   AOI21_X1 i_8_0_6569 (.A(n_8_0_6322), .B1(n_8_0_6691), .B2(n_8_0_6781), 
      .ZN(n_8_0_6320));
   NAND2_X1 i_8_0_6570 (.A1(n_8_0_6781), .A2(\out_bs[1] [5]), .ZN(n_8_0_6321));
   AOI21_X1 i_8_0_6571 (.A(n_8_0_119), .B1(n_8_0_6782), .B2(n_8_0_6692), 
      .ZN(n_8_0_6322));
   NAND2_X1 i_8_0_6572 (.A1(n_8_0_6563), .A2(n_8_0_6324), .ZN(n_8_0_6323));
   OAI21_X1 i_8_0_6573 (.A(n_8_0_245), .B1(n_8_0_6837), .B2(n_8_0_6645), 
      .ZN(n_8_0_6324));
   NAND2_X1 i_8_0_6574 (.A1(\out_bs[3] [5]), .A2(n_8_0_6838), .ZN(n_8_0_6325));
   NOR2_X1 i_8_0_6575 (.A1(n_8_0_7046), .A2(n_8_0_6837), .ZN(n_8_0_6326));
   NOR2_X1 i_8_0_6576 (.A1(n_8_0_6327), .A2(n_8_0_6853), .ZN(n_182));
   NOR3_X1 i_8_0_6577 (.A1(n_8_0_6358), .A2(n_8_0_6330), .A3(n_8_0_6328), 
      .ZN(n_8_0_6327));
   OR4_X1 i_8_0_6578 (.A1(n_8_0_6346), .A2(n_8_0_6337), .A3(n_8_0_6331), 
      .A4(n_8_0_6329), .ZN(n_8_0_6328));
   OAI21_X1 i_8_0_6579 (.A(n_8_0_6353), .B1(n_8_0_6811), .B2(n_8_0_57), .ZN(
      n_8_0_6329));
   AOI211_X1 i_8_0_6580 (.A(n_8_0_6345), .B(n_8_0_6660), .C1(n_8_0_6811), 
      .C2(n_8_0_57), .ZN(n_8_0_6330));
   AOI21_X1 i_8_0_6581 (.A(n_8_0_6332), .B1(n_8_0_6772), .B2(n_8_0_183), 
      .ZN(n_8_0_6331));
   AOI22_X1 i_8_0_6582 (.A1(n_8_0_6773), .A2(n_8_0_6941), .B1(n_8_0_6334), 
      .B2(n_8_0_6712), .ZN(n_8_0_6332));
   NAND2_X1 i_8_0_6583 (.A1(n_8_0_6335), .A2(n_8_0_6709), .ZN(n_8_0_6333));
   NOR2_X1 i_8_0_6584 (.A1(n_8_0_6336), .A2(n_8_0_6708), .ZN(n_8_0_6334));
   NAND2_X1 i_8_0_6585 (.A1(n_8_0_6400), .A2(n_8_0_7054), .ZN(n_8_0_6335));
   NOR2_X1 i_8_0_6586 (.A1(n_8_0_6399), .A2(\out_bs[2] [0]), .ZN(n_8_0_6336));
   OAI22_X1 i_8_0_6587 (.A1(n_8_0_120), .A2(n_8_0_6338), .B1(n_8_0_6339), 
      .B2(n_8_0_6525), .ZN(n_8_0_6337));
   AOI21_X1 i_8_0_6588 (.A(n_8_0_6781), .B1(n_8_0_6694), .B2(n_8_0_6340), 
      .ZN(n_8_0_6338));
   NAND2_X1 i_8_0_6589 (.A1(\out_bs[1] [4]), .A2(n_8_0_6341), .ZN(n_8_0_6339));
   NOR2_X1 i_8_0_6590 (.A1(n_8_0_6342), .A2(n_8_0_6695), .ZN(n_8_0_6340));
   NOR2_X1 i_8_0_6591 (.A1(n_8_0_6342), .A2(n_8_0_7069), .ZN(n_8_0_6341));
   NOR2_X1 i_8_0_6592 (.A1(n_8_0_6394), .A2(\out_bs[1] [0]), .ZN(n_8_0_6342));
   NOR2_X1 i_8_0_6593 (.A1(n_8_0_6345), .A2(n_8_0_6662), .ZN(n_8_0_6343));
   NAND2_X1 i_8_0_6594 (.A1(n_8_0_6421), .A2(n_8_0_7079), .ZN(n_8_0_6344));
   NOR2_X1 i_8_0_6595 (.A1(n_8_0_6420), .A2(\out_bs[0] [0]), .ZN(n_8_0_6345));
   OAI22_X1 i_8_0_6596 (.A1(n_8_0_309), .A2(n_8_0_6347), .B1(n_8_0_6348), 
      .B2(n_8_0_6554), .ZN(n_8_0_6346));
   AOI21_X1 i_8_0_6597 (.A(n_8_0_6794), .B1(n_8_0_6624), .B2(n_8_0_6352), 
      .ZN(n_8_0_6347));
   NAND2_X1 i_8_0_6598 (.A1(n_8_0_6352), .A2(n_8_0_6633), .ZN(n_8_0_6348));
   NOR2_X1 i_8_0_6599 (.A1(n_8_0_7033), .A2(n_8_0_6350), .ZN(n_8_0_6349));
   INV_X1 i_8_0_6600 (.A(n_8_0_6351), .ZN(n_8_0_6350));
   AND2_X1 i_8_0_6601 (.A1(n_8_0_6352), .A2(\out_bs[4] [3]), .ZN(n_8_0_6351));
   OR2_X1 i_8_0_6602 (.A1(n_8_0_6382), .A2(\out_bs[4] [0]), .ZN(n_8_0_6352));
   OAI211_X1 i_8_0_6603 (.A(n_8_0_6563), .B(n_8_0_6354), .C1(n_8_0_6357), 
      .C2(n_8_0_6838), .ZN(n_8_0_6353));
   OAI21_X1 i_8_0_6604 (.A(n_8_0_246), .B1(n_8_0_6575), .B2(n_8_0_6355), 
      .ZN(n_8_0_6354));
   NAND2_X1 i_8_0_6605 (.A1(n_8_0_6357), .A2(n_8_0_6648), .ZN(n_8_0_6355));
   AOI21_X1 i_8_0_6606 (.A(n_8_0_6647), .B1(n_8_0_6414), .B2(n_8_0_7041), 
      .ZN(n_8_0_6356));
   NAND2_X1 i_8_0_6607 (.A1(n_8_0_6414), .A2(n_8_0_7041), .ZN(n_8_0_6357));
   NAND3_X1 i_8_0_6608 (.A1(n_8_0_6370), .A2(n_8_0_6364), .A3(n_8_0_6359), 
      .ZN(n_8_0_6358));
   OAI21_X1 i_8_0_6609 (.A(n_8_0_6360), .B1(n_8_0_6729), .B2(n_8_0_6867), 
      .ZN(n_8_0_6359));
   OAI22_X1 i_8_0_6610 (.A1(n_8_0_498), .A2(n_8_0_6730), .B1(n_8_0_6715), 
      .B2(n_8_0_6361), .ZN(n_8_0_6360));
   NAND2_X1 i_8_0_6613 (.A1(n_8_0_6544), .A2(n_8_0_6996), .ZN(n_8_0_6363));
   OAI211_X1 i_8_0_6614 (.A(n_8_0_6583), .B(n_8_0_6365), .C1(n_8_0_6369), 
      .C2(n_8_0_6754), .ZN(n_8_0_6364));
   OAI21_X1 i_8_0_6615 (.A(n_8_0_435), .B1(n_8_0_6588), .B2(n_8_0_6366), 
      .ZN(n_8_0_6365));
   NAND2_X1 i_8_0_6616 (.A1(n_8_0_6369), .A2(n_8_0_6751), .ZN(n_8_0_6366));
   AOI21_X1 i_8_0_6617 (.A(n_8_0_6750), .B1(n_8_0_6387), .B2(n_8_0_7006), 
      .ZN(n_8_0_6367));
   AOI21_X1 i_8_0_6618 (.A(n_8_0_7009), .B1(n_8_0_6387), .B2(n_8_0_7006), 
      .ZN(n_8_0_6368));
   NAND2_X1 i_8_0_6619 (.A1(n_8_0_6387), .A2(n_8_0_7006), .ZN(n_8_0_6369));
   OAI211_X1 i_8_0_6620 (.A(n_8_0_6375), .B(n_8_0_6371), .C1(n_8_0_6373), 
      .C2(n_8_0_6825), .ZN(n_8_0_6370));
   OAI21_X1 i_8_0_6621 (.A(n_8_0_372), .B1(n_8_0_6511), .B2(n_8_0_6372), 
      .ZN(n_8_0_6371));
   NAND2_X1 i_8_0_6622 (.A1(n_8_0_6374), .A2(\out_bs[5] [4]), .ZN(n_8_0_6372));
   AOI21_X1 i_8_0_6623 (.A(n_8_0_7022), .B1(n_8_0_6680), .B2(n_8_0_6408), 
      .ZN(n_8_0_6373));
   NAND2_X1 i_8_0_6624 (.A1(n_8_0_6680), .A2(n_8_0_6408), .ZN(n_8_0_6374));
   NAND2_X1 i_8_0_6625 (.A1(n_8_0_6824), .A2(n_8_0_6685), .ZN(n_8_0_6375));
   AND2_X1 i_8_0_6626 (.A1(n_8_0_6824), .A2(n_8_0_6685), .ZN(n_8_0_6376));
   AOI22_X1 i_8_0_6630 (.A1(n_8_0_6908), .A2(n_8_0_6794), .B1(n_8_0_6636), 
      .B2(n_8_0_6380), .ZN(n_8_0_6379));
   AND2_X1 i_8_0_6631 (.A1(n_8_0_6382), .A2(n_8_0_6633), .ZN(n_8_0_6380));
   AND2_X1 i_8_0_6632 (.A1(n_8_0_6382), .A2(\out_bs[4] [3]), .ZN(n_8_0_6381));
   OR2_X1 i_8_0_6633 (.A1(\out_bs[4] [2]), .A2(\out_bs[4] [1]), .ZN(n_8_0_6382));
   NAND2_X1 i_8_0_6635 (.A1(n_8_0_6589), .A2(n_8_0_6385), .ZN(n_8_0_6384));
   NOR2_X1 i_8_0_6636 (.A1(n_8_0_6387), .A2(n_8_0_6750), .ZN(n_8_0_6385));
   NAND2_X1 i_8_0_6637 (.A1(n_8_0_7008), .A2(n_8_0_7007), .ZN(n_8_0_6386));
   NOR2_X1 i_8_0_6638 (.A1(\out_bs[6] [2]), .A2(\out_bs[6] [1]), .ZN(n_8_0_6387));
   NOR2_X1 i_8_0_6641 (.A1(n_8_0_121), .A2(n_8_0_6782), .ZN(n_8_0_6390));
   AOI21_X1 i_8_0_6642 (.A(n_8_0_6395), .B1(n_8_0_6782), .B2(n_8_0_121), 
      .ZN(n_8_0_6391));
   NAND2_X1 i_8_0_6643 (.A1(n_8_0_6696), .A2(n_8_0_6394), .ZN(n_8_0_6392));
   NOR2_X1 i_8_0_6644 (.A1(n_8_0_6395), .A2(n_8_0_6695), .ZN(n_8_0_6393));
   NAND2_X1 i_8_0_6645 (.A1(n_8_0_7068), .A2(n_8_0_7067), .ZN(n_8_0_6394));
   NOR2_X1 i_8_0_6646 (.A1(\out_bs[1] [2]), .A2(\out_bs[1] [1]), .ZN(n_8_0_6395));
   OAI22_X1 i_8_0_6648 (.A1(n_8_0_184), .A2(n_8_0_6772), .B1(n_8_0_6609), 
      .B2(n_8_0_6400), .ZN(n_8_0_6397));
   NOR2_X1 i_8_0_6649 (.A1(n_8_0_6400), .A2(n_8_0_6708), .ZN(n_8_0_6398));
   NAND2_X1 i_8_0_6650 (.A1(n_8_0_7056), .A2(n_8_0_7055), .ZN(n_8_0_6399));
   NOR2_X1 i_8_0_6651 (.A1(\out_bs[2] [2]), .A2(\out_bs[2] [1]), .ZN(n_8_0_6400));
   NOR2_X1 i_8_0_6656 (.A1(\out_bs[7] [2]), .A2(\out_bs[7] [1]), .ZN(n_8_0_6405));
   OAI22_X1 i_8_0_6658 (.A1(n_8_0_6824), .A2(n_8_0_373), .B1(n_8_0_6408), 
      .B2(n_8_0_6683), .ZN(n_8_0_6407));
   OAI21_X1 i_8_0_6659 (.A(\out_bs[5] [3]), .B1(\out_bs[5] [2]), .B2(
      \out_bs[5] [1]), .ZN(n_8_0_6408));
   AOI21_X1 i_8_0_6660 (.A(n_8_0_7021), .B1(n_8_0_7020), .B2(n_8_0_7019), 
      .ZN(n_8_0_6409));
   AOI22_X1 i_8_0_6662 (.A1(n_8_0_6838), .A2(n_8_0_6921), .B1(n_8_0_6412), 
      .B2(n_8_0_6659), .ZN(n_8_0_6411));
   NOR2_X1 i_8_0_6663 (.A1(n_8_0_6414), .A2(n_8_0_6647), .ZN(n_8_0_6412));
   NAND2_X1 i_8_0_6664 (.A1(n_8_0_7043), .A2(n_8_0_7042), .ZN(n_8_0_6413));
   NOR2_X1 i_8_0_6665 (.A1(\out_bs[3] [2]), .A2(\out_bs[3] [1]), .ZN(n_8_0_6414));
   OAI21_X1 i_8_0_6667 (.A(n_8_0_6811), .B1(n_8_0_6660), .B2(n_8_0_6421), 
      .ZN(n_8_0_6416));
   NOR2_X1 i_8_0_6668 (.A1(n_8_0_6810), .A2(n_8_0_6661), .ZN(n_8_0_6417));
   OAI21_X1 i_8_0_6669 (.A(n_8_0_58), .B1(n_8_0_6599), .B2(n_8_0_6421), .ZN(
      n_8_0_6418));
   NOR3_X1 i_8_0_6670 (.A1(n_8_0_6662), .A2(n_8_0_6596), .A3(n_8_0_6421), 
      .ZN(n_8_0_6419));
   NAND2_X1 i_8_0_6671 (.A1(n_8_0_7081), .A2(n_8_0_7080), .ZN(n_8_0_6420));
   NOR2_X1 i_8_0_6672 (.A1(\out_bs[0] [2]), .A2(\out_bs[0] [1]), .ZN(n_8_0_6421));
   AOI21_X1 i_8_0_6673 (.A(n_8_0_6853), .B1(n_8_0_6422), .B2(n_8_0_6463), 
      .ZN(n_183));
   AND4_X1 i_8_0_6674 (.A1(n_8_0_6423), .A2(n_8_0_6436), .A3(n_8_0_6449), 
      .A4(n_8_0_6476), .ZN(n_8_0_6422));
   AOI211_X1 i_8_0_6675 (.A(n_8_0_6443), .B(n_8_0_6424), .C1(n_8_0_6458), 
      .C2(n_8_0_6455), .ZN(n_8_0_6423));
   NAND2_X1 i_8_0_6676 (.A1(n_8_0_6430), .A2(n_8_0_6425), .ZN(n_8_0_6424));
   AOI21_X1 i_8_0_6677 (.A(n_8_0_6426), .B1(n_8_0_6838), .B2(n_8_0_6920), 
      .ZN(n_8_0_6425));
   AOI211_X1 i_8_0_6678 (.A(n_8_0_6645), .B(n_8_0_6429), .C1(n_8_0_6844), 
      .C2(n_8_0_248), .ZN(n_8_0_6426));
   NOR2_X1 i_8_0_6679 (.A1(n_8_0_6429), .A2(n_8_0_7044), .ZN(n_8_0_6427));
   NAND2_X1 i_8_0_6680 (.A1(n_8_0_7043), .A2(n_8_0_6651), .ZN(n_8_0_6428));
   AOI21_X1 i_8_0_6681 (.A(\out_bs[3] [2]), .B1(\out_bs[3] [1]), .B2(
      \out_bs[3] [0]), .ZN(n_8_0_6429));
   OAI21_X1 i_8_0_6682 (.A(n_8_0_6431), .B1(n_8_0_6435), .B2(n_8_0_6794), 
      .ZN(n_8_0_6430));
   OAI22_X1 i_8_0_6683 (.A1(n_8_0_311), .A2(n_8_0_6432), .B1(n_8_0_6433), 
      .B2(n_8_0_6554), .ZN(n_8_0_6431));
   NOR2_X1 i_8_0_6684 (.A1(n_8_0_6794), .A2(n_8_0_6624), .ZN(n_8_0_6432));
   NAND2_X1 i_8_0_6685 (.A1(n_8_0_6435), .A2(n_8_0_6633), .ZN(n_8_0_6433));
   AOI21_X1 i_8_0_6686 (.A(n_8_0_7032), .B1(n_8_0_7031), .B2(n_8_0_6639), 
      .ZN(n_8_0_6434));
   NAND2_X1 i_8_0_6687 (.A1(n_8_0_7031), .A2(n_8_0_6639), .ZN(n_8_0_6435));
   OAI211_X1 i_8_0_6688 (.A(n_8_0_6594), .B(n_8_0_6440), .C1(n_8_0_6439), 
      .C2(n_8_0_6810), .ZN(n_8_0_6436));
   NAND2_X1 i_8_0_6689 (.A1(\out_bs[0] [6]), .A2(n_8_0_6663), .ZN(n_8_0_6437));
   NOR2_X1 i_8_0_6690 (.A1(n_8_0_7085), .A2(n_8_0_6662), .ZN(n_8_0_6438));
   NOR2_X1 i_8_0_6691 (.A1(n_8_0_6442), .A2(n_8_0_6662), .ZN(n_8_0_6439));
   OAI21_X1 i_8_0_6692 (.A(n_8_0_59), .B1(n_8_0_6599), .B2(n_8_0_6442), .ZN(
      n_8_0_6440));
   INV_X1 i_8_0_6693 (.A(n_8_0_6442), .ZN(n_8_0_6441));
   AOI21_X1 i_8_0_6694 (.A(\out_bs[0] [2]), .B1(\out_bs[0] [1]), .B2(
      \out_bs[0] [0]), .ZN(n_8_0_6442));
   OAI21_X1 i_8_0_6695 (.A(n_8_0_6444), .B1(n_8_0_6782), .B2(n_8_0_122), 
      .ZN(n_8_0_6443));
   INV_X1 i_8_0_6696 (.A(n_8_0_6445), .ZN(n_8_0_6444));
   AOI211_X1 i_8_0_6697 (.A(n_8_0_6692), .B(n_8_0_6448), .C1(n_8_0_6784), 
      .C2(n_8_0_122), .ZN(n_8_0_6445));
   NOR2_X1 i_8_0_6698 (.A1(n_8_0_6448), .A2(n_8_0_6695), .ZN(n_8_0_6446));
   NAND2_X1 i_8_0_6699 (.A1(n_8_0_7068), .A2(n_8_0_6690), .ZN(n_8_0_6447));
   AOI21_X1 i_8_0_6700 (.A(\out_bs[1] [2]), .B1(\out_bs[1] [1]), .B2(
      \out_bs[1] [0]), .ZN(n_8_0_6448));
   OAI21_X1 i_8_0_6701 (.A(n_8_0_6450), .B1(n_8_0_6773), .B2(n_8_0_6939), 
      .ZN(n_8_0_6449));
   OAI22_X1 i_8_0_6702 (.A1(n_8_0_6772), .A2(n_8_0_185), .B1(n_8_0_6452), 
      .B2(n_8_0_6702), .ZN(n_8_0_6450));
   NOR2_X1 i_8_0_6703 (.A1(n_8_0_6453), .A2(n_8_0_6708), .ZN(n_8_0_6451));
   OAI21_X1 i_8_0_6704 (.A(\out_bs[2] [3]), .B1(\out_bs[2] [2]), .B2(n_8_0_6710), 
      .ZN(n_8_0_6452));
   NOR2_X1 i_8_0_6705 (.A1(\out_bs[2] [2]), .A2(n_8_0_6710), .ZN(n_8_0_6453));
   NAND2_X1 i_8_0_6706 (.A1(n_8_0_6458), .A2(n_8_0_6455), .ZN(n_8_0_6454));
   INV_X1 i_8_0_6707 (.A(n_8_0_6456), .ZN(n_8_0_6455));
   NOR2_X1 i_8_0_6708 (.A1(n_8_0_6825), .A2(n_8_0_6457), .ZN(n_8_0_6456));
   NOR3_X1 i_8_0_6709 (.A1(n_8_0_6459), .A2(n_8_0_374), .A3(n_8_0_6683), 
      .ZN(n_8_0_6457));
   OAI21_X1 i_8_0_6710 (.A(n_8_0_374), .B1(n_8_0_6683), .B2(n_8_0_6459), 
      .ZN(n_8_0_6458));
   NAND2_X1 i_8_0_6711 (.A1(n_8_0_6461), .A2(\out_bs[5] [3]), .ZN(n_8_0_6459));
   AOI21_X1 i_8_0_6712 (.A(n_8_0_7021), .B1(n_8_0_7020), .B2(n_8_0_6677), 
      .ZN(n_8_0_6460));
   NAND2_X1 i_8_0_6713 (.A1(n_8_0_7020), .A2(n_8_0_6677), .ZN(n_8_0_6461));
   INV_X1 i_8_0_6714 (.A(n_8_0_6463), .ZN(n_8_0_6462));
   OAI21_X1 i_8_0_6715 (.A(n_8_0_6472), .B1(n_8_0_6729), .B2(n_8_0_6865), 
      .ZN(n_8_0_6463));
   NAND2_X1 i_8_0_6716 (.A1(n_8_0_6729), .A2(n_8_0_6728), .ZN(n_8_0_6464));
   OAI22_X1 i_8_0_6724 (.A1(n_8_0_500), .A2(n_8_0_6730), .B1(n_8_0_6727), 
      .B2(n_8_0_6473), .ZN(n_8_0_6472));
   NAND2_X1 i_8_0_6725 (.A1(\out_bs[7] [4]), .A2(n_8_0_6474), .ZN(n_8_0_6473));
   AND2_X1 i_8_0_6726 (.A1(n_8_0_6475), .A2(\out_bs[7] [3]), .ZN(n_8_0_6474));
   OR2_X1 i_8_0_6727 (.A1(\out_bs[7] [2]), .A2(n_8_0_6726), .ZN(n_8_0_6475));
   OAI211_X1 i_8_0_6728 (.A(n_8_0_6583), .B(n_8_0_6477), .C1(n_8_0_6480), 
      .C2(n_8_0_6754), .ZN(n_8_0_6476));
   OAI21_X1 i_8_0_6729 (.A(n_8_0_437), .B1(n_8_0_6588), .B2(n_8_0_6478), 
      .ZN(n_8_0_6477));
   NAND2_X1 i_8_0_6730 (.A1(n_8_0_6480), .A2(n_8_0_6751), .ZN(n_8_0_6478));
   NOR2_X1 i_8_0_6731 (.A1(n_8_0_6481), .A2(n_8_0_6750), .ZN(n_8_0_6479));
   NAND2_X1 i_8_0_6732 (.A1(n_8_0_7008), .A2(n_8_0_6745), .ZN(n_8_0_6480));
   NOR2_X1 i_8_0_6733 (.A1(\out_bs[6] [2]), .A2(n_8_0_6746), .ZN(n_8_0_6481));
   AOI21_X1 i_8_0_6734 (.A(n_8_0_6853), .B1(n_8_0_6490), .B2(n_8_0_6482), 
      .ZN(n_184));
   AND3_X1 i_8_0_6735 (.A1(n_8_0_6488), .A2(n_8_0_6486), .A3(n_8_0_6483), 
      .ZN(n_8_0_6482));
   AOI21_X1 i_8_0_6736 (.A(n_8_0_6485), .B1(n_8_0_6484), .B2(\out_bs[1] [2]), 
      .ZN(n_8_0_6483));
   AOI21_X1 i_8_0_6737 (.A(n_8_0_6692), .B1(n_8_0_6782), .B2(n_8_0_123), 
      .ZN(n_8_0_6484));
   NOR2_X1 i_8_0_6738 (.A1(n_8_0_123), .A2(n_8_0_6782), .ZN(n_8_0_6485));
   OAI21_X1 i_8_0_6739 (.A(n_8_0_6487), .B1(n_8_0_6810), .B2(n_8_0_6978), 
      .ZN(n_8_0_6486));
   OAI22_X1 i_8_0_6740 (.A1(n_8_0_60), .A2(n_8_0_6811), .B1(n_8_0_6660), 
      .B2(n_8_0_7081), .ZN(n_8_0_6487));
   OAI21_X1 i_8_0_6741 (.A(n_8_0_6489), .B1(n_8_0_6729), .B2(n_8_0_6863), 
      .ZN(n_8_0_6488));
   OAI22_X1 i_8_0_6742 (.A1(n_8_0_501), .A2(n_8_0_6730), .B1(n_8_0_6714), 
      .B2(n_8_0_6996), .ZN(n_8_0_6489));
   AND4_X1 i_8_0_6743 (.A1(n_8_0_6497), .A2(n_8_0_6492), .A3(n_8_0_6491), 
      .A4(n_8_0_6495), .ZN(n_8_0_6490));
   AOI21_X1 i_8_0_6744 (.A(n_8_0_6501), .B1(n_8_0_6500), .B2(n_8_0_6499), 
      .ZN(n_8_0_6491));
   NAND2_X1 i_8_0_6745 (.A1(n_8_0_6494), .A2(n_8_0_6493), .ZN(n_8_0_6492));
   OAI21_X1 i_8_0_6746 (.A(n_8_0_6824), .B1(n_8_0_6683), .B2(n_8_0_6678), 
      .ZN(n_8_0_6493));
   OAI21_X1 i_8_0_6747 (.A(n_8_0_375), .B1(n_8_0_6678), .B2(n_8_0_6509), 
      .ZN(n_8_0_6494));
   OAI21_X1 i_8_0_6748 (.A(n_8_0_6496), .B1(n_8_0_6838), .B2(n_8_0_6919), 
      .ZN(n_8_0_6495));
   OAI22_X1 i_8_0_6749 (.A1(n_8_0_6837), .A2(n_8_0_249), .B1(n_8_0_7043), 
      .B2(n_8_0_6645), .ZN(n_8_0_6496));
   AOI21_X1 i_8_0_6750 (.A(n_8_0_6498), .B1(n_8_0_6794), .B2(n_8_0_6906), 
      .ZN(n_8_0_6497));
   AOI211_X1 i_8_0_6751 (.A(n_8_0_6641), .B(n_8_0_6634), .C1(n_8_0_6797), 
      .C2(n_8_0_312), .ZN(n_8_0_6498));
   NAND2_X1 i_8_0_6752 (.A1(n_8_0_6772), .A2(n_8_0_186), .ZN(n_8_0_6499));
   OAI22_X1 i_8_0_6753 (.A1(n_8_0_6772), .A2(n_8_0_186), .B1(n_8_0_6706), 
      .B2(n_8_0_6711), .ZN(n_8_0_6500));
   OAI21_X1 i_8_0_6754 (.A(n_8_0_6502), .B1(n_8_0_6755), .B2(n_8_0_438), 
      .ZN(n_8_0_6501));
   OAI211_X1 i_8_0_6755 (.A(n_8_0_6753), .B(n_8_0_6749), .C1(n_8_0_6759), 
      .C2(n_8_0_6876), .ZN(n_8_0_6502));
   NOR2_X1 i_8_0_6756 (.A1(n_8_0_6503), .A2(n_8_0_6853), .ZN(n_185));
   NOR3_X1 i_8_0_6757 (.A1(n_8_0_6504), .A2(n_8_0_6545), .A3(n_8_0_6552), 
      .ZN(n_8_0_6503));
   NAND4_X1 i_8_0_6758 (.A1(n_8_0_6505), .A2(n_8_0_6519), .A3(n_8_0_6533), 
      .A4(n_8_0_6538), .ZN(n_8_0_6504));
   NOR3_X1 i_8_0_6759 (.A1(n_8_0_6561), .A2(n_8_0_6524), .A3(n_8_0_6506), 
      .ZN(n_8_0_6505));
   AOI21_X1 i_8_0_6760 (.A(n_8_0_6507), .B1(n_8_0_6508), .B2(n_8_0_376), 
      .ZN(n_8_0_6506));
   AOI21_X1 i_8_0_6761 (.A(n_8_0_6825), .B1(n_8_0_6684), .B2(n_8_0_6516), 
      .ZN(n_8_0_6507));
   NAND2_X1 i_8_0_6762 (.A1(n_8_0_6516), .A2(n_8_0_6510), .ZN(n_8_0_6508));
   NAND2_X1 i_8_0_6763 (.A1(\out_bs[5] [4]), .A2(n_8_0_6512), .ZN(n_8_0_6509));
   NOR2_X1 i_8_0_6764 (.A1(n_8_0_6683), .A2(n_8_0_6619), .ZN(n_8_0_6510));
   NAND2_X1 i_8_0_6765 (.A1(\out_bs[5] [5]), .A2(n_8_0_6514), .ZN(n_8_0_6511));
   NOR2_X1 i_8_0_6766 (.A1(n_8_0_6685), .A2(n_8_0_6619), .ZN(n_8_0_6512));
   NAND2_X1 i_8_0_6767 (.A1(\out_bs[5] [6]), .A2(n_8_0_6825), .ZN(n_8_0_6513));
   NOR2_X1 i_8_0_6768 (.A1(n_8_0_7024), .A2(n_8_0_6619), .ZN(n_8_0_6514));
   NAND2_X1 i_8_0_6769 (.A1(\out_bs[5] [3]), .A2(n_8_0_6517), .ZN(n_8_0_6515));
   NOR2_X1 i_8_0_6770 (.A1(n_8_0_6518), .A2(n_8_0_6678), .ZN(n_8_0_6516));
   NOR2_X1 i_8_0_6771 (.A1(n_8_0_6518), .A2(n_8_0_7020), .ZN(n_8_0_6517));
   NOR2_X1 i_8_0_6772 (.A1(\out_bs[5] [1]), .A2(\out_bs[5] [0]), .ZN(n_8_0_6518));
   OAI211_X1 i_8_0_6773 (.A(n_8_0_6594), .B(n_8_0_6521), .C1(n_8_0_6520), 
      .C2(n_8_0_6810), .ZN(n_8_0_6519));
   OAI21_X1 i_8_0_6775 (.A(n_8_0_61), .B1(n_8_0_6599), .B2(n_8_0_6523), .ZN(
      n_8_0_6521));
   AOI21_X1 i_8_0_6776 (.A(n_8_0_7081), .B1(n_8_0_7080), .B2(n_8_0_7079), 
      .ZN(n_8_0_6522));
   OAI21_X1 i_8_0_6777 (.A(\out_bs[0] [2]), .B1(\out_bs[0] [1]), .B2(
      \out_bs[0] [0]), .ZN(n_8_0_6523));
   OAI21_X1 i_8_0_6778 (.A(n_8_0_6528), .B1(n_8_0_6782), .B2(n_8_0_124), 
      .ZN(n_8_0_6524));
   NAND2_X1 i_8_0_6779 (.A1(n_8_0_6783), .A2(n_8_0_6694), .ZN(n_8_0_6525));
   NAND2_X1 i_8_0_6780 (.A1(\out_bs[1] [6]), .A2(n_8_0_6783), .ZN(n_8_0_6526));
   NOR2_X1 i_8_0_6781 (.A1(n_8_0_7072), .A2(n_8_0_6784), .ZN(n_8_0_6527));
   INV_X1 i_8_0_6782 (.A(n_8_0_6529), .ZN(n_8_0_6528));
   AOI211_X1 i_8_0_6783 (.A(n_8_0_6693), .B(n_8_0_6530), .C1(n_8_0_6784), 
      .C2(n_8_0_124), .ZN(n_8_0_6529));
   NAND2_X1 i_8_0_6784 (.A1(n_8_0_6531), .A2(n_8_0_6696), .ZN(n_8_0_6530));
   NAND2_X1 i_8_0_6785 (.A1(n_8_0_6699), .A2(n_8_0_6698), .ZN(n_8_0_6531));
   OAI21_X1 i_8_0_6786 (.A(\out_bs[1] [2]), .B1(\out_bs[1] [1]), .B2(
      \out_bs[1] [0]), .ZN(n_8_0_6532));
   OAI21_X1 i_8_0_6787 (.A(n_8_0_6534), .B1(n_8_0_6773), .B2(n_8_0_6938), 
      .ZN(n_8_0_6533));
   OAI22_X1 i_8_0_6788 (.A1(n_8_0_187), .A2(n_8_0_6772), .B1(n_8_0_6609), 
      .B2(n_8_0_6537), .ZN(n_8_0_6534));
   NOR2_X1 i_8_0_6789 (.A1(n_8_0_6537), .A2(n_8_0_6708), .ZN(n_8_0_6535));
   INV_X1 i_8_0_6790 (.A(n_8_0_6537), .ZN(n_8_0_6536));
   OAI21_X1 i_8_0_6791 (.A(\out_bs[2] [2]), .B1(\out_bs[2] [1]), .B2(
      \out_bs[2] [0]), .ZN(n_8_0_6537));
   OAI21_X1 i_8_0_6792 (.A(n_8_0_6539), .B1(n_8_0_6729), .B2(n_8_0_6862), 
      .ZN(n_8_0_6538));
   OAI22_X1 i_8_0_6793 (.A1(n_8_0_502), .A2(n_8_0_6730), .B1(n_8_0_6715), 
      .B2(n_8_0_6540), .ZN(n_8_0_6539));
   NOR2_X1 i_8_0_6796 (.A1(n_8_0_6544), .A2(n_8_0_6996), .ZN(n_8_0_6542));
   NAND2_X1 i_8_0_6797 (.A1(\out_bs[7] [3]), .A2(n_8_0_6717), .ZN(n_8_0_6543));
   NOR2_X1 i_8_0_6798 (.A1(\out_bs[7] [1]), .A2(\out_bs[7] [0]), .ZN(n_8_0_6544));
   INV_X1 i_8_0_6799 (.A(n_8_0_6546), .ZN(n_8_0_6545));
   OAI211_X1 i_8_0_6800 (.A(n_8_0_6583), .B(n_8_0_6547), .C1(n_8_0_6550), 
      .C2(n_8_0_6754), .ZN(n_8_0_6546));
   OAI21_X1 i_8_0_6801 (.A(n_8_0_439), .B1(n_8_0_6588), .B2(n_8_0_6548), 
      .ZN(n_8_0_6547));
   NAND2_X1 i_8_0_6802 (.A1(n_8_0_6550), .A2(n_8_0_6751), .ZN(n_8_0_6548));
   NOR2_X1 i_8_0_6803 (.A1(n_8_0_6551), .A2(n_8_0_6750), .ZN(n_8_0_6549));
   AOI21_X1 i_8_0_6804 (.A(n_8_0_7008), .B1(n_8_0_7007), .B2(n_8_0_7006), 
      .ZN(n_8_0_6550));
   OAI21_X1 i_8_0_6805 (.A(\out_bs[6] [2]), .B1(\out_bs[6] [1]), .B2(
      \out_bs[6] [0]), .ZN(n_8_0_6551));
   OAI21_X1 i_8_0_6806 (.A(n_8_0_6553), .B1(n_8_0_6795), .B2(n_8_0_313), 
      .ZN(n_8_0_6552));
   OAI211_X1 i_8_0_6807 (.A(n_8_0_6636), .B(n_8_0_6558), .C1(n_8_0_6796), 
      .C2(n_8_0_6905), .ZN(n_8_0_6553));
   NAND2_X1 i_8_0_6808 (.A1(n_8_0_6796), .A2(n_8_0_6636), .ZN(n_8_0_6554));
   NOR2_X1 i_8_0_6809 (.A1(n_8_0_6797), .A2(n_8_0_6635), .ZN(n_8_0_6555));
   NAND2_X1 i_8_0_6810 (.A1(\out_bs[4] [6]), .A2(n_8_0_6796), .ZN(n_8_0_6556));
   NOR2_X1 i_8_0_6811 (.A1(n_8_0_7035), .A2(n_8_0_6797), .ZN(n_8_0_6557));
   AOI21_X1 i_8_0_6812 (.A(n_8_0_6632), .B1(n_8_0_6630), .B2(n_8_0_6642), 
      .ZN(n_8_0_6558));
   AOI21_X1 i_8_0_6813 (.A(n_8_0_7032), .B1(n_8_0_6642), .B2(n_8_0_6630), 
      .ZN(n_8_0_6559));
   NAND2_X1 i_8_0_6814 (.A1(n_8_0_6642), .A2(n_8_0_6630), .ZN(n_8_0_6560));
   OAI22_X1 i_8_0_6815 (.A1(n_8_0_250), .A2(n_8_0_6562), .B1(n_8_0_6566), 
      .B2(n_8_0_6574), .ZN(n_8_0_6561));
   AOI21_X1 i_8_0_6816 (.A(n_8_0_6838), .B1(n_8_0_6646), .B2(n_8_0_6565), 
      .ZN(n_8_0_6562));
   INV_X1 i_8_0_6817 (.A(n_8_0_6564), .ZN(n_8_0_6563));
   NOR2_X1 i_8_0_6818 (.A1(n_8_0_6838), .A2(n_8_0_6646), .ZN(n_8_0_6564));
   AOI21_X1 i_8_0_6819 (.A(n_8_0_7043), .B1(n_8_0_7042), .B2(n_8_0_7041), 
      .ZN(n_8_0_6565));
   OAI21_X1 i_8_0_6820 (.A(\out_bs[3] [2]), .B1(\out_bs[3] [1]), .B2(
      \out_bs[3] [0]), .ZN(n_8_0_6566));
   NAND3_X1 i_8_0_6824 (.A1(n_8_0_6617), .A2(n_8_0_6600), .A3(n_8_0_6570), 
      .ZN(n_8_0_6569));
   OAI211_X1 i_8_0_6825 (.A(n_8_0_6573), .B(n_8_0_6571), .C1(n_8_0_6838), 
      .C2(n_8_0_6580), .ZN(n_8_0_6570));
   NAND2_X1 i_8_0_6826 (.A1(n_8_0_6837), .A2(n_8_0_6658), .ZN(n_8_0_6571));
   NOR2_X1 i_8_0_6827 (.A1(n_8_0_6838), .A2(n_8_0_6659), .ZN(n_8_0_6572));
   OAI21_X1 i_8_0_6828 (.A(n_8_0_251), .B1(n_8_0_6579), .B2(n_8_0_6575), 
      .ZN(n_8_0_6573));
   NAND2_X1 i_8_0_6829 (.A1(n_8_0_6648), .A2(n_8_0_6576), .ZN(n_8_0_6574));
   NAND2_X1 i_8_0_6830 (.A1(n_8_0_6843), .A2(n_8_0_6659), .ZN(n_8_0_6575));
   NOR2_X1 i_8_0_6831 (.A1(n_8_0_6844), .A2(n_8_0_6658), .ZN(n_8_0_6576));
   NAND2_X1 i_8_0_6832 (.A1(\out_bs[3] [6]), .A2(n_8_0_6843), .ZN(n_8_0_6577));
   NOR2_X1 i_8_0_6833 (.A1(n_8_0_7047), .A2(n_8_0_6844), .ZN(n_8_0_6578));
   NAND2_X1 i_8_0_6834 (.A1(n_8_0_6653), .A2(n_8_0_6648), .ZN(n_8_0_6579));
   NOR2_X1 i_8_0_6835 (.A1(n_8_0_6652), .A2(n_8_0_6647), .ZN(n_8_0_6580));
   INV_X1 i_8_0_6836 (.A(n_8_0_6582), .ZN(n_8_0_6581));
   OAI21_X1 i_8_0_6838 (.A(n_8_0_6755), .B1(n_8_0_6752), .B2(n_8_0_6750), 
      .ZN(n_8_0_6583));
   AOI21_X1 i_8_0_6839 (.A(n_8_0_6754), .B1(n_8_0_6753), .B2(n_8_0_6751), 
      .ZN(n_8_0_6584));
   NAND2_X1 i_8_0_6840 (.A1(n_8_0_6742), .A2(n_8_0_6589), .ZN(n_8_0_6585));
   NAND2_X1 i_8_0_6841 (.A1(n_8_0_6751), .A2(n_8_0_6589), .ZN(n_8_0_6586));
   NAND2_X1 i_8_0_6842 (.A1(\out_bs[6] [4]), .A2(n_8_0_6589), .ZN(n_8_0_6587));
   NAND2_X1 i_8_0_6843 (.A1(n_8_0_6759), .A2(n_8_0_6753), .ZN(n_8_0_6588));
   NOR2_X1 i_8_0_6844 (.A1(n_8_0_6758), .A2(n_8_0_6752), .ZN(n_8_0_6589));
   NAND2_X1 i_8_0_6845 (.A1(\out_bs[6] [6]), .A2(n_8_0_6759), .ZN(n_8_0_6590));
   NOR2_X1 i_8_0_6846 (.A1(n_8_0_7012), .A2(n_8_0_6758), .ZN(n_8_0_6591));
   AOI221_X1 i_8_0_6847 (.A(n_8_0_6595), .B1(n_8_0_6593), .B2(n_8_0_6811), 
      .C1(n_8_0_6598), .C2(n_8_0_62), .ZN(n_8_0_6592));
   NAND2_X1 i_8_0_6849 (.A1(n_8_0_6811), .A2(n_8_0_6670), .ZN(n_8_0_6594));
   NAND2_X1 i_8_0_6851 (.A1(n_8_0_6810), .A2(\out_bs[0] [5]), .ZN(n_8_0_6596));
   NAND3_X1 i_8_0_6853 (.A1(n_8_0_6810), .A2(n_8_0_6668), .A3(n_8_0_6661), 
      .ZN(n_8_0_6598));
   NAND2_X1 i_8_0_6854 (.A1(n_8_0_6810), .A2(n_8_0_6661), .ZN(n_8_0_6599));
   OAI21_X1 i_8_0_6855 (.A(n_8_0_6601), .B1(n_8_0_6781), .B2(n_8_0_6963), 
      .ZN(n_8_0_6600));
   OAI22_X1 i_8_0_6856 (.A1(n_8_0_125), .A2(n_8_0_6782), .B1(n_8_0_6699), 
      .B2(n_8_0_6692), .ZN(n_8_0_6601));
   AOI21_X1 i_8_0_6858 (.A(n_8_0_6773), .B1(n_8_0_6712), .B2(n_8_0_6611), 
      .ZN(n_8_0_6603));
   NAND2_X1 i_8_0_6859 (.A1(n_8_0_6773), .A2(n_8_0_6712), .ZN(n_8_0_6604));
   NOR2_X1 i_8_0_6860 (.A1(n_8_0_6772), .A2(n_8_0_6711), .ZN(n_8_0_6605));
   NAND2_X1 i_8_0_6861 (.A1(\out_bs[2] [6]), .A2(n_8_0_6773), .ZN(n_8_0_6606));
   NOR2_X1 i_8_0_6862 (.A1(n_8_0_7060), .A2(n_8_0_6772), .ZN(n_8_0_6607));
   INV_X1 i_8_0_6863 (.A(n_8_0_6609), .ZN(n_8_0_6608));
   NAND2_X1 i_8_0_6864 (.A1(n_8_0_6712), .A2(n_8_0_6709), .ZN(n_8_0_6609));
   NAND2_X1 i_8_0_6865 (.A1(n_8_0_6709), .A2(n_8_0_6613), .ZN(n_8_0_6610));
   NOR2_X1 i_8_0_6866 (.A1(n_8_0_6708), .A2(n_8_0_6612), .ZN(n_8_0_6611));
   NAND2_X1 i_8_0_6867 (.A1(\out_bs[2] [2]), .A2(\out_bs[2] [1]), .ZN(n_8_0_6612));
   NOR2_X1 i_8_0_6868 (.A1(n_8_0_7056), .A2(n_8_0_7055), .ZN(n_8_0_6613));
   AOI22_X1 i_8_0_6872 (.A1(n_8_0_6825), .A2(n_8_0_6895), .B1(n_8_0_6618), 
      .B2(n_8_0_6684), .ZN(n_8_0_6617));
   AOI21_X1 i_8_0_6873 (.A(n_8_0_6675), .B1(n_8_0_6619), .B2(n_8_0_377), 
      .ZN(n_8_0_6618));
   NAND2_X1 i_8_0_6874 (.A1(n_8_0_6830), .A2(\out_as[5] [6]), .ZN(n_8_0_6619));
   AOI21_X1 i_8_0_6875 (.A(n_8_0_6621), .B1(n_8_0_6795), .B2(n_8_0_314), 
      .ZN(n_8_0_6620));
   AOI22_X1 i_8_0_6876 (.A1(n_8_0_6904), .A2(n_8_0_6794), .B1(n_8_0_6643), 
      .B2(n_8_0_6624), .ZN(n_8_0_6621));
   NAND2_X1 i_8_0_6877 (.A1(n_8_0_6794), .A2(\out_bs[4] [4]), .ZN(n_8_0_6622));
   NOR2_X1 i_8_0_6878 (.A1(n_8_0_6795), .A2(n_8_0_7033), .ZN(n_8_0_6623));
   NOR2_X1 i_8_0_6879 (.A1(n_8_0_6635), .A2(n_8_0_6632), .ZN(n_8_0_6624));
   AOI21_X1 i_8_0_6880 (.A(n_8_0_6853), .B1(n_8_0_6770), .B2(n_8_0_6625), 
      .ZN(n_186));
   NOR4_X1 i_8_0_6881 (.A1(n_8_0_6713), .A2(n_8_0_6626), .A3(n_8_0_6687), 
      .A4(n_8_0_6644), .ZN(n_8_0_6625));
   NAND4_X1 i_8_0_6882 (.A1(n_8_0_6739), .A2(n_8_0_6701), .A3(n_8_0_6672), 
      .A4(n_8_0_6627), .ZN(n_8_0_6626));
   NAND2_X1 i_8_0_6883 (.A1(n_8_0_6636), .A2(n_8_0_6628), .ZN(n_8_0_6627));
   NOR2_X1 i_8_0_6884 (.A1(n_8_0_6632), .A2(n_8_0_6629), .ZN(n_8_0_6628));
   NAND2_X1 i_8_0_6885 (.A1(\out_bs[4] [0]), .A2(n_8_0_6643), .ZN(n_8_0_6629));
   NAND2_X1 i_8_0_6886 (.A1(\out_bs[4] [2]), .A2(\out_bs[4] [0]), .ZN(n_8_0_6630));
   NOR2_X1 i_8_0_6887 (.A1(n_8_0_7031), .A2(n_8_0_6632), .ZN(n_8_0_6631));
   NAND2_X1 i_8_0_6888 (.A1(\out_bs[4] [4]), .A2(\out_bs[4] [3]), .ZN(n_8_0_6632));
   NOR2_X1 i_8_0_6889 (.A1(n_8_0_7033), .A2(n_8_0_7032), .ZN(n_8_0_6633));
   NAND2_X1 i_8_0_6890 (.A1(\out_bs[4] [6]), .A2(n_8_0_6637), .ZN(n_8_0_6634));
   NAND2_X1 i_8_0_6891 (.A1(\out_bs[4] [6]), .A2(\out_bs[4] [5]), .ZN(n_8_0_6635));
   NOR2_X1 i_8_0_6892 (.A1(n_8_0_7035), .A2(n_8_0_7034), .ZN(n_8_0_6636));
   INV_X1 i_8_0_6893 (.A(n_8_0_6638), .ZN(n_8_0_6637));
   NAND2_X1 i_8_0_6894 (.A1(\out_bs[4] [5]), .A2(\out_bs[4] [4]), .ZN(n_8_0_6638));
   NAND2_X1 i_8_0_6895 (.A1(\out_bs[4] [1]), .A2(\out_bs[4] [0]), .ZN(n_8_0_6639));
   NOR2_X1 i_8_0_6896 (.A1(n_8_0_7032), .A2(n_8_0_6642), .ZN(n_8_0_6640));
   NAND2_X1 i_8_0_6897 (.A1(\out_bs[4] [3]), .A2(\out_bs[4] [2]), .ZN(n_8_0_6641));
   NAND2_X1 i_8_0_6898 (.A1(\out_bs[4] [2]), .A2(\out_bs[4] [1]), .ZN(n_8_0_6642));
   AND2_X1 i_8_0_6899 (.A1(\out_bs[4] [2]), .A2(\out_bs[4] [1]), .ZN(n_8_0_6643));
   OAI22_X1 i_8_0_6900 (.A1(n_8_0_6665), .A2(n_8_0_6660), .B1(n_8_0_6649), 
      .B2(n_8_0_6645), .ZN(n_8_0_6644));
   NAND2_X1 i_8_0_6901 (.A1(n_8_0_6659), .A2(n_8_0_6648), .ZN(n_8_0_6645));
   NOR2_X1 i_8_0_6902 (.A1(n_8_0_6658), .A2(n_8_0_6647), .ZN(n_8_0_6646));
   NAND2_X1 i_8_0_6903 (.A1(\out_bs[3] [4]), .A2(\out_bs[3] [3]), .ZN(n_8_0_6647));
   NOR2_X1 i_8_0_6904 (.A1(n_8_0_7045), .A2(n_8_0_7044), .ZN(n_8_0_6648));
   NAND2_X1 i_8_0_6905 (.A1(\out_bs[3] [0]), .A2(n_8_0_6653), .ZN(n_8_0_6649));
   NOR2_X1 i_8_0_6906 (.A1(n_8_0_7041), .A2(n_8_0_6652), .ZN(n_8_0_6650));
   NAND2_X1 i_8_0_6907 (.A1(\out_bs[3] [1]), .A2(\out_bs[3] [0]), .ZN(n_8_0_6651));
   NAND2_X1 i_8_0_6908 (.A1(\out_bs[3] [2]), .A2(\out_bs[3] [1]), .ZN(n_8_0_6652));
   NOR2_X1 i_8_0_6909 (.A1(n_8_0_7043), .A2(n_8_0_7042), .ZN(n_8_0_6653));
   NAND2_X1 i_8_0_6910 (.A1(\out_bs[3] [4]), .A2(n_8_0_6659), .ZN(n_8_0_6654));
   NOR2_X1 i_8_0_6911 (.A1(n_8_0_7045), .A2(n_8_0_6658), .ZN(n_8_0_6655));
   NAND2_X1 i_8_0_6912 (.A1(\out_bs[3] [6]), .A2(\out_bs[3] [4]), .ZN(n_8_0_6656));
   NOR2_X1 i_8_0_6913 (.A1(n_8_0_7047), .A2(n_8_0_7045), .ZN(n_8_0_6657));
   NAND2_X1 i_8_0_6914 (.A1(\out_bs[3] [6]), .A2(\out_bs[3] [5]), .ZN(n_8_0_6658));
   NOR2_X1 i_8_0_6915 (.A1(n_8_0_7047), .A2(n_8_0_7046), .ZN(n_8_0_6659));
   NAND2_X1 i_8_0_6916 (.A1(n_8_0_6671), .A2(n_8_0_6663), .ZN(n_8_0_6660));
   NOR2_X1 i_8_0_6917 (.A1(n_8_0_6670), .A2(n_8_0_6662), .ZN(n_8_0_6661));
   NAND2_X1 i_8_0_6918 (.A1(\out_bs[0] [4]), .A2(\out_bs[0] [3]), .ZN(n_8_0_6662));
   NOR2_X1 i_8_0_6919 (.A1(n_8_0_7083), .A2(n_8_0_7082), .ZN(n_8_0_6663));
   NOR2_X1 i_8_0_6920 (.A1(n_8_0_7082), .A2(n_8_0_6665), .ZN(n_8_0_6664));
   NAND2_X1 i_8_0_6921 (.A1(\out_bs[0] [0]), .A2(n_8_0_6668), .ZN(n_8_0_6665));
   NOR2_X1 i_8_0_6922 (.A1(n_8_0_7079), .A2(n_8_0_6667), .ZN(n_8_0_6666));
   NAND2_X1 i_8_0_6923 (.A1(\out_bs[0] [2]), .A2(\out_bs[0] [1]), .ZN(n_8_0_6667));
   NOR2_X1 i_8_0_6924 (.A1(n_8_0_7081), .A2(n_8_0_7080), .ZN(n_8_0_6668));
   NAND2_X1 i_8_0_6925 (.A1(\out_bs[0] [4]), .A2(n_8_0_6671), .ZN(n_8_0_6669));
   NAND2_X1 i_8_0_6926 (.A1(\out_bs[0] [6]), .A2(\out_bs[0] [5]), .ZN(n_8_0_6670));
   NOR2_X1 i_8_0_6927 (.A1(n_8_0_7085), .A2(n_8_0_7084), .ZN(n_8_0_6671));
   NAND2_X1 i_8_0_6928 (.A1(n_8_0_6684), .A2(n_8_0_6674), .ZN(n_8_0_6672));
   NAND2_X1 i_8_0_6929 (.A1(\out_bs[5] [0]), .A2(n_8_0_6676), .ZN(n_8_0_6673));
   NOR2_X1 i_8_0_6930 (.A1(n_8_0_6678), .A2(n_8_0_6677), .ZN(n_8_0_6674));
   NAND2_X1 i_8_0_6931 (.A1(\out_bs[5] [1]), .A2(n_8_0_6679), .ZN(n_8_0_6675));
   NOR2_X1 i_8_0_6932 (.A1(n_8_0_7019), .A2(n_8_0_6678), .ZN(n_8_0_6676));
   NAND2_X1 i_8_0_6933 (.A1(\out_bs[5] [1]), .A2(\out_bs[5] [0]), .ZN(n_8_0_6677));
   NAND2_X1 i_8_0_6934 (.A1(\out_bs[5] [3]), .A2(\out_bs[5] [2]), .ZN(n_8_0_6678));
   NOR2_X1 i_8_0_6935 (.A1(n_8_0_7021), .A2(n_8_0_7020), .ZN(n_8_0_6679));
   NAND2_X1 i_8_0_6936 (.A1(\out_bs[5] [3]), .A2(\out_bs[5] [0]), .ZN(n_8_0_6680));
   NAND2_X1 i_8_0_6937 (.A1(\out_bs[5] [2]), .A2(\out_bs[5] [1]), .ZN(n_8_0_6681));
   NOR2_X1 i_8_0_6938 (.A1(n_8_0_7020), .A2(n_8_0_7019), .ZN(n_8_0_6682));
   NAND2_X1 i_8_0_6939 (.A1(\out_bs[5] [5]), .A2(n_8_0_6686), .ZN(n_8_0_6683));
   NOR2_X1 i_8_0_6940 (.A1(n_8_0_7022), .A2(n_8_0_6685), .ZN(n_8_0_6684));
   NAND2_X1 i_8_0_6941 (.A1(\out_bs[5] [6]), .A2(\out_bs[5] [5]), .ZN(n_8_0_6685));
   NOR2_X1 i_8_0_6942 (.A1(n_8_0_7024), .A2(n_8_0_7022), .ZN(n_8_0_6686));
   NOR2_X1 i_8_0_6943 (.A1(n_8_0_6697), .A2(n_8_0_6692), .ZN(n_8_0_6687));
   NOR2_X1 i_8_0_6944 (.A1(n_8_0_6697), .A2(n_8_0_6695), .ZN(n_8_0_6688));
   NAND2_X1 i_8_0_6945 (.A1(\out_bs[1] [2]), .A2(n_8_0_6696), .ZN(n_8_0_6689));
   NAND2_X1 i_8_0_6946 (.A1(\out_bs[1] [1]), .A2(\out_bs[1] [0]), .ZN(n_8_0_6690));
   INV_X1 i_8_0_6947 (.A(n_8_0_6692), .ZN(n_8_0_6691));
   NAND2_X1 i_8_0_6948 (.A1(n_8_0_6696), .A2(n_8_0_6694), .ZN(n_8_0_6692));
   NAND2_X1 i_8_0_6949 (.A1(\out_bs[1] [6]), .A2(\out_bs[1] [5]), .ZN(n_8_0_6693));
   NOR2_X1 i_8_0_6950 (.A1(n_8_0_7072), .A2(n_8_0_7071), .ZN(n_8_0_6694));
   NAND2_X1 i_8_0_6951 (.A1(\out_bs[1] [4]), .A2(\out_bs[1] [3]), .ZN(n_8_0_6695));
   NOR2_X1 i_8_0_6952 (.A1(n_8_0_7070), .A2(n_8_0_7069), .ZN(n_8_0_6696));
   NAND2_X1 i_8_0_6953 (.A1(\out_bs[1] [0]), .A2(n_8_0_6700), .ZN(n_8_0_6697));
   NAND2_X1 i_8_0_6954 (.A1(\out_bs[1] [2]), .A2(\out_bs[1] [0]), .ZN(n_8_0_6698));
   NAND2_X1 i_8_0_6955 (.A1(\out_bs[1] [2]), .A2(\out_bs[1] [1]), .ZN(n_8_0_6699));
   NOR2_X1 i_8_0_6956 (.A1(n_8_0_7068), .A2(n_8_0_7067), .ZN(n_8_0_6700));
   NAND2_X1 i_8_0_6957 (.A1(n_8_0_6712), .A2(n_8_0_6704), .ZN(n_8_0_6701));
   NAND2_X1 i_8_0_6958 (.A1(\out_bs[2] [4]), .A2(n_8_0_6712), .ZN(n_8_0_6702));
   INV_X1 i_8_0_6959 (.A(n_8_0_6704), .ZN(n_8_0_6703));
   AND2_X1 i_8_0_6960 (.A1(n_8_0_6710), .A2(n_8_0_6707), .ZN(n_8_0_6704));
   NAND2_X1 i_8_0_6961 (.A1(\out_bs[2] [4]), .A2(n_8_0_6710), .ZN(n_8_0_6705));
   NAND2_X1 i_8_0_6962 (.A1(\out_bs[2] [2]), .A2(n_8_0_6709), .ZN(n_8_0_6706));
   NOR2_X1 i_8_0_6963 (.A1(n_8_0_7056), .A2(n_8_0_6708), .ZN(n_8_0_6707));
   NAND2_X1 i_8_0_6964 (.A1(\out_bs[2] [4]), .A2(\out_bs[2] [3]), .ZN(n_8_0_6708));
   NOR2_X1 i_8_0_6965 (.A1(n_8_0_7058), .A2(n_8_0_7057), .ZN(n_8_0_6709));
   NOR2_X1 i_8_0_6966 (.A1(n_8_0_7055), .A2(n_8_0_7054), .ZN(n_8_0_6710));
   NAND2_X1 i_8_0_6967 (.A1(\out_bs[2] [6]), .A2(\out_bs[2] [5]), .ZN(n_8_0_6711));
   NOR2_X1 i_8_0_6968 (.A1(n_8_0_7060), .A2(n_8_0_7059), .ZN(n_8_0_6712));
   OAI21_X1 i_8_0_6969 (.A(n_8_0_6730), .B1(n_8_0_6722), .B2(n_8_0_6714), 
      .ZN(n_8_0_6713));
   NAND2_X1 i_8_0_6972 (.A1(\out_bs[7] [6]), .A2(\out_bs[7] [4]), .ZN(n_8_0_6716));
   NOR2_X1 i_8_0_6973 (.A1(n_8_0_7000), .A2(n_8_0_6998), .ZN(n_8_0_6717));
   NOR2_X1 i_8_0_6974 (.A1(n_8_0_6729), .A2(n_8_0_6728), .ZN(n_8_0_6718));
   NAND2_X1 i_8_0_6978 (.A1(\out_bs[7] [0]), .A2(n_8_0_6725), .ZN(n_8_0_6722));
   AND2_X1 i_8_0_6979 (.A1(\out_bs[7] [0]), .A2(n_8_0_6725), .ZN(n_8_0_6723));
   AND2_X1 i_8_0_6981 (.A1(\out_bs[7] [2]), .A2(\out_bs[7] [1]), .ZN(n_8_0_6725));
   AND2_X1 i_8_0_6982 (.A1(\out_bs[7] [1]), .A2(\out_bs[7] [0]), .ZN(n_8_0_6726));
   NOR2_X1 i_8_0_6984 (.A1(n_8_0_7000), .A2(n_8_0_6999), .ZN(n_8_0_6728));
   NOR2_X1 i_8_0_6995 (.A1(n_8_0_6754), .A2(n_8_0_6740), .ZN(n_8_0_6739));
   NOR3_X1 i_8_0_6996 (.A1(n_8_0_6752), .A2(n_8_0_6748), .A3(n_8_0_6745), 
      .ZN(n_8_0_6740));
   NAND2_X1 i_8_0_6997 (.A1(n_8_0_6751), .A2(n_8_0_6744), .ZN(n_8_0_6741));
   NOR2_X1 i_8_0_6998 (.A1(n_8_0_6750), .A2(n_8_0_6743), .ZN(n_8_0_6742));
   NAND2_X1 i_8_0_6999 (.A1(\out_bs[6] [2]), .A2(\out_bs[6] [1]), .ZN(n_8_0_6743));
   NOR2_X1 i_8_0_7000 (.A1(n_8_0_7008), .A2(n_8_0_7007), .ZN(n_8_0_6744));
   NAND2_X1 i_8_0_7001 (.A1(\out_bs[6] [1]), .A2(\out_bs[6] [0]), .ZN(n_8_0_6745));
   NOR2_X1 i_8_0_7002 (.A1(n_8_0_7007), .A2(n_8_0_7006), .ZN(n_8_0_6746));
   NAND2_X1 i_8_0_7003 (.A1(\out_bs[6] [4]), .A2(n_8_0_6753), .ZN(n_8_0_6747));
   NAND2_X1 i_8_0_7004 (.A1(\out_bs[6] [2]), .A2(n_8_0_6751), .ZN(n_8_0_6748));
   NOR2_X1 i_8_0_7005 (.A1(n_8_0_7008), .A2(n_8_0_6750), .ZN(n_8_0_6749));
   NAND2_X1 i_8_0_7006 (.A1(\out_bs[6] [4]), .A2(\out_bs[6] [3]), .ZN(n_8_0_6750));
   NOR2_X1 i_8_0_7007 (.A1(n_8_0_7010), .A2(n_8_0_7009), .ZN(n_8_0_6751));
   NOR2_X1 i_8_0_7009 (.A1(n_8_0_7012), .A2(n_8_0_7011), .ZN(n_8_0_6753));
   NAND2_X1 i_8_0_7010 (.A1(n_8_0_6758), .A2(n_8_0_6756), .ZN(n_8_0_6754));
   INV_X1 i_8_0_7012 (.A(n_8_0_6757), .ZN(n_8_0_6756));
   NOR2_X1 i_8_0_7013 (.A1(\out_bs[6] [6]), .A2(n_8_0_6761), .ZN(n_8_0_6757));
   NAND2_X1 i_8_0_7014 (.A1(n_8_0_6760), .A2(\out_as[6] [6]), .ZN(n_8_0_6758));
   NOR2_X1 i_8_0_7015 (.A1(n_8_0_6761), .A2(n_8_0_7018), .ZN(n_8_0_6759));
   OAI21_X1 i_8_0_7016 (.A(n_8_0_6763), .B1(\out_bs[6] [6]), .B2(n_8_0_7018), 
      .ZN(n_8_0_6760));
   AOI21_X1 i_8_0_7017 (.A(n_8_0_6762), .B1(n_8_0_7012), .B2(\out_as[6] [6]), 
      .ZN(n_8_0_6761));
   NAND2_X1 i_8_0_7018 (.A1(n_8_0_6765), .A2(n_8_0_6764), .ZN(n_8_0_6762));
   AND2_X1 i_8_0_7019 (.A1(n_8_0_6765), .A2(n_8_0_6764), .ZN(n_8_0_6763));
   NAND2_X1 i_8_0_7020 (.A1(n_8_0_7011), .A2(\out_as[6] [5]), .ZN(n_8_0_6764));
   OAI221_X1 i_8_0_7021 (.A(n_8_0_6766), .B1(n_8_0_7010), .B2(\out_as[6] [4]), 
      .C1(\out_as[6] [5]), .C2(n_8_0_7011), .ZN(n_8_0_6765));
   OAI221_X1 i_8_0_7022 (.A(n_8_0_6767), .B1(\out_bs[6] [3]), .B2(n_8_0_7015), 
      .C1(n_8_0_7016), .C2(\out_bs[6] [4]), .ZN(n_8_0_6766));
   OAI221_X1 i_8_0_7023 (.A(n_8_0_6768), .B1(n_8_0_7008), .B2(\out_as[6] [2]), 
      .C1(\out_as[6] [3]), .C2(n_8_0_7009), .ZN(n_8_0_6767));
   OAI221_X1 i_8_0_7024 (.A(n_8_0_6769), .B1(\out_bs[6] [1]), .B2(n_8_0_7013), 
      .C1(n_8_0_7014), .C2(\out_bs[6] [2]), .ZN(n_8_0_6768));
   OAI211_X1 i_8_0_7025 (.A(\out_as[6] [0]), .B(n_8_0_7006), .C1(n_8_0_7007), 
      .C2(\out_as[6] [1]), .ZN(n_8_0_6769));
   NOR4_X1 i_8_0_7026 (.A1(n_8_0_6825), .A2(n_8_0_6810), .A3(n_8_0_6781), 
      .A4(n_8_0_6771), .ZN(n_8_0_6770));
   NAND3_X1 i_8_0_7027 (.A1(n_8_0_6795), .A2(n_8_0_6772), .A3(n_8_0_6837), 
      .ZN(n_8_0_6771));
   OAI21_X1 i_8_0_7028 (.A(n_8_0_6775), .B1(n_8_0_7060), .B2(\out_as[2] [6]), 
      .ZN(n_8_0_6772));
   AOI21_X1 i_8_0_7029 (.A(n_8_0_6774), .B1(\out_bs[2] [6]), .B2(n_8_0_7066), 
      .ZN(n_8_0_6773));
   INV_X1 i_8_0_7030 (.A(n_8_0_6775), .ZN(n_8_0_6774));
   OAI221_X1 i_8_0_7031 (.A(n_8_0_6776), .B1(\out_bs[2] [5]), .B2(n_8_0_7065), 
      .C1(n_8_0_7066), .C2(\out_bs[2] [6]), .ZN(n_8_0_6775));
   OAI221_X1 i_8_0_7032 (.A(n_8_0_6777), .B1(n_8_0_7058), .B2(\out_as[2] [4]), 
      .C1(\out_as[2] [5]), .C2(n_8_0_7059), .ZN(n_8_0_6776));
   OAI221_X1 i_8_0_7033 (.A(n_8_0_6778), .B1(\out_bs[2] [3]), .B2(n_8_0_7063), 
      .C1(n_8_0_7064), .C2(\out_bs[2] [4]), .ZN(n_8_0_6777));
   OAI221_X1 i_8_0_7034 (.A(n_8_0_6779), .B1(n_8_0_7056), .B2(\out_as[2] [2]), 
      .C1(\out_as[2] [3]), .C2(n_8_0_7057), .ZN(n_8_0_6778));
   OAI221_X1 i_8_0_7035 (.A(n_8_0_6780), .B1(\out_bs[2] [1]), .B2(n_8_0_7061), 
      .C1(n_8_0_7062), .C2(\out_bs[2] [2]), .ZN(n_8_0_6779));
   OAI211_X1 i_8_0_7036 (.A(\out_as[2] [0]), .B(n_8_0_7054), .C1(n_8_0_7055), 
      .C2(\out_as[2] [1]), .ZN(n_8_0_6780));
   OAI21_X1 i_8_0_7037 (.A(n_8_0_6784), .B1(\out_bs[1] [6]), .B2(n_8_0_7078), 
      .ZN(n_8_0_6781));
   AOI21_X1 i_8_0_7038 (.A(n_8_0_6783), .B1(n_8_0_7072), .B2(\out_as[1] [6]), 
      .ZN(n_8_0_6782));
   INV_X1 i_8_0_7039 (.A(n_8_0_6784), .ZN(n_8_0_6783));
   OAI21_X1 i_8_0_7040 (.A(n_8_0_6785), .B1(n_8_0_7072), .B2(\out_as[1] [6]), 
      .ZN(n_8_0_6784));
   OAI21_X1 i_8_0_7041 (.A(n_8_0_6787), .B1(\out_bs[1] [5]), .B2(n_8_0_7077), 
      .ZN(n_8_0_6785));
   AOI21_X1 i_8_0_7042 (.A(n_8_0_6788), .B1(n_8_0_7071), .B2(\out_as[1] [5]), 
      .ZN(n_8_0_6786));
   INV_X1 i_8_0_7043 (.A(n_8_0_6788), .ZN(n_8_0_6787));
   AOI21_X1 i_8_0_7044 (.A(n_8_0_6789), .B1(n_8_0_6791), .B2(n_8_0_6792), 
      .ZN(n_8_0_6788));
   OAI222_X1 i_8_0_7045 (.A1(n_8_0_6790), .A2(\out_as[1] [3]), .B1(n_8_0_7070), 
      .B2(\out_as[1] [4]), .C1(\out_as[1] [5]), .C2(n_8_0_7071), .ZN(n_8_0_6789));
   OAI21_X1 i_8_0_7046 (.A(\out_bs[1] [3]), .B1(n_8_0_7076), .B2(\out_bs[1] [4]), 
      .ZN(n_8_0_6790));
   AOI222_X1 i_8_0_7047 (.A1(\out_as[1] [4]), .A2(n_8_0_7070), .B1(n_8_0_7069), 
      .B2(\out_as[1] [3]), .C1(n_8_0_7068), .C2(\out_as[1] [2]), .ZN(n_8_0_6791));
   OAI221_X1 i_8_0_7048 (.A(n_8_0_6793), .B1(n_8_0_7067), .B2(\out_as[1] [1]), 
      .C1(\out_as[1] [2]), .C2(n_8_0_7068), .ZN(n_8_0_6792));
   OAI22_X1 i_8_0_7049 (.A1(n_8_0_7074), .A2(\out_bs[1] [1]), .B1(n_8_0_7073), 
      .B2(\out_bs[1] [0]), .ZN(n_8_0_6793));
   NAND2_X1 i_8_0_7050 (.A1(n_8_0_6798), .A2(n_8_0_6797), .ZN(n_8_0_6794));
   NOR2_X1 i_8_0_7051 (.A1(n_8_0_6799), .A2(n_8_0_6796), .ZN(n_8_0_6795));
   INV_X1 i_8_0_7052 (.A(n_8_0_6797), .ZN(n_8_0_6796));
   NAND2_X1 i_8_0_7053 (.A1(n_8_0_6800), .A2(\out_as[4] [6]), .ZN(n_8_0_6797));
   INV_X1 i_8_0_7054 (.A(n_8_0_6799), .ZN(n_8_0_6798));
   NOR2_X1 i_8_0_7055 (.A1(\out_bs[4] [6]), .A2(n_8_0_6801), .ZN(n_8_0_6799));
   NAND3_X1 i_8_0_7056 (.A1(n_8_0_6809), .A2(n_8_0_6803), .A3(n_8_0_6802), 
      .ZN(n_8_0_6800));
   AND3_X1 i_8_0_7057 (.A1(n_8_0_6809), .A2(n_8_0_6803), .A3(n_8_0_6802), 
      .ZN(n_8_0_6801));
   NAND2_X1 i_8_0_7058 (.A1(n_8_0_7034), .A2(\out_as[4] [5]), .ZN(n_8_0_6802));
   OAI221_X1 i_8_0_7059 (.A(n_8_0_6804), .B1(n_8_0_7033), .B2(\out_as[4] [4]), 
      .C1(\out_as[4] [5]), .C2(n_8_0_7034), .ZN(n_8_0_6803));
   OAI221_X1 i_8_0_7060 (.A(n_8_0_6805), .B1(\out_bs[4] [3]), .B2(n_8_0_7038), 
      .C1(n_8_0_7039), .C2(\out_bs[4] [4]), .ZN(n_8_0_6804));
   OAI221_X1 i_8_0_7061 (.A(n_8_0_6806), .B1(n_8_0_7031), .B2(\out_as[4] [2]), 
      .C1(\out_as[4] [3]), .C2(n_8_0_7032), .ZN(n_8_0_6805));
   OAI221_X1 i_8_0_7062 (.A(n_8_0_6807), .B1(\out_bs[4] [1]), .B2(n_8_0_7036), 
      .C1(n_8_0_7037), .C2(\out_bs[4] [2]), .ZN(n_8_0_6806));
   NAND2_X1 i_8_0_7063 (.A1(\out_as[4] [0]), .A2(n_8_0_6808), .ZN(n_8_0_6807));
   AOI21_X1 i_8_0_7064 (.A(\out_bs[4] [0]), .B1(n_8_0_7036), .B2(\out_bs[4] [1]), 
      .ZN(n_8_0_6808));
   NAND2_X1 i_8_0_7065 (.A1(n_8_0_7035), .A2(\out_as[4] [6]), .ZN(n_8_0_6809));
   AOI21_X1 i_8_0_7066 (.A(n_8_0_6816), .B1(\out_bs[0] [6]), .B2(n_8_0_7089), 
      .ZN(n_8_0_6810));
   NAND2_X1 i_8_0_7068 (.A1(n_8_0_6815), .A2(\out_as[0] [6]), .ZN(n_8_0_6812));
   NOR2_X1 i_8_0_7069 (.A1(n_8_0_6816), .A2(n_8_0_7089), .ZN(n_8_0_6813));
   NOR2_X1 i_8_0_7070 (.A1(\out_bs[0] [6]), .A2(n_8_0_6816), .ZN(n_8_0_6814));
   OR2_X1 i_8_0_7071 (.A1(n_8_0_6817), .A2(n_8_0_6823), .ZN(n_8_0_6815));
   NOR2_X1 i_8_0_7072 (.A1(n_8_0_6817), .A2(n_8_0_6823), .ZN(n_8_0_6816));
   OAI22_X1 i_8_0_7073 (.A1(n_8_0_6819), .A2(n_8_0_6818), .B1(n_8_0_7088), 
      .B2(\out_bs[0] [5]), .ZN(n_8_0_6817));
   OAI22_X1 i_8_0_7074 (.A1(\out_as[0] [5]), .A2(n_8_0_7084), .B1(n_8_0_7083), 
      .B2(\out_as[0] [4]), .ZN(n_8_0_6818));
   AOI221_X1 i_8_0_7075 (.A(n_8_0_6820), .B1(n_8_0_7082), .B2(\out_as[0] [3]), 
      .C1(\out_as[0] [4]), .C2(n_8_0_7083), .ZN(n_8_0_6819));
   AOI222_X1 i_8_0_7076 (.A1(n_8_0_6821), .A2(n_8_0_6822), .B1(\out_bs[0] [3]), 
      .B2(n_8_0_7087), .C1(\out_bs[0] [2]), .C2(n_8_0_7086), .ZN(n_8_0_6820));
   AOI22_X1 i_8_0_7077 (.A1(\out_as[0] [2]), .A2(n_8_0_7081), .B1(n_8_0_7080), 
      .B2(\out_as[0] [1]), .ZN(n_8_0_6821));
   OAI211_X1 i_8_0_7078 (.A(\out_as[0] [0]), .B(n_8_0_7079), .C1(n_8_0_7080), 
      .C2(\out_as[0] [1]), .ZN(n_8_0_6822));
   NOR2_X1 i_8_0_7079 (.A1(n_8_0_7089), .A2(\out_bs[0] [6]), .ZN(n_8_0_6823));
   NAND2_X1 i_8_0_7080 (.A1(n_8_0_6826), .A2(n_8_0_6829), .ZN(n_8_0_6824));
   AND2_X1 i_8_0_7081 (.A1(n_8_0_6826), .A2(n_8_0_6829), .ZN(n_8_0_6825));
   OAI21_X1 i_8_0_7082 (.A(n_8_0_7030), .B1(\out_bs[5] [6]), .B2(n_8_0_6831), 
      .ZN(n_8_0_6826));
   NAND2_X1 i_8_0_7083 (.A1(n_8_0_6831), .A2(n_8_0_7030), .ZN(n_8_0_6827));
   NOR2_X1 i_8_0_7084 (.A1(n_8_0_6830), .A2(\out_as[5] [6]), .ZN(n_8_0_6828));
   NAND2_X1 i_8_0_7085 (.A1(\out_bs[5] [6]), .A2(n_8_0_6831), .ZN(n_8_0_6829));
   INV_X1 i_8_0_7086 (.A(n_8_0_6831), .ZN(n_8_0_6830));
   AOI21_X1 i_8_0_7087 (.A(n_8_0_6832), .B1(n_8_0_7023), .B2(\out_as[5] [5]), 
      .ZN(n_8_0_6831));
   AOI221_X1 i_8_0_7088 (.A(n_8_0_6833), .B1(\out_bs[5] [4]), .B2(n_8_0_7028), 
      .C1(n_8_0_7029), .C2(\out_bs[5] [5]), .ZN(n_8_0_6832));
   AOI221_X1 i_8_0_7089 (.A(n_8_0_6834), .B1(n_8_0_7021), .B2(\out_as[5] [3]), 
      .C1(\out_as[5] [4]), .C2(n_8_0_7022), .ZN(n_8_0_6833));
   AOI221_X1 i_8_0_7090 (.A(n_8_0_6835), .B1(\out_bs[5] [2]), .B2(n_8_0_7026), 
      .C1(n_8_0_7027), .C2(\out_bs[5] [3]), .ZN(n_8_0_6834));
   AOI222_X1 i_8_0_7091 (.A1(\out_as[5] [0]), .A2(n_8_0_6836), .B1(n_8_0_7020), 
      .B2(\out_as[5] [2]), .C1(n_8_0_7019), .C2(\out_as[5] [1]), .ZN(n_8_0_6835));
   AOI21_X1 i_8_0_7092 (.A(\out_bs[5] [0]), .B1(n_8_0_7025), .B2(\out_bs[5] [1]), 
      .ZN(n_8_0_6836));
   OAI21_X1 i_8_0_7093 (.A(n_8_0_6839), .B1(n_8_0_6841), .B2(\out_as[3] [6]), 
      .ZN(n_8_0_6837));
   OAI21_X1 i_8_0_7094 (.A(n_8_0_6842), .B1(\out_bs[3] [6]), .B2(n_8_0_7053), 
      .ZN(n_8_0_6838));
   NAND2_X1 i_8_0_7095 (.A1(n_8_0_6845), .A2(\out_bs[3] [6]), .ZN(n_8_0_6839));
   NOR2_X1 i_8_0_7096 (.A1(n_8_0_6841), .A2(\out_as[3] [6]), .ZN(n_8_0_6840));
   AOI21_X1 i_8_0_7097 (.A(n_8_0_6845), .B1(\out_bs[3] [6]), .B2(n_8_0_7053), 
      .ZN(n_8_0_6841));
   OAI21_X1 i_8_0_7098 (.A(n_8_0_6846), .B1(n_8_0_7047), .B2(\out_as[3] [6]), 
      .ZN(n_8_0_6842));
   INV_X1 i_8_0_7099 (.A(n_8_0_6844), .ZN(n_8_0_6843));
   NAND2_X1 i_8_0_7100 (.A1(\out_as[3] [6]), .A2(n_8_0_6846), .ZN(n_8_0_6844));
   INV_X1 i_8_0_7101 (.A(n_8_0_6846), .ZN(n_8_0_6845));
   AOI21_X1 i_8_0_7102 (.A(n_8_0_6847), .B1(\out_bs[3] [5]), .B2(n_8_0_7052), 
      .ZN(n_8_0_6846));
   AOI222_X1 i_8_0_7103 (.A1(n_8_0_6849), .A2(n_8_0_6848), .B1(\out_as[3] [5]), 
      .B2(n_8_0_7046), .C1(n_8_0_7045), .C2(\out_as[3] [4]), .ZN(n_8_0_6847));
   AOI22_X1 i_8_0_7104 (.A1(n_8_0_7051), .A2(\out_bs[3] [4]), .B1(n_8_0_7050), 
      .B2(\out_bs[3] [3]), .ZN(n_8_0_6848));
   OAI21_X1 i_8_0_7105 (.A(n_8_0_6850), .B1(\out_bs[3] [3]), .B2(n_8_0_7050), 
      .ZN(n_8_0_6849));
   OAI21_X1 i_8_0_7106 (.A(n_8_0_6851), .B1(n_8_0_7043), .B2(\out_as[3] [2]), 
      .ZN(n_8_0_6850));
   OAI221_X1 i_8_0_7107 (.A(n_8_0_6852), .B1(\out_bs[3] [1]), .B2(n_8_0_7048), 
      .C1(n_8_0_7049), .C2(\out_bs[3] [2]), .ZN(n_8_0_6851));
   OAI211_X1 i_8_0_7108 (.A(\out_as[3] [0]), .B(n_8_0_7041), .C1(n_8_0_7042), 
      .C2(\out_as[3] [1]), .ZN(n_8_0_6852));
   INV_X1 i_8_0_7111 (.A(n_8_0_659), .ZN(n_8_0_6855));
   INV_X1 i_8_0_7112 (.A(n_8_0_623), .ZN(n_8_0_6856));
   INV_X1 i_8_0_7113 (.A(n_8_0_597), .ZN(n_8_0_6857));
   INV_X1 i_8_0_7114 (.A(n_8_0_590), .ZN(n_8_0_6858));
   INV_X1 i_8_0_7116 (.A(n_8_0_570), .ZN(n_8_0_6860));
   INV_X1 i_8_0_7117 (.A(n_8_0_529), .ZN(n_8_0_6861));
   INV_X1 i_8_0_7118 (.A(n_8_0_502), .ZN(n_8_0_6862));
   INV_X1 i_8_0_7119 (.A(n_8_0_501), .ZN(n_8_0_6863));
   INV_X1 i_8_0_7120 (.A(n_8_0_610), .ZN(n_8_0_6864));
   INV_X1 i_8_0_7121 (.A(n_8_0_500), .ZN(n_8_0_6865));
   INV_X1 i_8_0_7123 (.A(n_8_0_498), .ZN(n_8_0_6867));
   INV_X1 i_8_0_7125 (.A(n_8_0_493), .ZN(n_8_0_6869));
   INV_X1 i_8_0_7129 (.A(n_8_0_461), .ZN(n_8_0_6873));
   INV_X1 i_8_0_7130 (.A(n_8_0_445), .ZN(n_8_0_6874));
   INV_X1 i_8_0_7131 (.A(n_8_0_444), .ZN(n_8_0_6875));
   INV_X1 i_8_0_7132 (.A(n_8_0_438), .ZN(n_8_0_6876));
   INV_X1 i_8_0_7133 (.A(n_8_0_433), .ZN(n_8_0_6877));
   INV_X1 i_8_0_7134 (.A(n_8_0_787), .ZN(n_8_0_6878));
   INV_X1 i_8_0_7135 (.A(n_8_0_425), .ZN(n_8_0_6879));
   INV_X1 i_8_0_7136 (.A(n_8_0_424), .ZN(n_8_0_6880));
   INV_X1 i_8_0_7137 (.A(n_8_0_422), .ZN(n_8_0_6881));
   INV_X1 i_8_0_7138 (.A(n_8_0_421), .ZN(n_8_0_6882));
   INV_X1 i_8_0_7139 (.A(n_8_0_419), .ZN(n_8_0_6883));
   INV_X1 i_8_0_7140 (.A(n_8_0_417), .ZN(n_8_0_6884));
   INV_X1 i_8_0_7141 (.A(n_8_0_416), .ZN(n_8_0_6885));
   INV_X1 i_8_0_7142 (.A(n_8_0_415), .ZN(n_8_0_6886));
   INV_X1 i_8_0_7143 (.A(n_8_0_921), .ZN(n_8_0_6887));
   INV_X1 i_8_0_7144 (.A(n_8_0_413), .ZN(n_8_0_6888));
   INV_X1 i_8_0_7145 (.A(n_8_0_412), .ZN(n_8_0_6889));
   INV_X1 i_8_0_7146 (.A(n_8_0_411), .ZN(n_8_0_6890));
   INV_X1 i_8_0_7147 (.A(n_8_0_953), .ZN(n_8_0_6891));
   INV_X1 i_8_0_7148 (.A(n_8_0_386), .ZN(n_8_0_6892));
   INV_X1 i_8_0_7149 (.A(n_8_0_382), .ZN(n_8_0_6893));
   INV_X1 i_8_0_7150 (.A(n_8_0_380), .ZN(n_8_0_6894));
   INV_X1 i_8_0_7151 (.A(n_8_0_377), .ZN(n_8_0_6895));
   INV_X1 i_8_0_7152 (.A(n_8_0_373), .ZN(n_8_0_6896));
   INV_X1 i_8_0_7153 (.A(n_8_0_371), .ZN(n_8_0_6897));
   INV_X1 i_8_0_7154 (.A(n_8_0_773), .ZN(n_8_0_6898));
   INV_X1 i_8_0_7155 (.A(n_8_0_821), .ZN(n_8_0_6899));
   INV_X1 i_8_0_7156 (.A(n_8_0_361), .ZN(n_8_0_6900));
   INV_X1 i_8_0_7157 (.A(n_8_0_866), .ZN(n_8_0_6901));
   INV_X1 i_8_0_7158 (.A(n_8_0_348), .ZN(n_8_0_6902));
   INV_X1 i_8_0_7159 (.A(n_8_0_317), .ZN(n_8_0_6903));
   INV_X1 i_8_0_7160 (.A(n_8_0_314), .ZN(n_8_0_6904));
   INV_X1 i_8_0_7161 (.A(n_8_0_313), .ZN(n_8_0_6905));
   INV_X1 i_8_0_7162 (.A(n_8_0_312), .ZN(n_8_0_6906));
   INV_X1 i_8_0_7163 (.A(n_8_0_619), .ZN(n_8_0_6907));
   INV_X1 i_8_0_7164 (.A(n_8_0_310), .ZN(n_8_0_6908));
   INV_X1 i_8_0_7165 (.A(n_8_0_307), .ZN(n_8_0_6909));
   INV_X1 i_8_0_7166 (.A(n_8_0_301), .ZN(n_8_0_6910));
   INV_X1 i_8_0_7167 (.A(n_8_0_835), .ZN(n_8_0_6911));
   INV_X1 i_8_0_7168 (.A(n_8_0_297), .ZN(n_8_0_6912));
   INV_X1 i_8_0_7169 (.A(n_8_0_296), .ZN(n_8_0_6913));
   INV_X1 i_8_0_7170 (.A(n_8_0_294), .ZN(n_8_0_6914));
   INV_X1 i_8_0_7171 (.A(n_8_0_289), .ZN(n_8_0_6915));
   INV_X1 i_8_0_7172 (.A(n_8_0_263), .ZN(n_8_0_6916));
   INV_X1 i_8_0_7173 (.A(n_8_0_260), .ZN(n_8_0_6917));
   INV_X1 i_8_0_7174 (.A(n_8_0_254), .ZN(n_8_0_6918));
   INV_X1 i_8_0_7175 (.A(n_8_0_249), .ZN(n_8_0_6919));
   INV_X1 i_8_0_7176 (.A(n_8_0_248), .ZN(n_8_0_6920));
   INV_X1 i_8_0_7177 (.A(n_8_0_247), .ZN(n_8_0_6921));
   INV_X1 i_8_0_7178 (.A(n_8_0_235), .ZN(n_8_0_6922));
   INV_X1 i_8_0_7179 (.A(n_8_0_234), .ZN(n_8_0_6923));
   INV_X1 i_8_0_7180 (.A(n_8_0_231), .ZN(n_8_0_6924));
   INV_X1 i_8_0_7181 (.A(n_8_0_220), .ZN(n_8_0_6925));
   INV_X1 i_8_0_7182 (.A(n_8_0_219), .ZN(n_8_0_6926));
   INV_X1 i_8_0_7183 (.A(n_8_0_216), .ZN(n_8_0_6927));
   INV_X1 i_8_0_7184 (.A(n_8_0_213), .ZN(n_8_0_6928));
   INV_X1 i_8_0_7185 (.A(n_8_0_211), .ZN(n_8_0_6929));
   INV_X1 i_8_0_7186 (.A(n_8_0_205), .ZN(n_8_0_6930));
   INV_X1 i_8_0_7187 (.A(n_8_0_203), .ZN(n_8_0_6931));
   INV_X1 i_8_0_7188 (.A(n_8_0_202), .ZN(n_8_0_6932));
   INV_X1 i_8_0_7189 (.A(n_8_0_201), .ZN(n_8_0_6933));
   INV_X1 i_8_0_7190 (.A(n_8_0_197), .ZN(n_8_0_6934));
   INV_X1 i_8_0_7191 (.A(n_8_0_195), .ZN(n_8_0_6935));
   INV_X1 i_8_0_7192 (.A(n_8_0_194), .ZN(n_8_0_6936));
   INV_X1 i_8_0_7193 (.A(n_8_0_193), .ZN(n_8_0_6937));
   INV_X1 i_8_0_7194 (.A(n_8_0_187), .ZN(n_8_0_6938));
   INV_X1 i_8_0_7195 (.A(n_8_0_185), .ZN(n_8_0_6939));
   INV_X1 i_8_0_7196 (.A(n_8_0_184), .ZN(n_8_0_6940));
   INV_X1 i_8_0_7197 (.A(n_8_0_183), .ZN(n_8_0_6941));
   INV_X1 i_8_0_7198 (.A(n_8_0_180), .ZN(n_8_0_6942));
   INV_X1 i_8_0_7199 (.A(n_8_0_179), .ZN(n_8_0_6943));
   INV_X1 i_8_0_7200 (.A(n_8_0_178), .ZN(n_8_0_6944));
   INV_X1 i_8_0_7201 (.A(n_8_0_177), .ZN(n_8_0_6945));
   INV_X1 i_8_0_7202 (.A(n_8_0_172), .ZN(n_8_0_6946));
   INV_X1 i_8_0_7203 (.A(n_8_0_171), .ZN(n_8_0_6947));
   INV_X1 i_8_0_7204 (.A(n_8_0_168), .ZN(n_8_0_6948));
   INV_X1 i_8_0_7205 (.A(n_8_0_167), .ZN(n_8_0_6949));
   INV_X1 i_8_0_7206 (.A(n_8_0_166), .ZN(n_8_0_6950));
   INV_X1 i_8_0_7207 (.A(n_8_0_165), .ZN(n_8_0_6951));
   INV_X1 i_8_0_7208 (.A(n_8_0_164), .ZN(n_8_0_6952));
   INV_X1 i_8_0_7209 (.A(n_8_0_925), .ZN(n_8_0_6953));
   INV_X1 i_8_0_7210 (.A(n_8_0_162), .ZN(n_8_0_6954));
   INV_X1 i_8_0_7211 (.A(n_8_0_159), .ZN(n_8_0_6955));
   INV_X1 i_8_0_7212 (.A(n_8_0_155), .ZN(n_8_0_6956));
   INV_X1 i_8_0_7213 (.A(n_8_0_152), .ZN(n_8_0_6957));
   INV_X1 i_8_0_7214 (.A(n_8_0_149), .ZN(n_8_0_6958));
   INV_X1 i_8_0_7215 (.A(n_8_0_141), .ZN(n_8_0_6959));
   INV_X1 i_8_0_7216 (.A(n_8_0_136), .ZN(n_8_0_6960));
   INV_X1 i_8_0_7217 (.A(n_8_0_134), .ZN(n_8_0_6961));
   INV_X1 i_8_0_7218 (.A(n_8_0_538), .ZN(n_8_0_6962));
   INV_X1 i_8_0_7219 (.A(n_8_0_125), .ZN(n_8_0_6963));
   INV_X1 i_8_0_7220 (.A(n_8_0_628), .ZN(n_8_0_6964));
   INV_X1 i_8_0_7221 (.A(n_8_0_117), .ZN(n_8_0_6965));
   INV_X1 i_8_0_7222 (.A(n_8_0_114), .ZN(n_8_0_6966));
   INV_X1 i_8_0_7223 (.A(n_8_0_113), .ZN(n_8_0_6967));
   INV_X1 i_8_0_7224 (.A(n_8_0_112), .ZN(n_8_0_6968));
   INV_X1 i_8_0_7225 (.A(n_8_0_111), .ZN(n_8_0_6969));
   INV_X1 i_8_0_7226 (.A(n_8_0_110), .ZN(n_8_0_6970));
   INV_X1 i_8_0_7227 (.A(n_8_0_846), .ZN(n_8_0_6971));
   INV_X1 i_8_0_7228 (.A(n_8_0_98), .ZN(n_8_0_6972));
   INV_X1 i_8_0_7229 (.A(n_8_0_94), .ZN(n_8_0_6973));
   INV_X1 i_8_0_7230 (.A(n_8_0_92), .ZN(n_8_0_6974));
   INV_X1 i_8_0_7231 (.A(n_8_0_90), .ZN(n_8_0_6975));
   INV_X1 i_8_0_7232 (.A(n_8_0_89), .ZN(n_8_0_6976));
   INV_X1 i_8_0_7233 (.A(n_8_0_78), .ZN(n_8_0_6977));
   INV_X1 i_8_0_7234 (.A(n_8_0_60), .ZN(n_8_0_6978));
   INV_X1 i_8_0_7235 (.A(n_8_0_719), .ZN(n_8_0_6979));
   INV_X1 i_8_0_7236 (.A(n_8_0_54), .ZN(n_8_0_6980));
   INV_X1 i_8_0_7237 (.A(n_8_0_767), .ZN(n_8_0_6981));
   INV_X1 i_8_0_7238 (.A(n_8_0_831), .ZN(n_8_0_6982));
   INV_X1 i_8_0_7239 (.A(n_8_0_41), .ZN(n_8_0_6983));
   INV_X1 i_8_0_7240 (.A(n_8_0_38), .ZN(n_8_0_6984));
   INV_X1 i_8_0_7241 (.A(n_8_0_35), .ZN(n_8_0_6985));
   INV_X1 i_8_0_7242 (.A(n_8_0_18), .ZN(n_8_0_6986));
   INV_X1 i_8_0_7246 (.A(in_data[8]), .ZN(n_8_0_6990));
   INV_X1 i_8_0_7247 (.A(in_data[12]), .ZN(n_8_0_6991));
   INV_X1 i_8_0_7248 (.A(in_data[16]), .ZN(n_8_0_6992));
   INV_X1 i_8_0_7249 (.A(in_data[20]), .ZN(n_8_0_6993));
   INV_X1 i_8_0_7250 (.A(in_data[24]), .ZN(n_8_0_6994));
   INV_X1 i_8_0_7251 (.A(in_data[28]), .ZN(n_8_0_6995));
   INV_X1 i_8_0_7258 (.A(\out_as[7] [2]), .ZN(n_8_0_7002));
   INV_X1 i_8_0_7262 (.A(\out_bs[6] [0]), .ZN(n_8_0_7006));
   INV_X1 i_8_0_7263 (.A(\out_bs[6] [1]), .ZN(n_8_0_7007));
   INV_X1 i_8_0_7264 (.A(\out_bs[6] [2]), .ZN(n_8_0_7008));
   INV_X1 i_8_0_7265 (.A(\out_bs[6] [3]), .ZN(n_8_0_7009));
   INV_X1 i_8_0_7266 (.A(\out_bs[6] [4]), .ZN(n_8_0_7010));
   INV_X1 i_8_0_7267 (.A(\out_bs[6] [5]), .ZN(n_8_0_7011));
   INV_X1 i_8_0_7268 (.A(\out_bs[6] [6]), .ZN(n_8_0_7012));
   INV_X1 i_8_0_7269 (.A(\out_as[6] [1]), .ZN(n_8_0_7013));
   INV_X1 i_8_0_7270 (.A(\out_as[6] [2]), .ZN(n_8_0_7014));
   INV_X1 i_8_0_7271 (.A(\out_as[6] [3]), .ZN(n_8_0_7015));
   INV_X1 i_8_0_7272 (.A(\out_as[6] [4]), .ZN(n_8_0_7016));
   INV_X1 i_8_0_7273 (.A(\out_as[6] [5]), .ZN(n_8_0_7017));
   INV_X1 i_8_0_7274 (.A(\out_as[6] [6]), .ZN(n_8_0_7018));
   INV_X1 i_8_0_7275 (.A(\out_bs[5] [1]), .ZN(n_8_0_7019));
   INV_X1 i_8_0_7276 (.A(\out_bs[5] [2]), .ZN(n_8_0_7020));
   INV_X1 i_8_0_7277 (.A(\out_bs[5] [3]), .ZN(n_8_0_7021));
   INV_X1 i_8_0_7278 (.A(\out_bs[5] [4]), .ZN(n_8_0_7022));
   INV_X1 i_8_0_7279 (.A(\out_bs[5] [5]), .ZN(n_8_0_7023));
   INV_X1 i_8_0_7280 (.A(\out_bs[5] [6]), .ZN(n_8_0_7024));
   INV_X1 i_8_0_7281 (.A(\out_as[5] [1]), .ZN(n_8_0_7025));
   INV_X1 i_8_0_7282 (.A(\out_as[5] [2]), .ZN(n_8_0_7026));
   INV_X1 i_8_0_7283 (.A(\out_as[5] [3]), .ZN(n_8_0_7027));
   INV_X1 i_8_0_7284 (.A(\out_as[5] [4]), .ZN(n_8_0_7028));
   INV_X1 i_8_0_7285 (.A(\out_as[5] [5]), .ZN(n_8_0_7029));
   INV_X1 i_8_0_7286 (.A(\out_as[5] [6]), .ZN(n_8_0_7030));
   INV_X1 i_8_0_7287 (.A(\out_bs[4] [2]), .ZN(n_8_0_7031));
   INV_X1 i_8_0_7288 (.A(\out_bs[4] [3]), .ZN(n_8_0_7032));
   INV_X1 i_8_0_7289 (.A(\out_bs[4] [4]), .ZN(n_8_0_7033));
   INV_X1 i_8_0_7290 (.A(\out_bs[4] [5]), .ZN(n_8_0_7034));
   INV_X1 i_8_0_7291 (.A(\out_bs[4] [6]), .ZN(n_8_0_7035));
   INV_X1 i_8_0_7292 (.A(\out_as[4] [1]), .ZN(n_8_0_7036));
   INV_X1 i_8_0_7293 (.A(\out_as[4] [2]), .ZN(n_8_0_7037));
   INV_X1 i_8_0_7294 (.A(\out_as[4] [3]), .ZN(n_8_0_7038));
   INV_X1 i_8_0_7295 (.A(\out_as[4] [4]), .ZN(n_8_0_7039));
   INV_X1 i_8_0_7296 (.A(\out_as[4] [6]), .ZN(n_8_0_7040));
   INV_X1 i_8_0_7297 (.A(\out_bs[3] [0]), .ZN(n_8_0_7041));
   INV_X1 i_8_0_7298 (.A(\out_bs[3] [1]), .ZN(n_8_0_7042));
   INV_X1 i_8_0_7299 (.A(\out_bs[3] [2]), .ZN(n_8_0_7043));
   INV_X1 i_8_0_7300 (.A(\out_bs[3] [3]), .ZN(n_8_0_7044));
   INV_X1 i_8_0_7301 (.A(\out_bs[3] [4]), .ZN(n_8_0_7045));
   INV_X1 i_8_0_7302 (.A(\out_bs[3] [5]), .ZN(n_8_0_7046));
   INV_X1 i_8_0_7303 (.A(\out_bs[3] [6]), .ZN(n_8_0_7047));
   INV_X1 i_8_0_7304 (.A(\out_as[3] [1]), .ZN(n_8_0_7048));
   INV_X1 i_8_0_7305 (.A(\out_as[3] [2]), .ZN(n_8_0_7049));
   INV_X1 i_8_0_7306 (.A(\out_as[3] [3]), .ZN(n_8_0_7050));
   INV_X1 i_8_0_7307 (.A(\out_as[3] [4]), .ZN(n_8_0_7051));
   INV_X1 i_8_0_7308 (.A(\out_as[3] [5]), .ZN(n_8_0_7052));
   INV_X1 i_8_0_7309 (.A(\out_as[3] [6]), .ZN(n_8_0_7053));
   INV_X1 i_8_0_7310 (.A(\out_bs[2] [0]), .ZN(n_8_0_7054));
   INV_X1 i_8_0_7311 (.A(\out_bs[2] [1]), .ZN(n_8_0_7055));
   INV_X1 i_8_0_7312 (.A(\out_bs[2] [2]), .ZN(n_8_0_7056));
   INV_X1 i_8_0_7313 (.A(\out_bs[2] [3]), .ZN(n_8_0_7057));
   INV_X1 i_8_0_7314 (.A(\out_bs[2] [4]), .ZN(n_8_0_7058));
   INV_X1 i_8_0_7315 (.A(\out_bs[2] [5]), .ZN(n_8_0_7059));
   INV_X1 i_8_0_7316 (.A(\out_bs[2] [6]), .ZN(n_8_0_7060));
   INV_X1 i_8_0_7317 (.A(\out_as[2] [1]), .ZN(n_8_0_7061));
   INV_X1 i_8_0_7318 (.A(\out_as[2] [2]), .ZN(n_8_0_7062));
   INV_X1 i_8_0_7319 (.A(\out_as[2] [3]), .ZN(n_8_0_7063));
   INV_X1 i_8_0_7320 (.A(\out_as[2] [4]), .ZN(n_8_0_7064));
   INV_X1 i_8_0_7321 (.A(\out_as[2] [5]), .ZN(n_8_0_7065));
   INV_X1 i_8_0_7322 (.A(\out_as[2] [6]), .ZN(n_8_0_7066));
   INV_X1 i_8_0_7323 (.A(\out_bs[1] [1]), .ZN(n_8_0_7067));
   INV_X1 i_8_0_7324 (.A(\out_bs[1] [2]), .ZN(n_8_0_7068));
   INV_X1 i_8_0_7325 (.A(\out_bs[1] [3]), .ZN(n_8_0_7069));
   INV_X1 i_8_0_7326 (.A(\out_bs[1] [4]), .ZN(n_8_0_7070));
   INV_X1 i_8_0_7327 (.A(\out_bs[1] [5]), .ZN(n_8_0_7071));
   INV_X1 i_8_0_7328 (.A(\out_bs[1] [6]), .ZN(n_8_0_7072));
   INV_X1 i_8_0_7329 (.A(\out_as[1] [0]), .ZN(n_8_0_7073));
   INV_X1 i_8_0_7330 (.A(\out_as[1] [1]), .ZN(n_8_0_7074));
   INV_X1 i_8_0_7331 (.A(\out_as[1] [2]), .ZN(n_8_0_7075));
   INV_X1 i_8_0_7332 (.A(\out_as[1] [4]), .ZN(n_8_0_7076));
   INV_X1 i_8_0_7333 (.A(\out_as[1] [5]), .ZN(n_8_0_7077));
   INV_X1 i_8_0_7334 (.A(\out_as[1] [6]), .ZN(n_8_0_7078));
   INV_X1 i_8_0_7335 (.A(\out_bs[0] [0]), .ZN(n_8_0_7079));
   INV_X1 i_8_0_7336 (.A(\out_bs[0] [1]), .ZN(n_8_0_7080));
   INV_X1 i_8_0_7337 (.A(\out_bs[0] [2]), .ZN(n_8_0_7081));
   INV_X1 i_8_0_7338 (.A(\out_bs[0] [3]), .ZN(n_8_0_7082));
   INV_X1 i_8_0_7339 (.A(\out_bs[0] [4]), .ZN(n_8_0_7083));
   INV_X1 i_8_0_7340 (.A(\out_bs[0] [5]), .ZN(n_8_0_7084));
   INV_X1 i_8_0_7341 (.A(\out_bs[0] [6]), .ZN(n_8_0_7085));
   INV_X1 i_8_0_7342 (.A(\out_as[0] [2]), .ZN(n_8_0_7086));
   INV_X1 i_8_0_7343 (.A(\out_as[0] [3]), .ZN(n_8_0_7087));
   INV_X1 i_8_0_7344 (.A(\out_as[0] [5]), .ZN(n_8_0_7088));
   INV_X1 i_8_0_7345 (.A(\out_as[0] [6]), .ZN(n_8_0_7089));
   INV_X1 i_8_0_1242 (.A(n_8_0_4315), .ZN(n_8_0_4314));
   OAI221_X1 i_8_0_1243 (.A(n_8_0_1528), .B1(n_8_0_6853), .B2(n_8_0_1529), 
      .C1(n_8_0_6469), .C2(n_8_0_1484), .ZN(n_187));
   NAND3_X1 i_8_0_1289 (.A1(n_8_0_1527), .A2(n_8_0_3885), .A3(n_8_0_6278), 
      .ZN(n_8_0_1484));
   INV_X1 i_8_0_1290 (.A(n_8_0_6998), .ZN(n_8_0_1527));
   OR3_X1 i_8_0_1291 (.A1(n_8_0_6730), .A2(n_8_0_7000), .A3(n_8_0_6853), 
      .ZN(n_8_0_1528));
   AND3_X1 i_8_0_1292 (.A1(n_8_0_1607), .A2(n_8_0_4312), .A3(n_8_0_1589), 
      .ZN(n_8_0_1529));
   NOR4_X1 i_8_0_1358 (.A1(n_8_0_4315), .A2(n_8_0_4328), .A3(n_8_0_4303), 
      .A4(n_8_0_1590), .ZN(n_8_0_1589));
   NAND2_X1 i_8_0_1359 (.A1(n_8_0_1600), .A2(n_8_0_1599), .ZN(n_8_0_1590));
   AOI21_X1 i_8_0_1360 (.A(n_8_0_4319), .B1(n_8_0_4326), .B2(n_8_0_6979), 
      .ZN(n_8_0_1599));
   INV_X1 i_8_0_1369 (.A(n_8_0_4330), .ZN(n_8_0_1600));
   OAI221_X1 i_8_0_1370 (.A(n_8_0_6606), .B1(n_8_0_6282), .B2(n_8_0_6286), 
      .C1(n_8_0_4331), .C2(n_8_0_715), .ZN(n_8_0_4330));
   OAI211_X1 i_8_0_1371 (.A(n_8_0_4304), .B(n_8_0_6577), .C1(n_8_0_4307), 
      .C2(n_8_0_5698), .ZN(n_8_0_4303));
   OAI221_X1 i_8_0_1378 (.A(n_8_0_6556), .B1(n_8_0_4484), .B2(n_8_0_6274), 
      .C1(n_8_0_4329), .C2(n_8_0_711), .ZN(n_8_0_4328));
   OAI211_X1 i_8_0_1379 (.A(n_8_0_1656), .B(n_8_0_1617), .C1(n_8_0_7422), 
      .C2(n_8_0_1616), .ZN(n_8_0_1607));
   OAI211_X1 i_8_0_1388 (.A(n_8_0_7000), .B(n_8_0_3885), .C1(n_8_0_4532), 
      .C2(n_8_0_6279), .ZN(n_8_0_1616));
   OAI21_X1 i_8_0_1389 (.A(\out_as[7] [6]), .B1(n_8_0_4532), .B2(n_8_0_6279), 
      .ZN(n_8_0_1617));
   INV_X1 i_8_0_1390 (.A(n_8_0_705), .ZN(n_8_0_1656));
   INV_X1 i_8_0_1432 (.A(n_8_0_1657), .ZN(n_8_0_4600));
   NAND2_X1 i_8_0_1433 (.A1(\out_bs[7] [5]), .A2(n_8_0_7232), .ZN(n_8_0_1657));
   INV_X1 i_8_0_1434 (.A(n_8_0_4532), .ZN(n_8_0_4531));
   INV_X1 i_8_0_1518 (.A(n_8_0_7230), .ZN(n_8_0_4597));
   INV_X1 i_8_0_1519 (.A(n_8_0_3602), .ZN(n_8_0_4501));
   OAI21_X1 i_8_0_1520 (.A(n_8_0_3375), .B1(n_8_0_4307), .B2(n_8_0_6218), 
      .ZN(n_8_0_4292));
   INV_X1 i_8_0_1521 (.A(n_8_0_3460), .ZN(n_8_0_4290));
   INV_X1 i_8_0_1522 (.A(n_8_0_3282), .ZN(n_8_0_4257));
   INV_X1 i_8_0_1539 (.A(n_8_0_3214), .ZN(n_8_0_4050));
   INV_X1 i_8_0_1540 (.A(n_8_0_3140), .ZN(n_8_0_4022));
   INV_X1 i_8_0_1541 (.A(n_8_0_1734), .ZN(n_8_0_3939));
   NAND3_X1 i_8_0_1542 (.A1(n_8_0_6467), .A2(n_8_0_6465), .A3(n_8_0_3081), 
      .ZN(n_8_0_1734));
   INV_X1 i_8_0_1562 (.A(n_8_0_3007), .ZN(n_8_0_3008));
   NOR2_X1 i_8_0_1563 (.A1(n_8_0_3006), .A2(n_8_0_3005), .ZN(n_8_0_3004));
   OAI21_X1 i_8_0_1571 (.A(n_8_0_1754), .B1(n_8_0_2755), .B2(n_8_0_1735), 
      .ZN(n_188));
   MUX2_X1 i_8_0_1572 (.A(n_8_0_1736), .B(n_8_0_6989), .S(n_8_0_2754), .Z(
      n_8_0_1735));
   OAI21_X1 i_8_0_1573 (.A(n_8_0_1737), .B1(n_8_0_3763), .B2(n_8_0_1756), 
      .ZN(n_8_0_1736));
   NAND2_X1 i_8_0_1672 (.A1(n_8_0_3763), .A2(n_8_0_1753), .ZN(n_8_0_1737));
   INV_X1 i_8_0_1673 (.A(in_data[8]), .ZN(n_8_0_1753));
   NAND2_X1 i_8_0_1683 (.A1(n_8_0_2755), .A2(in_data[0]), .ZN(n_8_0_1754));
   INV_X1 i_8_0_1684 (.A(n_8_0_1755), .ZN(n_189));
   OAI21_X1 i_8_0_1685 (.A(n_8_0_1774), .B1(n_8_0_1883), .B2(n_8_0_1782), 
      .ZN(n_8_0_1755));
   NAND2_X1 i_8_0_1706 (.A1(n_8_0_1883), .A2(n_8_0_6988), .ZN(n_8_0_1774));
   INV_X1 i_8_0_1707 (.A(n_8_0_1783), .ZN(n_8_0_1782));
   OAI21_X1 i_8_0_1708 (.A(n_8_0_1873), .B1(in_data[4]), .B2(n_8_0_4312), 
      .ZN(n_8_0_1783));
   OAI221_X1 i_8_0_1750 (.A(n_8_0_4312), .B1(n_8_0_6990), .B2(n_8_0_4314), 
      .C1(n_8_0_1947), .C2(n_8_0_1948), .ZN(n_8_0_1873));
   AOI211_X1 i_8_0_1751 (.A(n_8_0_6591), .B(n_8_0_4313), .C1(n_8_0_6291), 
      .C2(n_8_0_4349), .ZN(n_8_0_4312));
   NAND3_X1 i_8_0_1752 (.A1(n_8_0_1884), .A2(n_8_0_1607), .A3(n_8_0_6465), 
      .ZN(n_8_0_1883));
   NAND2_X1 i_8_0_1753 (.A1(n_8_0_6468), .A2(n_8_0_6278), .ZN(n_8_0_1884));
   NAND2_X1 i_8_0_1781 (.A1(n_8_0_6997), .A2(n_8_0_6722), .ZN(n_8_0_6278));
   INV_X1 i_8_0_1782 (.A(n_8_0_1904), .ZN(n_190));
   OAI21_X1 i_8_0_1783 (.A(n_8_0_3885), .B1(n_8_0_3007), .B2(n_8_0_1905), 
      .ZN(n_8_0_1904));
   OR4_X1 i_8_0_2403 (.A1(n_8_0_3006), .A2(n_8_0_3005), .A3(n_8_0_2992), 
      .A4(n_8_0_1944), .ZN(n_8_0_1905));
   NAND4_X1 i_8_0_2404 (.A1(n_8_0_2541), .A2(n_8_0_3017), .A3(n_8_0_2998), 
      .A4(n_8_0_1945), .ZN(n_8_0_1944));
   AND3_X1 i_8_0_2405 (.A1(n_8_0_3011), .A2(n_8_0_1972), .A3(n_8_0_1946), 
      .ZN(n_8_0_1945));
   OR2_X1 i_8_0_2407 (.A1(n_8_0_6811), .A2(n_8_0_3016), .ZN(n_8_0_1946));
   NAND2_X1 i_8_0_2408 (.A1(n_8_0_3003), .A2(n_8_0_1973), .ZN(n_8_0_1972));
   NOR2_X1 i_8_0_2634 (.A1(n_8_0_3206), .A2(n_8_0_701), .ZN(n_8_0_1973));
   NAND2_X1 i_8_0_2635 (.A1(n_8_0_6811), .A2(n_8_0_3016), .ZN(n_8_0_3003));
   OAI22_X1 i_8_0_2658 (.A1(n_8_0_3013), .A2(n_8_0_3012), .B1(n_8_0_4198), 
      .B2(n_8_0_5983), .ZN(n_8_0_3011));
   AOI21_X1 i_8_0_2659 (.A(n_8_0_2999), .B1(n_8_0_6838), .B2(n_8_0_3001), 
      .ZN(n_8_0_2998));
   INV_X1 i_8_0_2660 (.A(n_8_0_2994), .ZN(n_8_0_2541));
   OAI21_X1 i_8_0_2661 (.A(n_8_0_2995), .B1(n_8_0_6795), .B2(n_8_0_2997), 
      .ZN(n_8_0_2994));
   OAI221_X1 i_8_0_2662 (.A(n_8_0_3227), .B1(n_8_0_6824), .B2(n_8_0_7021), 
      .C1(n_8_0_2993), .C2(n_8_0_686), .ZN(n_8_0_2992));
   AND2_X1 i_8_0_2666 (.A1(n_8_0_2544), .A2(n_8_0_2542), .ZN(n_8_0_3007));
   NAND3_X1 i_8_0_2671 (.A1(n_8_0_6730), .A2(n_8_0_5976), .A3(n_8_0_4424), 
      .ZN(n_8_0_2542));
   OAI21_X1 i_8_0_2677 (.A(n_8_0_3010), .B1(n_8_0_680), .B2(n_8_0_3211), 
      .ZN(n_8_0_2544));
   INV_X1 i_8_0_2904 (.A(n_8_0_2545), .ZN(n_191));
   OAI21_X1 i_8_0_2905 (.A(n_8_0_3885), .B1(n_8_0_2755), .B2(n_8_0_2737), 
      .ZN(n_8_0_2545));
   OR3_X1 i_8_0_2906 (.A1(n_8_0_2754), .A2(n_8_0_3763), .A3(n_8_0_2752), 
      .ZN(n_8_0_2737));
   OR4_X1 i_8_0_2907 (.A1(n_8_0_3767), .A2(n_8_0_3752), .A3(n_8_0_3776), 
      .A4(n_8_0_3771), .ZN(n_8_0_2752));
   OAI211_X1 i_8_0_2921 (.A(n_8_0_3753), .B(n_8_0_6556), .C1(n_8_0_5573), 
      .C2(n_8_0_4484), .ZN(n_8_0_3752));
   OAI211_X1 i_8_0_2933 (.A(n_8_0_3760), .B(n_8_0_3916), .C1(n_8_0_929), 
      .C2(n_8_0_3994), .ZN(n_8_0_2754));
   OAI211_X1 i_8_0_2940 (.A(n_8_0_2756), .B(n_8_0_6465), .C1(n_8_0_928), 
      .C2(n_8_0_4595), .ZN(n_8_0_2755));
   NAND3_X1 i_8_0_2947 (.A1(n_8_0_2918), .A2(n_8_0_4598), .A3(n_8_0_5594), 
      .ZN(n_8_0_2756));
   NAND2_X1 i_8_0_2948 (.A1(n_8_0_6998), .A2(n_8_0_6117), .ZN(n_8_0_5594));
   NAND2_X1 i_8_0_2952 (.A1(n_8_0_6469), .A2(n_8_0_928), .ZN(n_8_0_2918));
   AOI21_X1 i_8_0_2995 (.A(n_8_0_6853), .B1(n_8_0_3883), .B2(n_8_0_2919), 
      .ZN(n_192));
   NOR4_X1 i_8_0_2996 (.A1(n_8_0_3871), .A2(n_8_0_3867), .A3(n_8_0_3889), 
      .A4(n_8_0_2920), .ZN(n_8_0_2919));
   OR4_X1 i_8_0_2997 (.A1(n_8_0_3874), .A2(n_8_0_3887), .A3(n_8_0_3878), 
      .A4(n_8_0_2944), .ZN(n_8_0_2920));
   OAI211_X1 i_8_0_2998 (.A(n_8_0_2946), .B(n_8_0_6249), .C1(n_8_0_903), 
      .C2(n_8_0_4514), .ZN(n_8_0_2944));
   NAND2_X1 i_8_0_3007 (.A1(n_8_0_2980), .A2(n_8_0_5724), .ZN(n_8_0_2946));
   NAND2_X1 i_8_0_3008 (.A1(n_8_0_5944), .A2(n_8_0_6665), .ZN(n_8_0_5724));
   OAI21_X1 i_8_0_3009 (.A(n_8_0_6596), .B1(n_8_0_903), .B2(n_8_0_4512), 
      .ZN(n_8_0_2980));
   OAI211_X1 i_8_0_3010 (.A(n_8_0_6526), .B(n_8_0_3880), .C1(n_8_0_3879), 
      .C2(n_8_0_902), .ZN(n_8_0_3878));
   OAI221_X1 i_8_0_3011 (.A(n_8_0_6606), .B1(n_8_0_6282), .B2(n_8_0_5707), 
      .C1(n_8_0_3888), .C2(n_8_0_901), .ZN(n_8_0_3887));
   OAI211_X1 i_8_0_3014 (.A(n_8_0_3890), .B(n_8_0_6513), .C1(n_8_0_898), 
      .C2(n_8_0_4571), .ZN(n_8_0_3889));
   OAI21_X1 i_8_0_3019 (.A(n_8_0_2989), .B1(n_8_0_6729), .B2(n_8_0_2990), 
      .ZN(n_8_0_3883));
   OAI22_X1 i_8_0_3025 (.A1(n_8_0_6730), .A2(n_8_0_2991), .B1(\out_as[7] [6]), 
      .B2(n_8_0_896), .ZN(n_8_0_2989));
   INV_X1 i_8_0_3028 (.A(n_8_0_2991), .ZN(n_8_0_2990));
   AOI21_X1 i_8_0_3029 (.A(\out_bs[7] [6]), .B1(\out_bs[7] [5]), .B2(n_8_0_5716), 
      .ZN(n_8_0_2991));
   OR4_X1 i_8_0_3033 (.A1(n_8_0_3913), .A2(n_8_0_3910), .A3(n_8_0_3908), 
      .A4(n_8_0_3893), .ZN(n_8_0_3002));
   OAI221_X1 i_8_0_3034 (.A(n_8_0_6526), .B1(n_8_0_5984), .B2(n_8_0_6321), 
      .C1(n_8_0_3894), .C2(n_8_0_894), .ZN(n_8_0_3893));
   OAI21_X1 i_8_0_3035 (.A(n_8_0_3896), .B1(n_8_0_3898), .B2(n_8_0_3897), 
      .ZN(n_8_0_3895));
   OAI21_X1 i_8_0_3038 (.A(n_8_0_3009), .B1(n_8_0_3901), .B2(n_8_0_3014), 
      .ZN(n_8_0_3899));
   OR3_X1 i_8_0_3042 (.A1(n_8_0_6831), .A2(\out_as[5] [6]), .A3(n_8_0_890), 
      .ZN(n_8_0_3009));
   OR2_X1 i_8_0_3119 (.A1(n_8_0_3900), .A2(n_8_0_4110), .ZN(n_8_0_3014));
   NOR2_X1 i_8_0_3120 (.A1(\out_bs[7] [4]), .A2(\out_bs[7] [3]), .ZN(n_8_0_5976));
   INV_X1 i_8_0_3121 (.A(n_8_0_3074), .ZN(n_193));
   NAND2_X1 i_8_0_3125 (.A1(n_8_0_3075), .A2(n_8_0_3885), .ZN(n_8_0_3074));
   NAND4_X1 i_8_0_3126 (.A1(n_8_0_6467), .A2(n_8_0_6465), .A3(n_8_0_3081), 
      .A4(n_8_0_3079), .ZN(n_8_0_3075));
   NOR3_X1 i_8_0_3127 (.A1(n_8_0_3921), .A2(n_8_0_3931), .A3(n_8_0_3080), 
      .ZN(n_8_0_3079));
   OR4_X1 i_8_0_3134 (.A1(n_8_0_3920), .A2(n_8_0_3928), .A3(n_8_0_3923), 
      .A4(n_8_0_3934), .ZN(n_8_0_3080));
   OAI221_X1 i_8_0_3141 (.A(n_8_0_6606), .B1(n_8_0_885), .B2(n_8_0_4587), 
      .C1(n_8_0_3935), .C2(n_8_0_5779), .ZN(n_8_0_3934));
   OAI221_X1 i_8_0_3149 (.A(n_8_0_6577), .B1(n_8_0_3924), .B2(n_8_0_884), 
      .C1(n_8_0_6325), .C2(n_8_0_5788), .ZN(n_8_0_3923));
   OAI211_X1 i_8_0_3153 (.A(n_8_0_6556), .B(n_8_0_3929), .C1(n_8_0_4542), 
      .C2(n_8_0_883), .ZN(n_8_0_3928));
   OAI21_X1 i_8_0_3154 (.A(n_8_0_3099), .B1(n_8_0_7221), .B2(n_8_0_3090), 
      .ZN(n_8_0_3081));
   INV_X1 i_8_0_3155 (.A(n_8_0_3098), .ZN(n_8_0_3090));
   NAND4_X1 i_8_0_3156 (.A1(n_8_0_3710), .A2(\out_bs[7] [5]), .A3(\out_bs[7] [3]), 
      .A4(n_8_0_6363), .ZN(n_8_0_3098));
   OAI21_X1 i_8_0_3159 (.A(n_8_0_880), .B1(n_8_0_6469), .B2(n_8_0_6361), 
      .ZN(n_8_0_3099));
   OR3_X1 i_8_0_3175 (.A1(n_8_0_3998), .A2(n_8_0_4016), .A3(n_8_0_3997), 
      .ZN(n_8_0_3100));
   OAI221_X1 i_8_0_3176 (.A(n_8_0_6577), .B1(n_8_0_860), .B2(n_8_0_4590), 
      .C1(n_8_0_3999), .C2(n_8_0_4592), .ZN(n_8_0_3998));
   AOI211_X1 i_8_0_3177 (.A(n_8_0_4014), .B(n_8_0_4107), .C1(n_8_0_858), 
      .C2(n_8_0_4104), .ZN(n_8_0_4013));
   INV_X1 i_8_0_3179 (.A(n_8_0_3115), .ZN(n_194));
   OAI21_X1 i_8_0_3186 (.A(n_8_0_3885), .B1(n_8_0_3140), .B2(n_8_0_3116), 
      .ZN(n_8_0_3115));
   OR3_X1 i_8_0_3187 (.A1(n_8_0_4043), .A2(n_8_0_4040), .A3(n_8_0_3117), 
      .ZN(n_8_0_3116));
   NAND3_X1 i_8_0_3188 (.A1(n_8_0_4025), .A2(n_8_0_4033), .A3(n_8_0_3123), 
      .ZN(n_8_0_3117));
   INV_X1 i_8_0_3192 (.A(n_8_0_3124), .ZN(n_8_0_3123));
   OR2_X1 i_8_0_3208 (.A1(n_8_0_4035), .A2(n_8_0_4038), .ZN(n_8_0_3124));
   OAI221_X1 i_8_0_3209 (.A(n_8_0_6526), .B1(n_8_0_6321), .B2(n_8_0_5901), 
      .C1(n_8_0_4036), .C2(n_8_0_854), .ZN(n_8_0_4035));
   AOI211_X1 i_8_0_3210 (.A(n_8_0_6607), .B(n_8_0_4034), .C1(n_8_0_5905), 
      .C2(n_8_0_4498), .ZN(n_8_0_4033));
   INV_X1 i_8_0_3212 (.A(n_8_0_3128), .ZN(n_8_0_4025));
   NAND2_X1 i_8_0_3216 (.A1(n_8_0_4026), .A2(n_8_0_4030), .ZN(n_8_0_3128));
   AOI211_X1 i_8_0_3254 (.A(n_8_0_4041), .B(n_8_0_4107), .C1(n_8_0_850), 
      .C2(n_8_0_4104), .ZN(n_8_0_4040));
   NAND2_X1 i_8_0_3255 (.A1(n_8_0_4044), .A2(n_8_0_6590), .ZN(n_8_0_4043));
   NAND2_X1 i_8_0_3256 (.A1(n_8_0_3175), .A2(n_8_0_3141), .ZN(n_8_0_3140));
   INV_X1 i_8_0_3257 (.A(n_8_0_3174), .ZN(n_8_0_3141));
   OAI21_X1 i_8_0_3258 (.A(n_8_0_6465), .B1(n_8_0_4595), .B2(n_8_0_848), 
      .ZN(n_8_0_3174));
   NAND3_X1 i_8_0_3270 (.A1(n_8_0_3176), .A2(n_8_0_4598), .A3(n_8_0_5914), 
      .ZN(n_8_0_3175));
   NAND2_X1 i_8_0_3281 (.A1(n_8_0_6469), .A2(n_8_0_848), .ZN(n_8_0_3176));
   INV_X1 i_8_0_3286 (.A(n_8_0_3205), .ZN(n_195));
   OAI21_X1 i_8_0_3292 (.A(n_8_0_3885), .B1(n_8_0_3214), .B2(n_8_0_3210), 
      .ZN(n_8_0_3205));
   OR3_X1 i_8_0_3297 (.A1(n_8_0_4063), .A2(n_8_0_4067), .A3(n_8_0_3212), 
      .ZN(n_8_0_3210));
   NAND2_X1 i_8_0_3298 (.A1(n_8_0_4056), .A2(n_8_0_3213), .ZN(n_8_0_3212));
   NOR4_X1 i_8_0_3299 (.A1(n_8_0_4053), .A2(n_8_0_6250), .A3(n_8_0_4049), 
      .A4(n_8_0_4065), .ZN(n_8_0_3213));
   OAI221_X1 i_8_0_3300 (.A(n_8_0_6606), .B1(n_8_0_6282), .B2(n_8_0_5947), 
      .C1(n_8_0_4066), .C2(n_8_0_845), .ZN(n_8_0_4065));
   AOI21_X1 i_8_0_3302 (.A(n_8_0_4054), .B1(n_8_0_844), .B2(n_8_0_6840), 
      .ZN(n_8_0_4053));
   AOI21_X1 i_8_0_3303 (.A(n_8_0_4061), .B1(n_8_0_4057), .B2(n_8_0_4060), 
      .ZN(n_8_0_4056));
   NAND2_X1 i_8_0_3304 (.A1(n_8_0_3239), .A2(n_8_0_3215), .ZN(n_8_0_3214));
   INV_X1 i_8_0_3305 (.A(n_8_0_3238), .ZN(n_8_0_3215));
   OAI21_X1 i_8_0_3310 (.A(n_8_0_6465), .B1(n_8_0_4595), .B2(n_8_0_840), 
      .ZN(n_8_0_3238));
   NAND3_X1 i_8_0_3320 (.A1(n_8_0_3242), .A2(n_8_0_4598), .A3(n_8_0_5952), 
      .ZN(n_8_0_3239));
   OAI21_X1 i_8_0_3324 (.A(n_8_0_6998), .B1(n_8_0_6997), .B2(n_8_0_6724), 
      .ZN(n_8_0_5952));
   NAND2_X1 i_8_0_3329 (.A1(n_8_0_6469), .A2(n_8_0_840), .ZN(n_8_0_3242));
   INV_X1 i_8_0_3333 (.A(n_8_0_3276), .ZN(n_196));
   OAI21_X1 i_8_0_3334 (.A(n_8_0_3885), .B1(n_8_0_3282), .B2(n_8_0_3277), 
      .ZN(n_8_0_3276));
   OR4_X1 i_8_0_3336 (.A1(n_8_0_4252), .A2(n_8_0_4250), .A3(n_8_0_4247), 
      .A4(n_8_0_3278), .ZN(n_8_0_3277));
   NAND3_X1 i_8_0_3337 (.A1(n_8_0_4272), .A2(n_8_0_4260), .A3(n_8_0_3279), 
      .ZN(n_8_0_3278));
   AOI211_X1 i_8_0_3339 (.A(n_8_0_4267), .B(n_8_0_4269), .C1(n_8_0_6185), 
      .C2(n_8_0_4268), .ZN(n_8_0_3279));
   NAND3_X1 i_8_0_3340 (.A1(n_8_0_4261), .A2(n_8_0_4263), .A3(n_8_0_4264), 
      .ZN(n_8_0_4260));
   INV_X1 i_8_0_3378 (.A(n_8_0_4273), .ZN(n_8_0_4272));
   OAI211_X1 i_8_0_3379 (.A(n_8_0_4248), .B(n_8_0_6556), .C1(n_8_0_6192), 
      .C2(n_8_0_4338), .ZN(n_8_0_4247));
   OAI221_X1 i_8_0_3380 (.A(n_8_0_6513), .B1(n_8_0_6211), .B2(n_8_0_4552), 
      .C1(n_8_0_4251), .C2(n_8_0_741), .ZN(n_8_0_4250));
   OAI211_X1 i_8_0_3381 (.A(n_8_0_4253), .B(n_8_0_6590), .C1(n_8_0_739), 
      .C2(n_8_0_4610), .ZN(n_8_0_4252));
   NAND3_X1 i_8_0_3382 (.A1(n_8_0_3309), .A2(n_8_0_3303), .A3(n_8_0_6465), 
      .ZN(n_8_0_3282));
   NAND2_X1 i_8_0_3383 (.A1(n_8_0_6468), .A2(n_8_0_6201), .ZN(n_8_0_3303));
   OAI21_X1 i_8_0_3385 (.A(n_8_0_3330), .B1(n_8_0_4596), .B2(n_8_0_3328), 
      .ZN(n_8_0_3309));
   INV_X1 i_8_0_3388 (.A(n_8_0_4259), .ZN(n_8_0_3328));
   INV_X1 i_8_0_3402 (.A(n_8_0_737), .ZN(n_8_0_3330));
   INV_X1 i_8_0_3404 (.A(n_8_0_3336), .ZN(n_197));
   OAI21_X1 i_8_0_3409 (.A(n_8_0_3885), .B1(n_8_0_3460), .B2(n_8_0_3337), 
      .ZN(n_8_0_3336));
   NAND4_X1 i_8_0_3410 (.A1(n_8_0_4298), .A2(n_8_0_4295), .A3(n_8_0_3377), 
      .A4(n_8_0_3354), .ZN(n_8_0_3337));
   INV_X1 i_8_0_3416 (.A(n_8_0_3355), .ZN(n_8_0_3354));
   OAI211_X1 i_8_0_3438 (.A(n_8_0_3375), .B(n_8_0_3357), .C1(n_8_0_4307), 
      .C2(n_8_0_6218), .ZN(n_8_0_3355));
   AOI21_X1 i_8_0_3439 (.A(n_8_0_4286), .B1(n_8_0_6253), .B2(n_8_0_4285), 
      .ZN(n_8_0_3357));
   AND2_X1 i_8_0_3441 (.A1(n_8_0_3376), .A2(n_8_0_6577), .ZN(n_8_0_3375));
   OR2_X1 i_8_0_3447 (.A1(n_8_0_4293), .A2(n_8_0_729), .ZN(n_8_0_3376));
   INV_X1 i_8_0_3448 (.A(n_8_0_4278), .ZN(n_8_0_3377));
   NAND3_X1 i_8_0_3465 (.A1(n_8_0_3474), .A2(n_8_0_3461), .A3(n_8_0_6465), 
      .ZN(n_8_0_3460));
   NAND2_X1 i_8_0_3467 (.A1(n_8_0_6468), .A2(n_8_0_6237), .ZN(n_8_0_3461));
   NAND2_X1 i_8_0_3468 (.A1(n_8_0_6997), .A2(n_8_0_6724), .ZN(n_8_0_6237));
   OAI21_X1 i_8_0_3469 (.A(n_8_0_3484), .B1(n_8_0_4596), .B2(n_8_0_3475), 
      .ZN(n_8_0_3474));
   AOI21_X1 i_8_0_3471 (.A(n_8_0_4532), .B1(n_8_0_6997), .B2(n_8_0_3476), 
      .ZN(n_8_0_3475));
   INV_X1 i_8_0_3480 (.A(n_8_0_6725), .ZN(n_8_0_3476));
   INV_X1 i_8_0_3487 (.A(n_8_0_4595), .ZN(n_8_0_4596));
   INV_X1 i_8_0_3490 (.A(n_8_0_721), .ZN(n_8_0_3484));
   INV_X1 i_8_0_3491 (.A(n_8_0_3544), .ZN(n_198));
   OAI21_X1 i_8_0_3492 (.A(n_8_0_3885), .B1(n_8_0_3602), .B2(n_8_0_3545), 
      .ZN(n_8_0_3544));
   NAND4_X1 i_8_0_3589 (.A1(n_8_0_4504), .A2(n_8_0_4481), .A3(n_8_0_4477), 
      .A4(n_8_0_3546), .ZN(n_8_0_3545));
   INV_X1 i_8_0_3590 (.A(n_8_0_3555), .ZN(n_8_0_3546));
   OAI211_X1 i_8_0_3591 (.A(n_8_0_4495), .B(n_8_0_3556), .C1(n_8_0_4511), 
      .C2(n_8_0_3569), .ZN(n_8_0_3555));
   NAND2_X1 i_8_0_3598 (.A1(n_8_0_6597), .A2(n_8_0_6520), .ZN(n_8_0_3556));
   NOR2_X1 i_8_0_3604 (.A1(n_8_0_6662), .A2(n_8_0_6523), .ZN(n_8_0_6520));
   NOR2_X1 i_8_0_3605 (.A1(n_8_0_6811), .A2(n_8_0_7084), .ZN(n_8_0_6597));
   OAI21_X1 i_8_0_3606 (.A(n_8_0_3581), .B1(n_8_0_3570), .B2(n_8_0_3573), 
      .ZN(n_8_0_3569));
   INV_X1 i_8_0_3607 (.A(n_8_0_4514), .ZN(n_8_0_3570));
   OAI21_X1 i_8_0_3608 (.A(n_8_0_7089), .B1(n_8_0_6817), .B2(\out_bs[0] [6]), 
      .ZN(n_8_0_4514));
   INV_X1 i_8_0_3615 (.A(n_8_0_6523), .ZN(n_8_0_3573));
   INV_X1 i_8_0_3686 (.A(n_8_0_575), .ZN(n_8_0_3581));
   INV_X1 i_8_0_3687 (.A(n_8_0_3582), .ZN(n_8_0_4504));
   NAND2_X1 i_8_0_3688 (.A1(n_8_0_3599), .A2(n_8_0_3600), .ZN(n_8_0_3582));
   NAND2_X1 i_8_0_3689 (.A1(n_8_0_4556), .A2(n_8_0_6549), .ZN(n_8_0_3599));
   INV_X1 i_8_0_3691 (.A(n_8_0_4505), .ZN(n_8_0_3600));
   NAND3_X1 i_8_0_3699 (.A1(n_8_0_3624), .A2(n_8_0_3603), .A3(n_8_0_6465), 
      .ZN(n_8_0_3602));
   NAND2_X1 i_8_0_3700 (.A1(n_8_0_6468), .A2(n_8_0_6541), .ZN(n_8_0_3603));
   INV_X1 i_8_0_3701 (.A(n_8_0_3604), .ZN(n_8_0_6541));
   NAND3_X1 i_8_0_3703 (.A1(\out_bs[7] [3]), .A2(\out_bs[7] [2]), .A3(n_8_0_3605), 
      .ZN(n_8_0_3604));
   INV_X1 i_8_0_3704 (.A(n_8_0_6544), .ZN(n_8_0_3605));
   NAND2_X1 i_8_0_3708 (.A1(n_8_0_3678), .A2(n_8_0_7221), .ZN(n_8_0_3624));
   AOI21_X1 i_8_0_3714 (.A(n_8_0_547), .B1(n_8_0_4595), .B2(n_8_0_6540), 
      .ZN(n_8_0_3678));
   AOI21_X1 i_8_0_3718 (.A(n_8_0_6853), .B1(n_8_0_4594), .B2(n_8_0_3679), 
      .ZN(n_199));
   NOR4_X1 i_8_0_3719 (.A1(n_8_0_4609), .A2(n_8_0_4570), .A3(n_8_0_4607), 
      .A4(n_8_0_3680), .ZN(n_8_0_3679));
   NAND3_X1 i_8_0_3720 (.A1(n_8_0_3698), .A2(n_8_0_4583), .A3(n_8_0_3690), 
      .ZN(n_8_0_3680));
   NOR2_X1 i_8_0_3723 (.A1(n_8_0_4578), .A2(n_8_0_4601), .ZN(n_8_0_3690));
   AOI21_X1 i_8_0_3724 (.A(n_8_0_4586), .B1(\out_bs[2] [5]), .B2(n_8_0_4584), 
      .ZN(n_8_0_4583));
   INV_X1 i_8_0_3728 (.A(n_8_0_4589), .ZN(n_8_0_3698));
   OAI211_X1 i_8_0_3731 (.A(n_8_0_6577), .B(n_8_0_4590), .C1(n_8_0_5466), 
      .C2(n_8_0_4592), .ZN(n_8_0_4589));
   INV_X1 i_8_0_3732 (.A(n_8_0_3708), .ZN(n_8_0_4594));
   NAND3_X1 i_8_0_3733 (.A1(n_8_0_3709), .A2(n_8_0_6465), .A3(n_8_0_4595), 
      .ZN(n_8_0_3708));
   NAND2_X1 i_8_0_3739 (.A1(n_8_0_4598), .A2(n_8_0_6719), .ZN(n_8_0_3709));
   NOR2_X1 i_8_0_3743 (.A1(n_8_0_6721), .A2(n_8_0_6722), .ZN(n_8_0_6719));
   NAND3_X1 i_8_0_3747 (.A1(n_8_0_7421), .A2(\out_as[7] [6]), .A3(n_8_0_3885), 
      .ZN(n_8_0_3710));
   AOI211_X1 i_8_0_3752 (.A(n_8_0_3751), .B(\out_bs[7] [0]), .C1(\out_bs[7] [1]), 
      .C2(n_8_0_3755), .ZN(n_8_0_3711));
   INV_X1 i_8_0_3753 (.A(\out_as[7] [0]), .ZN(n_8_0_3751));
   INV_X1 i_8_0_3754 (.A(\out_as[7] [1]), .ZN(n_8_0_3755));
   INV_X1 i_8_0_3755 (.A(\out_bs[7] [1]), .ZN(n_8_0_3756));
   AND3_X1 i_8_0_3756 (.A1(n_8_0_3853), .A2(n_8_0_3884), .A3(n_8_0_6465), 
      .ZN(n_8_0_4184));
   INV_X1 i_8_0_3757 (.A(in_data[4]), .ZN(n_8_0_6989));
   OAI21_X1 i_8_0_3759 (.A(n_8_0_3757), .B1(n_8_0_3819), .B2(n_8_0_7153), 
      .ZN(n_200));
   NAND3_X1 i_8_0_3760 (.A1(n_8_0_3811), .A2(n_8_0_3812), .A3(n_8_0_3758), 
      .ZN(n_8_0_3757));
   MUX2_X1 i_8_0_3772 (.A(n_8_0_3759), .B(in_data[4]), .S(n_8_0_3699), .Z(
      n_8_0_3758));
   NAND2_X1 i_8_0_3781 (.A1(n_8_0_3810), .A2(n_8_0_3762), .ZN(n_8_0_3759));
   NAND2_X1 i_8_0_3817 (.A1(n_8_0_3702), .A2(in_data[8]), .ZN(n_8_0_3762));
   OAI21_X1 i_8_0_3818 (.A(n_8_0_1738), .B1(n_8_0_1739), .B2(n_8_0_3721), 
      .ZN(n_8_0_3810));
   NAND2_X1 i_8_0_3819 (.A1(n_8_0_7155), .A2(n_8_0_7154), .ZN(n_8_0_3811));
   INV_X1 i_8_0_3838 (.A(n_8_0_4409), .ZN(n_8_0_3812));
   INV_X1 i_8_0_3839 (.A(in_data[0]), .ZN(n_8_0_3819));
   INV_X1 i_8_0_3840 (.A(n_8_0_3820), .ZN(n_201));
   NAND2_X1 i_8_0_3841 (.A1(n_8_0_3821), .A2(n_8_0_3885), .ZN(n_8_0_3820));
   NAND4_X1 i_8_0_3842 (.A1(n_8_0_3839), .A2(n_8_0_3884), .A3(n_8_0_6465), 
      .A4(n_8_0_4187), .ZN(n_8_0_3821));
   INV_X1 i_8_0_3843 (.A(n_8_0_3840), .ZN(n_8_0_3839));
   NAND4_X1 i_8_0_3848 (.A1(n_8_0_3853), .A2(n_8_0_3881), .A3(n_8_0_4178), 
      .A4(n_8_0_3866), .ZN(n_8_0_3840));
   NAND2_X1 i_8_0_3850 (.A1(n_8_0_3854), .A2(n_8_0_3863), .ZN(n_8_0_3853));
   NAND2_X1 i_8_0_3851 (.A1(n_8_0_4595), .A2(n_8_0_4186), .ZN(n_8_0_3854));
   INV_X1 i_8_0_3852 (.A(n_8_0_785), .ZN(n_8_0_3863));
   INV_X1 i_8_0_3853 (.A(n_8_0_3876), .ZN(n_8_0_3866));
   NAND2_X1 i_8_0_3855 (.A1(n_8_0_4181), .A2(n_8_0_3877), .ZN(n_8_0_3876));
   NOR2_X1 i_8_0_3859 (.A1(n_8_0_4165), .A2(n_8_0_4174), .ZN(n_8_0_3877));
   AOI21_X1 i_8_0_3860 (.A(n_8_0_4182), .B1(n_8_0_4308), .B2(n_8_0_5116), 
      .ZN(n_8_0_4181));
   AOI21_X1 i_8_0_3861 (.A(n_8_0_4179), .B1(n_8_0_4545), .B2(n_8_0_6092), 
      .ZN(n_8_0_4178));
   INV_X1 i_8_0_3864 (.A(n_8_0_4175), .ZN(n_8_0_3881));
   AOI21_X1 i_8_0_3867 (.A(n_8_0_4188), .B1(n_8_0_4611), .B2(n_8_0_6878), 
      .ZN(n_8_0_4187));
   NAND2_X1 i_8_0_3870 (.A1(n_8_0_7422), .A2(\out_as[7] [6]), .ZN(n_8_0_3882));
   NAND2_X1 i_8_0_3871 (.A1(n_8_0_6468), .A2(n_8_0_6080), .ZN(n_8_0_3884));
   INV_X1 i_8_0_3872 (.A(n_8_0_6853), .ZN(n_8_0_3885));
   INV_X1 i_8_0_3873 (.A(n_8_0_7222), .ZN(n_8_0_6404));
   NAND2_X1 i_8_0_3914 (.A1(\out_bs[7] [3]), .A2(n_8_0_6363), .ZN(n_8_0_6361));
   INV_X1 i_8_0_3915 (.A(n_8_0_7234), .ZN(n_8_0_6469));
   NAND2_X1 i_8_0_3916 (.A1(\out_bs[7] [4]), .A2(\out_bs[7] [3]), .ZN(n_8_0_6721));
   INV_X1 i_8_0_3919 (.A(n_8_0_7102), .ZN(n_8_0_6471));
   NAND2_X1 i_8_0_3920 (.A1(n_8_0_6729), .A2(n_8_0_3659), .ZN(n_8_0_3657));
   NAND2_X1 i_8_0_3921 (.A1(n_8_0_6998), .A2(n_8_0_6540), .ZN(n_8_0_5914));
   NAND2_X1 i_8_0_3922 (.A1(n_8_0_5358), .A2(n_8_0_6998), .ZN(n_8_0_5842));
   INV_X1 i_8_0_3923 (.A(n_8_0_7166), .ZN(n_8_0_5652));
   INV_X1 i_8_0_3926 (.A(n_8_0_4424), .ZN(n_8_0_4423));
   NAND3_X1 i_8_0_3975 (.A1(n_8_0_6728), .A2(\out_bs[7] [4]), .A3(\out_bs[7] [3]), 
      .ZN(n_8_0_6714));
   INV_X1 i_8_0_3976 (.A(n_8_0_7407), .ZN(n_8_0_6410));
   INV_X1 i_8_0_3977 (.A(n_8_0_7396), .ZN(n_8_0_6276));
   INV_X1 i_8_0_3978 (.A(n_8_0_7354), .ZN(n_8_0_5971));
   INV_X1 i_8_0_3985 (.A(n_8_0_7337), .ZN(n_8_0_5423));
   INV_X1 i_8_0_3986 (.A(n_8_0_7314), .ZN(n_8_0_5392));
   OAI21_X1 i_8_0_3987 (.A(n_8_0_7323), .B1(n_8_0_5406), .B2(n_8_0_344), 
      .ZN(n_8_0_5405));
   NAND2_X1 i_8_0_4001 (.A1(n_8_0_7305), .A2(n_8_0_5363), .ZN(n_8_0_5362));
   OAI21_X1 i_8_0_4005 (.A(n_8_0_5375), .B1(n_8_0_6837), .B2(n_8_0_217), 
      .ZN(n_8_0_5374));
   INV_X1 i_8_0_4006 (.A(n_8_0_7289), .ZN(n_8_0_5186));
   NAND2_X1 i_8_0_4007 (.A1(n_8_0_4376), .A2(n_8_0_7213), .ZN(n_8_0_4375));
   INV_X1 i_8_0_4020 (.A(n_8_0_4333), .ZN(n_8_0_4211));
   INV_X1 i_8_0_4021 (.A(n_8_0_4101), .ZN(n_8_0_4100));
   INV_X1 i_8_0_4022 (.A(n_8_0_7191), .ZN(n_8_0_4079));
   INV_X1 i_8_0_4030 (.A(n_8_0_7177), .ZN(n_8_0_3904));
   INV_X1 i_8_0_4033 (.A(n_8_0_7122), .ZN(n_8_0_3587));
   NAND2_X1 i_8_0_4034 (.A1(n_8_0_3593), .A2(n_8_0_7127), .ZN(n_8_0_3591));
   INV_X1 i_8_0_4044 (.A(n_8_0_7106), .ZN(n_8_0_3548));
   INV_X1 i_8_0_4045 (.A(n_8_0_7111), .ZN(n_8_0_3558));
   INV_X1 i_8_0_4046 (.A(n_8_0_3996), .ZN(n_8_0_3302));
   INV_X1 i_8_0_4049 (.A(n_8_0_6470), .ZN(n_8_0_3298));
   NAND2_X1 i_8_0_4050 (.A1(n_8_0_3201), .A2(n_8_0_6200), .ZN(n_8_0_3200));
   INV_X1 i_8_0_4051 (.A(n_8_0_5972), .ZN(n_8_0_3142));
   INV_X1 i_8_0_4052 (.A(n_8_0_5974), .ZN(n_8_0_3139));
   NAND2_X1 i_8_0_4053 (.A1(n_8_0_5412), .A2(n_8_0_5411), .ZN(n_8_0_3102));
   INV_X1 i_8_0_4054 (.A(n_8_0_5413), .ZN(n_8_0_3114));
   INV_X1 i_8_0_4055 (.A(n_8_0_5061), .ZN(n_8_0_3085));
   NAND2_X1 i_8_0_4057 (.A1(n_8_0_5172), .A2(n_8_0_5171), .ZN(n_8_0_3095));
   INV_X1 i_8_0_4060 (.A(n_8_0_4567), .ZN(n_8_0_2753));
   OAI21_X1 i_8_0_4061 (.A(n_8_0_3886), .B1(n_8_0_6988), .B2(n_8_0_2979), 
      .ZN(n_202));
   NAND2_X1 i_8_0_4062 (.A1(n_8_0_2979), .A2(n_8_0_3892), .ZN(n_8_0_3886));
   OAI21_X1 i_8_0_4064 (.A(n_8_0_1485), .B1(n_8_0_6989), .B2(n_8_0_2964), 
      .ZN(n_8_0_3892));
   AOI21_X1 i_8_0_4068 (.A(n_8_0_3903), .B1(n_8_0_6729), .B2(n_8_0_2982), 
      .ZN(n_8_0_2979));
   AOI22_X1 i_8_0_4072 (.A1(n_8_0_6730), .A2(n_8_0_2981), .B1(n_8_0_6279), 
      .B2(n_8_0_3244), .ZN(n_8_0_3903));
   MUX2_X1 i_8_0_4073 (.A(in_data[0]), .B(n_8_0_3905), .S(n_8_0_5174), .Z(n_203));
   INV_X1 i_8_0_4074 (.A(n_8_0_3906), .ZN(n_8_0_3905));
   OAI21_X1 i_8_0_4075 (.A(n_8_0_3907), .B1(n_8_0_4047), .B2(n_8_0_5173), 
      .ZN(n_8_0_3906));
   OAI211_X1 i_8_0_4076 (.A(n_8_0_5173), .B(n_8_0_1530), .C1(n_8_0_6990), 
      .C2(n_8_0_3087), .ZN(n_8_0_3907));
   OAI21_X1 i_8_0_4086 (.A(n_8_0_3917), .B1(n_8_0_6720), .B2(n_8_0_3918), 
      .ZN(n_204));
   NAND2_X1 i_8_0_4087 (.A1(n_8_0_6720), .A2(in_data[0]), .ZN(n_8_0_3917));
   AOI22_X1 i_8_0_4088 (.A1(n_8_0_1591), .A2(n_8_0_3919), .B1(in_data[4]), 
      .B2(n_8_0_3285), .ZN(n_8_0_3918));
   OAI21_X1 i_8_0_4089 (.A(n_8_0_3286), .B1(n_8_0_786), .B2(n_8_0_3287), 
      .ZN(n_8_0_3285));
   OR2_X1 i_8_0_4093 (.A1(n_8_0_3296), .A2(n_8_0_1592), .ZN(n_8_0_3919));
   OAI21_X1 i_8_0_4098 (.A(n_8_0_3940), .B1(n_8_0_6988), .B2(n_8_0_3996), 
      .ZN(n_205));
   NAND2_X1 i_8_0_4104 (.A1(n_8_0_3996), .A2(n_8_0_3941), .ZN(n_8_0_3940));
   OAI21_X1 i_8_0_4109 (.A(n_8_0_3995), .B1(n_8_0_4408), .B2(n_8_0_3310), 
      .ZN(n_8_0_3941));
   OAI211_X1 i_8_0_4110 (.A(n_8_0_3310), .B(n_8_0_1601), .C1(in_data[8]), 
      .C2(n_8_0_3306), .ZN(n_8_0_3995));
   NOR2_X1 i_8_0_4111 (.A1(n_8_0_4003), .A2(n_8_0_4002), .ZN(n_8_0_3996));
   OAI21_X1 i_8_0_4167 (.A(n_8_0_4422), .B1(n_8_0_3478), .B2(n_8_0_768), 
      .ZN(n_8_0_4002));
   INV_X1 i_8_0_4168 (.A(n_8_0_4020), .ZN(n_8_0_4003));
   NAND2_X1 i_8_0_4169 (.A1(n_8_0_3304), .A2(n_8_0_6118), .ZN(n_8_0_4020));
   INV_X1 i_8_0_4171 (.A(n_8_0_4021), .ZN(n_206));
   OAI21_X1 i_8_0_4174 (.A(n_8_0_4023), .B1(n_8_0_6736), .B2(in_data[0]), 
      .ZN(n_8_0_4021));
   NAND3_X1 i_8_0_4175 (.A1(n_8_0_4051), .A2(n_8_0_4048), .A3(n_8_0_4024), 
      .ZN(n_8_0_4023));
   OAI21_X1 i_8_0_4176 (.A(n_8_0_4037), .B1(n_8_0_4047), .B2(n_8_0_4046), 
      .ZN(n_8_0_4024));
   NAND2_X1 i_8_0_4186 (.A1(n_8_0_1610), .A2(n_8_0_1608), .ZN(n_8_0_4037));
   INV_X1 i_8_0_4193 (.A(n_8_0_3346), .ZN(n_8_0_4046));
   INV_X1 i_8_0_4194 (.A(n_8_0_6989), .ZN(n_8_0_4047));
   INV_X1 i_8_0_4195 (.A(n_8_0_6737), .ZN(n_8_0_4048));
   NAND2_X1 i_8_0_4196 (.A1(n_8_0_3338), .A2(n_8_0_6738), .ZN(n_8_0_4051));
   INV_X1 i_8_0_4197 (.A(n_8_0_4052), .ZN(n_207));
   OAI21_X1 i_8_0_4198 (.A(n_8_0_4075), .B1(n_8_0_6872), .B2(n_8_0_4076), 
      .ZN(n_8_0_4052));
   NAND2_X1 i_8_0_4199 (.A1(n_8_0_6872), .A2(n_8_0_6988), .ZN(n_8_0_4075));
   AOI21_X1 i_8_0_4207 (.A(n_8_0_4077), .B1(n_8_0_4081), .B2(n_8_0_4080), 
      .ZN(n_8_0_4076));
   NOR2_X1 i_8_0_4209 (.A1(n_8_0_3365), .A2(in_data[4]), .ZN(n_8_0_4077));
   NAND2_X1 i_8_0_4211 (.A1(n_8_0_3372), .A2(n_8_0_1619), .ZN(n_8_0_4080));
   INV_X1 i_8_0_4214 (.A(n_8_0_1618), .ZN(n_8_0_4081));
   INV_X1 i_8_0_4217 (.A(n_8_0_4116), .ZN(n_208));
   OAI21_X1 i_8_0_4220 (.A(n_8_0_4136), .B1(n_8_0_7097), .B2(n_8_0_4137), 
      .ZN(n_8_0_4116));
   NAND2_X1 i_8_0_4221 (.A1(n_8_0_7097), .A2(n_8_0_6988), .ZN(n_8_0_4136));
   MUX2_X1 i_8_0_4222 (.A(n_8_0_4156), .B(in_data[4]), .S(n_8_0_7095), .Z(
      n_8_0_4137));
   INV_X1 i_8_0_4223 (.A(n_8_0_1658), .ZN(n_8_0_4156));
   AOI21_X1 i_8_0_4225 (.A(n_8_0_4160), .B1(n_8_0_4164), .B2(n_8_0_4161), 
      .ZN(n_209));
   NOR2_X1 i_8_0_4226 (.A1(n_8_0_4164), .A2(in_data[0]), .ZN(n_8_0_4160));
   OAI21_X1 i_8_0_4227 (.A(n_8_0_4162), .B1(in_data[4]), .B2(n_8_0_3813), 
      .ZN(n_8_0_4161));
   NAND2_X1 i_8_0_4228 (.A1(n_8_0_3813), .A2(n_8_0_4163), .ZN(n_8_0_4162));
   INV_X1 i_8_0_4231 (.A(n_8_0_1775), .ZN(n_8_0_4163));
   INV_X1 i_8_0_4240 (.A(n_8_0_7163), .ZN(n_8_0_4164));
   OAI21_X1 i_8_0_4250 (.A(n_8_0_4185), .B1(n_8_0_7172), .B2(n_8_0_4190), 
      .ZN(n_210));
   NAND2_X1 i_8_0_4251 (.A1(n_8_0_7172), .A2(in_data[0]), .ZN(n_8_0_4185));
   AOI21_X1 i_8_0_4252 (.A(n_8_0_4206), .B1(n_8_0_4246), .B2(n_8_0_4207), 
      .ZN(n_8_0_4190));
   NOR2_X1 i_8_0_4253 (.A1(n_8_0_4246), .A2(n_8_0_4408), .ZN(n_8_0_4206));
   AOI22_X1 i_8_0_4255 (.A1(n_8_0_1784), .A2(n_8_0_1785), .B1(n_8_0_6990), 
      .B2(n_8_0_3855), .ZN(n_8_0_4207));
   INV_X1 i_8_0_4256 (.A(n_8_0_7171), .ZN(n_8_0_4246));
   OAI21_X1 i_8_0_4257 (.A(n_8_0_4256), .B1(n_8_0_6988), .B2(n_8_0_4115), 
      .ZN(n_211));
   NAND2_X1 i_8_0_4259 (.A1(n_8_0_4115), .A2(n_8_0_4258), .ZN(n_8_0_4256));
   OAI22_X1 i_8_0_4266 (.A1(n_8_0_1874), .A2(n_8_0_1882), .B1(n_8_0_6989), 
      .B2(n_8_0_4117), .ZN(n_8_0_4258));
   INV_X1 i_8_0_4272 (.A(n_8_0_4266), .ZN(n_8_0_4115));
   OAI211_X1 i_8_0_4276 (.A(n_8_0_6467), .B(n_8_0_6465), .C1(n_8_0_4503), 
      .C2(n_8_0_817), .ZN(n_8_0_4266));
   INV_X1 i_8_0_4292 (.A(n_8_0_4275), .ZN(n_212));
   OAI21_X1 i_8_0_4293 (.A(n_8_0_4276), .B1(in_data[0]), .B2(n_8_0_7197), 
      .ZN(n_8_0_4275));
   NAND2_X1 i_8_0_4313 (.A1(n_8_0_7197), .A2(n_8_0_4277), .ZN(n_8_0_4276));
   OAI21_X1 i_8_0_4314 (.A(n_8_0_4291), .B1(in_data[4]), .B2(n_8_0_7196), 
      .ZN(n_8_0_4277));
   NAND2_X1 i_8_0_4315 (.A1(n_8_0_7196), .A2(n_8_0_4294), .ZN(n_8_0_4291));
   AOI21_X1 i_8_0_4334 (.A(n_8_0_1885), .B1(in_data[8]), .B2(n_8_0_4150), 
      .ZN(n_8_0_4294));
   INV_X1 i_8_0_4338 (.A(n_8_0_4301), .ZN(n_213));
   OAI21_X1 i_8_0_4339 (.A(n_8_0_4302), .B1(n_8_0_7205), .B2(n_8_0_4318), 
      .ZN(n_8_0_4301));
   NAND2_X1 i_8_0_4340 (.A1(n_8_0_7205), .A2(n_8_0_6988), .ZN(n_8_0_4302));
   MUX2_X1 i_8_0_4341 (.A(n_8_0_4332), .B(in_data[4]), .S(n_8_0_4333), .Z(
      n_8_0_4318));
   OAI21_X1 i_8_0_4342 (.A(n_8_0_1906), .B1(n_8_0_1907), .B2(n_8_0_4204), 
      .ZN(n_8_0_4332));
   OAI21_X1 i_8_0_4343 (.A(n_8_0_4355), .B1(n_8_0_4356), .B2(n_8_0_4334), 
      .ZN(n_8_0_4333));
   INV_X1 i_8_0_4357 (.A(n_8_0_4213), .ZN(n_8_0_4334));
   INV_X1 i_8_0_4360 (.A(n_8_0_4212), .ZN(n_8_0_4355));
   INV_X1 i_8_0_4363 (.A(n_8_0_4559), .ZN(n_8_0_4356));
   INV_X1 i_8_0_4364 (.A(n_8_0_4371), .ZN(n_214));
   OAI21_X1 i_8_0_4366 (.A(n_8_0_4372), .B1(n_8_0_7218), .B2(n_8_0_4379), 
      .ZN(n_8_0_4371));
   NAND2_X1 i_8_0_4369 (.A1(n_8_0_7218), .A2(n_8_0_6988), .ZN(n_8_0_4372));
   INV_X1 i_8_0_4370 (.A(n_8_0_4388), .ZN(n_8_0_4379));
   MUX2_X1 i_8_0_4386 (.A(n_8_0_4404), .B(n_8_0_4408), .S(n_8_0_4405), .Z(
      n_8_0_4388));
   AOI21_X1 i_8_0_4387 (.A(n_8_0_1974), .B1(in_data[8]), .B2(n_8_0_4401), 
      .ZN(n_8_0_4404));
   INV_X1 i_8_0_4391 (.A(in_data[4]), .ZN(n_8_0_4408));
   AOI21_X1 i_8_0_4427 (.A(n_8_0_4410), .B1(n_8_0_4469), .B2(n_8_0_7350), 
      .ZN(n_215));
   NOR2_X1 i_8_0_4428 (.A1(n_8_0_7350), .A2(n_8_0_4444), .ZN(n_8_0_4410));
   OAI21_X1 i_8_0_4429 (.A(n_8_0_4459), .B1(n_8_0_6990), .B2(n_8_0_7349), 
      .ZN(n_8_0_4444));
   NAND2_X1 i_8_0_4432 (.A1(n_8_0_7349), .A2(n_8_0_4460), .ZN(n_8_0_4459));
   AOI22_X1 i_8_0_4434 (.A1(n_8_0_2546), .A2(n_8_0_2547), .B1(n_8_0_6991), 
      .B2(n_8_0_5993), .ZN(n_8_0_4460));
   NAND2_X1 i_8_0_4438 (.A1(n_8_0_2543), .A2(n_8_0_4470), .ZN(n_8_0_4469));
   NAND2_X1 i_8_0_4439 (.A1(n_8_0_7354), .A2(n_8_0_6988), .ZN(n_8_0_4470));
   INV_X1 i_8_0_4440 (.A(in_data[0]), .ZN(n_8_0_6988));
   AOI21_X1 i_8_0_4442 (.A(n_8_0_6853), .B1(n_8_0_4567), .B2(n_8_0_4474), 
      .ZN(n_216));
   INV_X1 i_8_0_4448 (.A(n_8_0_4475), .ZN(n_8_0_4474));
   NAND2_X1 i_8_0_4454 (.A1(n_8_0_2738), .A2(n_8_0_4476), .ZN(n_8_0_4475));
   NOR2_X1 i_8_0_4457 (.A1(n_8_0_2765), .A2(n_8_0_4500), .ZN(n_8_0_4476));
   NAND3_X1 i_8_0_4458 (.A1(n_8_0_2745), .A2(n_8_0_2741), .A3(n_8_0_4502), 
      .ZN(n_8_0_4500));
   NOR3_X1 i_8_0_4459 (.A1(n_8_0_2758), .A2(n_8_0_4566), .A3(n_8_0_2761), 
      .ZN(n_8_0_4502));
   OAI211_X1 i_8_0_4460 (.A(n_8_0_4231), .B(n_8_0_2762), .C1(n_8_0_6782), 
      .C2(n_8_0_5526), .ZN(n_8_0_2761));
   AOI21_X1 i_8_0_4473 (.A(n_8_0_2759), .B1(n_8_0_4127), .B2(n_8_0_5515), 
      .ZN(n_8_0_2758));
   INV_X1 i_8_0_4474 (.A(n_8_0_2749), .ZN(n_8_0_4566));
   AOI22_X1 i_8_0_4475 (.A1(n_8_0_6824), .A2(n_8_0_2768), .B1(n_8_0_2766), 
      .B2(n_8_0_5518), .ZN(n_8_0_2765));
   OAI21_X1 i_8_0_4477 (.A(n_8_0_4613), .B1(n_8_0_4569), .B2(n_8_0_4568), 
      .ZN(n_8_0_4567));
   NAND2_X1 i_8_0_4484 (.A1(n_8_0_3244), .A2(n_8_0_6041), .ZN(n_8_0_4568));
   NOR2_X1 i_8_0_4485 (.A1(n_8_0_6730), .A2(n_8_0_4614), .ZN(n_8_0_4569));
   NAND2_X1 i_8_0_4486 (.A1(n_8_0_6730), .A2(n_8_0_4614), .ZN(n_8_0_4613));
   NAND2_X1 i_8_0_4487 (.A1(n_8_0_2982), .A2(n_8_0_2757), .ZN(n_8_0_4614));
   INV_X1 i_8_0_4496 (.A(n_8_0_4615), .ZN(n_8_0_2982));
   OR2_X1 i_8_0_4498 (.A1(n_8_0_3658), .A2(n_8_0_1296), .ZN(n_8_0_4615));
   INV_X1 i_8_0_4502 (.A(n_8_0_4616), .ZN(n_217));
   OAI21_X1 i_8_0_4512 (.A(n_8_0_6854), .B1(n_8_0_4846), .B2(n_8_0_4814), 
      .ZN(n_8_0_4616));
   NAND3_X1 i_8_0_4514 (.A1(n_8_0_2924), .A2(n_8_0_2928), .A3(n_8_0_4815), 
      .ZN(n_8_0_4814));
   INV_X1 i_8_0_4516 (.A(n_8_0_4821), .ZN(n_8_0_4815));
   NAND3_X1 i_8_0_4517 (.A1(n_8_0_2921), .A2(n_8_0_2947), .A3(n_8_0_4822), 
      .ZN(n_8_0_4821));
   INV_X1 i_8_0_4518 (.A(n_8_0_4830), .ZN(n_8_0_4822));
   OR2_X1 i_8_0_4540 (.A1(n_8_0_2939), .A2(n_8_0_4844), .ZN(n_8_0_4830));
   NAND3_X1 i_8_0_4541 (.A1(n_8_0_2935), .A2(n_8_0_2933), .A3(n_8_0_4845), 
      .ZN(n_8_0_4844));
   OAI21_X1 i_8_0_4542 (.A(n_8_0_6810), .B1(n_8_0_3015), .B2(n_8_0_6668), 
      .ZN(n_8_0_4845));
   OAI22_X1 i_8_0_4549 (.A1(n_8_0_6781), .A2(n_8_0_2937), .B1(n_8_0_2936), 
      .B2(n_8_0_5668), .ZN(n_8_0_2935));
   OAI21_X1 i_8_0_4556 (.A(n_8_0_2940), .B1(n_8_0_6772), .B2(n_8_0_2941), 
      .ZN(n_8_0_2939));
   OAI21_X1 i_8_0_4557 (.A(n_8_0_2929), .B1(n_8_0_2930), .B2(n_8_0_6300), 
      .ZN(n_8_0_2928));
   INV_X1 i_8_0_4558 (.A(n_8_0_2943), .ZN(n_8_0_4846));
   OAI21_X1 i_8_0_4561 (.A(n_8_0_4847), .B1(n_8_0_5674), .B2(n_8_0_3691), 
      .ZN(n_8_0_2943));
   OAI21_X1 i_8_0_4565 (.A(n_8_0_2945), .B1(n_8_0_505), .B2(n_8_0_2981), 
      .ZN(n_8_0_4847));
   NAND2_X1 i_8_0_4574 (.A1(n_8_0_3659), .A2(n_8_0_2983), .ZN(n_8_0_2981));
   AOI21_X1 i_8_0_4575 (.A(n_8_0_6853), .B1(n_8_0_5174), .B2(n_8_0_4849), 
      .ZN(n_218));
   INV_X1 i_8_0_4591 (.A(n_8_0_4850), .ZN(n_8_0_4849));
   NAND4_X1 i_8_0_4595 (.A1(n_8_0_5173), .A2(n_8_0_3087), .A3(n_8_0_3093), 
      .A4(n_8_0_5059), .ZN(n_8_0_4850));
   INV_X1 i_8_0_4596 (.A(n_8_0_5060), .ZN(n_8_0_5059));
   NAND4_X1 i_8_0_4597 (.A1(n_8_0_5172), .A2(n_8_0_3076), .A3(n_8_0_5171), 
      .A4(n_8_0_5061), .ZN(n_8_0_5060));
   OAI221_X1 i_8_0_4610 (.A(n_8_0_5064), .B1(n_8_0_5068), .B2(n_8_0_7370), 
      .C1(n_8_0_5063), .C2(n_8_0_5062), .ZN(n_8_0_5061));
   INV_X1 i_8_0_4611 (.A(n_8_0_5846), .ZN(n_8_0_5062));
   INV_X1 i_8_0_4612 (.A(n_8_0_3086), .ZN(n_8_0_5063));
   INV_X1 i_8_0_4632 (.A(n_8_0_3639), .ZN(n_8_0_5064));
   INV_X1 i_8_0_4633 (.A(n_8_0_1326), .ZN(n_8_0_5068));
   INV_X1 i_8_0_4648 (.A(n_8_0_3096), .ZN(n_8_0_5171));
   INV_X1 i_8_0_4649 (.A(n_8_0_3097), .ZN(n_8_0_5172));
   AOI21_X1 i_8_0_4654 (.A(n_8_0_3091), .B1(n_8_0_3647), .B2(n_8_0_3092), 
      .ZN(n_8_0_5173));
   OAI21_X1 i_8_0_4657 (.A(n_8_0_5175), .B1(n_8_0_6729), .B2(n_8_0_5357), 
      .ZN(n_8_0_5174));
   OAI22_X1 i_8_0_4658 (.A1(n_8_0_6730), .A2(n_8_0_5356), .B1(n_8_0_608), 
      .B2(n_8_0_3211), .ZN(n_8_0_5175));
   INV_X1 i_8_0_4659 (.A(n_8_0_5357), .ZN(n_8_0_5356));
   NAND3_X1 i_8_0_4660 (.A1(n_8_0_4424), .A2(n_8_0_6998), .A3(n_8_0_5358), 
      .ZN(n_8_0_5357));
   INV_X1 i_8_0_4663 (.A(n_8_0_6474), .ZN(n_8_0_5358));
   AOI21_X1 i_8_0_4664 (.A(n_8_0_6853), .B1(n_8_0_5413), .B2(n_8_0_5359), 
      .ZN(n_219));
   INV_X1 i_8_0_4665 (.A(n_8_0_5361), .ZN(n_8_0_5359));
   NAND4_X1 i_8_0_4666 (.A1(n_8_0_5412), .A2(n_8_0_3121), .A3(n_8_0_5411), 
      .A4(n_8_0_5380), .ZN(n_8_0_5361));
   INV_X1 i_8_0_4690 (.A(n_8_0_5381), .ZN(n_8_0_5380));
   NAND4_X1 i_8_0_4691 (.A1(n_8_0_3105), .A2(n_8_0_3118), .A3(n_8_0_3111), 
      .A4(n_8_0_5391), .ZN(n_8_0_5381));
   INV_X1 i_8_0_4692 (.A(n_8_0_5401), .ZN(n_8_0_5391));
   OAI211_X1 i_8_0_4693 (.A(n_8_0_3108), .B(n_8_0_5402), .C1(n_8_0_605), 
      .C2(n_8_0_3101), .ZN(n_8_0_5401));
   NAND2_X1 i_8_0_4694 (.A1(n_8_0_7393), .A2(n_8_0_5410), .ZN(n_8_0_5402));
   NAND2_X1 i_8_0_4705 (.A1(n_8_0_4604), .A2(n_8_0_5941), .ZN(n_8_0_5410));
   INV_X1 i_8_0_4722 (.A(n_8_0_3103), .ZN(n_8_0_5411));
   INV_X1 i_8_0_4723 (.A(n_8_0_3104), .ZN(n_8_0_5412));
   OAI22_X1 i_8_0_4757 (.A1(n_8_0_5962), .A2(n_8_0_5437), .B1(n_8_0_3691), 
      .B2(n_8_0_7184), .ZN(n_8_0_5413));
   AOI21_X1 i_8_0_4758 (.A(n_8_0_6730), .B1(n_8_0_5954), .B2(n_8_0_4424), 
      .ZN(n_8_0_5437));
   INV_X1 i_8_0_4759 (.A(n_8_0_5963), .ZN(n_8_0_5962));
   NAND2_X1 i_8_0_4760 (.A1(n_8_0_6238), .A2(n_8_0_6859), .ZN(n_8_0_5963));
   INV_X1 i_8_0_4761 (.A(n_8_0_577), .ZN(n_8_0_6859));
   AOI21_X1 i_8_0_4775 (.A(n_8_0_6853), .B1(n_8_0_5974), .B2(n_8_0_5964), 
      .ZN(n_220));
   INV_X1 i_8_0_4781 (.A(n_8_0_5967), .ZN(n_8_0_5964));
   NAND4_X1 i_8_0_4786 (.A1(n_8_0_3131), .A2(n_8_0_3129), .A3(n_8_0_3145), 
      .A4(n_8_0_5968), .ZN(n_8_0_5967));
   AND3_X1 i_8_0_4787 (.A1(n_8_0_5972), .A2(n_8_0_3137), .A3(n_8_0_3125), 
      .ZN(n_8_0_5968));
   NAND2_X1 i_8_0_4788 (.A1(n_8_0_3144), .A2(n_8_0_3143), .ZN(n_8_0_5972));
   OAI211_X1 i_8_0_4789 (.A(n_8_0_3146), .B(n_8_0_3184), .C1(n_8_0_3183), 
      .C2(n_8_0_6516), .ZN(n_8_0_3145));
   OAI21_X1 i_8_0_4790 (.A(n_8_0_6104), .B1(n_8_0_6103), .B2(n_8_0_6102), 
      .ZN(n_8_0_5974));
   OAI22_X1 i_8_0_4791 (.A1(n_8_0_6730), .A2(n_8_0_3244), .B1(n_8_0_545), 
      .B2(n_8_0_3211), .ZN(n_8_0_6102));
   AND2_X1 i_8_0_4792 (.A1(n_8_0_6729), .A2(n_8_0_6541), .ZN(n_8_0_6103));
   NAND3_X1 i_8_0_4805 (.A1(n_8_0_3692), .A2(n_8_0_6998), .A3(n_8_0_6540), 
      .ZN(n_8_0_6104));
   AOI21_X1 i_8_0_4806 (.A(n_8_0_6853), .B1(n_8_0_3209), .B2(n_8_0_6116), 
      .ZN(n_221));
   AOI21_X1 i_8_0_4807 (.A(n_8_0_6119), .B1(n_8_0_3201), .B2(n_8_0_6200), 
      .ZN(n_8_0_6116));
   NAND4_X1 i_8_0_4808 (.A1(n_8_0_3182), .A2(n_8_0_3196), .A3(n_8_0_3177), 
      .A4(n_8_0_6137), .ZN(n_8_0_6119));
   AOI211_X1 i_8_0_4809 (.A(n_8_0_6178), .B(n_8_0_3187), .C1(n_8_0_6177), 
      .C2(n_8_0_6176), .ZN(n_8_0_6137));
   OAI211_X1 i_8_0_4810 (.A(n_8_0_4604), .B(n_8_0_6000), .C1(n_8_0_6816), 
      .C2(n_8_0_3206), .ZN(n_8_0_6176));
   NAND2_X1 i_8_0_4811 (.A1(n_8_0_6811), .A2(n_8_0_3206), .ZN(n_8_0_6177));
   AOI21_X1 i_8_0_4812 (.A(n_8_0_3188), .B1(n_8_0_6772), .B2(n_8_0_3190), 
      .ZN(n_8_0_3187));
   INV_X1 i_8_0_4816 (.A(n_8_0_3192), .ZN(n_8_0_6178));
   OAI21_X1 i_8_0_4817 (.A(n_8_0_3178), .B1(n_8_0_6838), .B2(n_8_0_3181), 
      .ZN(n_8_0_3177));
   NAND2_X1 i_8_0_4818 (.A1(n_8_0_3197), .A2(n_8_0_3198), .ZN(n_8_0_3196));
   OR2_X1 i_8_0_5014 (.A1(n_8_0_3202), .A2(n_8_0_5969), .ZN(n_8_0_6200));
   AOI21_X1 i_8_0_5015 (.A(n_8_0_6202), .B1(n_8_0_6729), .B2(n_8_0_6238), 
      .ZN(n_8_0_3209));
   AOI22_X1 i_8_0_5016 (.A1(n_8_0_6730), .A2(n_8_0_3211), .B1(n_8_0_7359), 
      .B2(n_8_0_4424), .ZN(n_8_0_6202));
   INV_X1 i_8_0_5017 (.A(n_8_0_3211), .ZN(n_8_0_6238));
   NAND2_X1 i_8_0_5021 (.A1(n_8_0_3659), .A2(n_8_0_7004), .ZN(n_8_0_3211));
   AOI21_X1 i_8_0_5022 (.A(n_8_0_6853), .B1(n_8_0_3241), .B2(n_8_0_6257), 
      .ZN(n_222));
   INV_X1 i_8_0_5023 (.A(n_8_0_6258), .ZN(n_8_0_6257));
   OR3_X1 i_8_0_5024 (.A1(n_8_0_3235), .A2(n_8_0_3224), .A3(n_8_0_6259), 
      .ZN(n_8_0_6258));
   NAND4_X1 i_8_0_5025 (.A1(n_8_0_3219), .A2(n_8_0_3228), .A3(n_8_0_3231), 
      .A4(n_8_0_6260), .ZN(n_8_0_6259));
   NOR3_X1 i_8_0_5028 (.A1(n_8_0_3216), .A2(n_8_0_6377), .A3(n_8_0_6277), 
      .ZN(n_8_0_6260));
   AOI211_X1 i_8_0_5031 (.A(n_8_0_830), .B(n_8_0_3643), .C1(n_8_0_6816), 
      .C2(n_8_0_3240), .ZN(n_8_0_6277));
   NOR2_X1 i_8_0_5045 (.A1(n_8_0_6811), .A2(n_8_0_3240), .ZN(n_8_0_6377));
   AOI21_X1 i_8_0_5046 (.A(n_8_0_3234), .B1(n_8_0_3233), .B2(n_8_0_3232), 
      .ZN(n_8_0_3231));
   OAI21_X1 i_8_0_5047 (.A(n_8_0_3230), .B1(\out_bs[3] [4]), .B2(n_8_0_3229), 
      .ZN(n_8_0_3228));
   OAI21_X1 i_8_0_5048 (.A(n_8_0_3221), .B1(n_8_0_4059), .B2(n_8_0_3220), 
      .ZN(n_8_0_3219));
   OAI22_X1 i_8_0_5049 (.A1(n_8_0_3236), .A2(n_8_0_818), .B1(n_8_0_3237), 
      .B2(n_8_0_6755), .ZN(n_8_0_3235));
   AOI21_X1 i_8_0_5050 (.A(n_8_0_6388), .B1(n_8_0_6729), .B2(n_8_0_3243), 
      .ZN(n_8_0_3241));
   AOI211_X1 i_8_0_5051 (.A(n_8_0_816), .B(n_8_0_3658), .C1(n_8_0_6730), 
      .C2(n_8_0_3244), .ZN(n_8_0_6388));
   INV_X1 i_8_0_5052 (.A(n_8_0_3243), .ZN(n_8_0_3244));
   NAND2_X1 i_8_0_5053 (.A1(n_8_0_4424), .A2(n_8_0_6998), .ZN(n_8_0_3243));
   INV_X1 i_8_0_5063 (.A(n_8_0_6402), .ZN(n_223));
   OAI21_X1 i_8_0_5066 (.A(n_8_0_6854), .B1(n_8_0_6720), .B2(n_8_0_6415), 
      .ZN(n_8_0_6402));
   OR4_X1 i_8_0_5069 (.A1(n_8_0_6616), .A2(n_8_0_3296), .A3(n_8_0_3280), 
      .A4(n_8_0_6470), .ZN(n_8_0_6415));
   OAI21_X1 i_8_0_5265 (.A(n_8_0_6567), .B1(n_8_0_6568), .B2(n_8_0_6615), 
      .ZN(n_8_0_6470));
   INV_X1 i_8_0_5268 (.A(n_8_0_3299), .ZN(n_8_0_6567));
   INV_X1 i_8_0_5269 (.A(n_8_0_6623), .ZN(n_8_0_6568));
   INV_X1 i_8_0_5270 (.A(n_8_0_6092), .ZN(n_8_0_6615));
   OAI221_X1 i_8_0_5271 (.A(n_8_0_3683), .B1(n_8_0_792), .B2(n_8_0_3281), 
      .C1(n_8_0_4309), .C2(n_8_0_5115), .ZN(n_8_0_3280));
   OAI221_X1 i_8_0_5272 (.A(n_8_0_3803), .B1(n_8_0_6098), .B2(n_8_0_3623), 
      .C1(n_8_0_3297), .C2(n_8_0_788), .ZN(n_8_0_3296));
   INV_X1 i_8_0_5273 (.A(n_8_0_3283), .ZN(n_8_0_6616));
   OAI211_X1 i_8_0_5274 (.A(n_8_0_6732), .B(n_8_0_4422), .C1(n_8_0_784), 
      .C2(n_8_0_3478), .ZN(n_8_0_6720));
   OAI21_X1 i_8_0_5275 (.A(n_8_0_6080), .B1(n_8_0_7102), .B2(n_8_0_6733), 
      .ZN(n_8_0_6732));
   INV_X1 i_8_0_5278 (.A(n_8_0_6734), .ZN(n_8_0_6733));
   OR2_X1 i_8_0_5281 (.A1(n_8_0_3477), .A2(n_8_0_784), .ZN(n_8_0_6734));
   NAND2_X1 i_8_0_5284 (.A1(n_8_0_6997), .A2(n_8_0_6405), .ZN(n_8_0_6080));
   AOI21_X1 i_8_0_5287 (.A(n_8_0_6853), .B1(n_8_0_6736), .B2(n_8_0_6735), 
      .ZN(n_224));
   NOR4_X1 i_8_0_5291 (.A1(n_8_0_3331), .A2(n_8_0_3350), .A3(n_8_0_3329), 
      .A4(n_8_0_3352), .ZN(n_8_0_6735));
   OAI221_X1 i_8_0_5292 (.A(n_8_0_4058), .B1(n_8_0_758), .B2(n_8_0_3353), 
      .C1(n_8_0_6622), .C2(n_8_0_6171), .ZN(n_8_0_3352));
   AOI21_X1 i_8_0_5384 (.A(n_8_0_6737), .B1(n_8_0_3338), .B2(n_8_0_6738), 
      .ZN(n_8_0_6736));
   OAI21_X1 i_8_0_5385 (.A(n_8_0_4422), .B1(n_8_0_3478), .B2(n_8_0_752), 
      .ZN(n_8_0_6737));
   INV_X1 i_8_0_5386 (.A(n_8_0_6157), .ZN(n_8_0_6738));
   INV_X1 i_8_0_5387 (.A(n_8_0_6866), .ZN(n_225));
   OAI21_X1 i_8_0_5388 (.A(n_8_0_6854), .B1(n_8_0_6872), .B2(n_8_0_6868), 
      .ZN(n_8_0_6866));
   NAND3_X1 i_8_0_5389 (.A1(n_8_0_3365), .A2(n_8_0_3372), .A3(n_8_0_6870), 
      .ZN(n_8_0_6868));
   AOI211_X1 i_8_0_5390 (.A(n_8_0_3356), .B(n_8_0_3367), .C1(n_8_0_3358), 
      .C2(n_8_0_6871), .ZN(n_8_0_6870));
   OR2_X1 i_8_0_5392 (.A1(n_8_0_3696), .A2(n_8_0_6185), .ZN(n_8_0_6871));
   AOI21_X1 i_8_0_5396 (.A(n_8_0_3373), .B1(n_8_0_6210), .B2(n_8_0_3622), 
      .ZN(n_8_0_3372));
   AOI211_X1 i_8_0_5400 (.A(n_8_0_3366), .B(n_8_0_4346), .C1(n_8_0_6754), 
      .C2(n_8_0_6197), .ZN(n_8_0_3365));
   OAI211_X1 i_8_0_5402 (.A(n_8_0_4422), .B(n_8_0_6987), .C1(n_8_0_7001), 
      .C2(n_8_0_736), .ZN(n_8_0_6872));
   NAND2_X1 i_8_0_5406 (.A1(n_8_0_7102), .A2(n_8_0_6201), .ZN(n_8_0_6987));
   NOR2_X1 i_8_0_5407 (.A1(n_8_0_7098), .A2(n_8_0_7005), .ZN(n_8_0_7001));
   INV_X1 i_8_0_5409 (.A(n_8_0_7090), .ZN(n_8_0_7005));
   NAND3_X1 i_8_0_5576 (.A1(n_8_0_6201), .A2(\out_bs[7] [4]), .A3(n_8_0_3659), 
      .ZN(n_8_0_7090));
   INV_X1 i_8_0_5577 (.A(n_8_0_7380), .ZN(n_8_0_6201));
   INV_X1 i_8_0_5578 (.A(n_8_0_7091), .ZN(n_226));
   OAI21_X1 i_8_0_5579 (.A(n_8_0_6854), .B1(n_8_0_7097), .B2(n_8_0_7092), 
      .ZN(n_8_0_7091));
   OR3_X1 i_8_0_5580 (.A1(n_8_0_7095), .A2(n_8_0_7096), .A3(n_8_0_7093), 
      .ZN(n_8_0_7092));
   NAND4_X1 i_8_0_5582 (.A1(n_8_0_3479), .A2(n_8_0_3466), .A3(n_8_0_3462), 
      .A4(n_8_0_7094), .ZN(n_8_0_7093));
   INV_X1 i_8_0_5583 (.A(n_8_0_3468), .ZN(n_8_0_7094));
   OAI211_X1 i_8_0_5586 (.A(n_8_0_4364), .B(n_8_0_3469), .C1(n_8_0_6772), 
      .C2(n_8_0_6333), .ZN(n_8_0_3468));
   OAI21_X1 i_8_0_5592 (.A(n_8_0_3486), .B1(n_8_0_660), .B2(n_8_0_3485), 
      .ZN(n_8_0_7095));
   INV_X1 i_8_0_5595 (.A(n_8_0_3481), .ZN(n_8_0_7096));
   OAI211_X1 i_8_0_5598 (.A(n_8_0_7099), .B(n_8_0_4422), .C1(n_8_0_657), 
      .C2(n_8_0_3478), .ZN(n_8_0_7097));
   INV_X1 i_8_0_5601 (.A(n_8_0_7098), .ZN(n_8_0_3478));
   NOR2_X1 i_8_0_5602 (.A1(n_8_0_3692), .A2(n_8_0_3658), .ZN(n_8_0_7098));
   INV_X1 i_8_0_5603 (.A(n_8_0_3691), .ZN(n_8_0_3692));
   OAI21_X1 i_8_0_5610 (.A(n_8_0_6362), .B1(n_8_0_7102), .B2(n_8_0_7100), 
      .ZN(n_8_0_7099));
   INV_X1 i_8_0_5613 (.A(n_8_0_7101), .ZN(n_8_0_7100));
   OR2_X1 i_8_0_5614 (.A1(n_8_0_3477), .A2(n_8_0_657), .ZN(n_8_0_7101));
   NAND2_X1 i_8_0_5620 (.A1(\out_bs[7] [4]), .A2(n_8_0_3659), .ZN(n_8_0_3477));
   NOR2_X1 i_8_0_5623 (.A1(n_8_0_6730), .A2(n_8_0_6998), .ZN(n_8_0_7102));
   INV_X1 i_8_0_5624 (.A(n_8_0_7149), .ZN(n_8_0_4422));
   AOI21_X1 i_8_0_5625 (.A(n_8_0_6853), .B1(n_8_0_3554), .B2(n_8_0_7103), 
      .ZN(n_227));
   NOR3_X1 i_8_0_5626 (.A1(n_8_0_3551), .A2(n_8_0_3557), .A3(n_8_0_7104), 
      .ZN(n_8_0_7103));
   OR4_X1 i_8_0_5627 (.A1(n_8_0_7111), .A2(n_8_0_3566), .A3(n_8_0_3561), 
      .A4(n_8_0_7105), .ZN(n_8_0_7104));
   OR4_X1 i_8_0_5629 (.A1(n_8_0_4133), .A2(n_8_0_7106), .A3(n_8_0_3564), 
      .A4(n_8_0_3547), .ZN(n_8_0_7105));
   NAND3_X1 i_8_0_5632 (.A1(n_8_0_7109), .A2(n_8_0_7108), .A3(n_8_0_7107), 
      .ZN(n_8_0_7106));
   INV_X1 i_8_0_5633 (.A(n_8_0_3549), .ZN(n_8_0_7107));
   INV_X1 i_8_0_5634 (.A(n_8_0_3550), .ZN(n_8_0_7108));
   INV_X1 i_8_0_5635 (.A(n_8_0_4232), .ZN(n_8_0_7109));
   NAND2_X1 i_8_0_5636 (.A1(n_8_0_3562), .A2(n_8_0_4364), .ZN(n_8_0_3561));
   INV_X1 i_8_0_5637 (.A(n_8_0_7110), .ZN(n_8_0_3566));
   NAND2_X1 i_8_0_5639 (.A1(n_8_0_3568), .A2(n_8_0_3567), .ZN(n_8_0_7110));
   NAND2_X1 i_8_0_5643 (.A1(n_8_0_7112), .A2(n_8_0_7113), .ZN(n_8_0_7111));
   AOI21_X1 i_8_0_5646 (.A(n_8_0_4059), .B1(n_8_0_3559), .B2(n_8_0_6858), 
      .ZN(n_8_0_7112));
   NAND2_X1 i_8_0_5653 (.A1(n_8_0_3560), .A2(n_8_0_6631), .ZN(n_8_0_7113));
   OAI211_X1 i_8_0_5659 (.A(n_8_0_3803), .B(n_8_0_3598), .C1(n_8_0_3596), 
      .C2(n_8_0_586), .ZN(n_8_0_3557));
   AOI21_X1 i_8_0_5660 (.A(n_8_0_7114), .B1(n_8_0_6729), .B2(n_8_0_7117), 
      .ZN(n_8_0_3554));
   AOI22_X1 i_8_0_5661 (.A1(n_8_0_6730), .A2(n_8_0_7115), .B1(n_8_0_7116), 
      .B2(n_8_0_4424), .ZN(n_8_0_7114));
   INV_X1 i_8_0_5704 (.A(n_8_0_7117), .ZN(n_8_0_7115));
   NAND2_X1 i_8_0_5822 (.A1(\out_bs[7] [4]), .A2(n_8_0_7433), .ZN(n_8_0_7116));
   NOR2_X1 i_8_0_5882 (.A1(n_8_0_578), .A2(n_8_0_3658), .ZN(n_8_0_7117));
   AOI21_X1 i_8_0_5905 (.A(n_8_0_6853), .B1(n_8_0_3580), .B2(n_8_0_7118), 
      .ZN(n_228));
   INV_X1 i_8_0_5956 (.A(n_8_0_7119), .ZN(n_8_0_7118));
   NAND4_X1 i_8_0_6078 (.A1(n_8_0_3574), .A2(n_8_0_7129), .A3(n_8_0_7128), 
      .A4(n_8_0_7120), .ZN(n_8_0_7119));
   AOI211_X1 i_8_0_6152 (.A(n_8_0_7122), .B(n_8_0_7121), .C1(n_8_0_3593), 
      .C2(n_8_0_7127), .ZN(n_8_0_7120));
   NAND4_X1 i_8_0_6191 (.A1(n_8_0_3583), .A2(n_8_0_4132), .A3(n_8_0_3572), 
      .A4(n_8_0_3571), .ZN(n_8_0_7121));
   OAI211_X1 i_8_0_6193 (.A(n_8_0_7126), .B(n_8_0_7125), .C1(n_8_0_7124), 
      .C2(n_8_0_7123), .ZN(n_8_0_7122));
   INV_X1 i_8_0_6201 (.A(n_8_0_5400), .ZN(n_8_0_7123));
   INV_X1 i_8_0_6202 (.A(n_8_0_3589), .ZN(n_8_0_7124));
   INV_X1 i_8_0_6203 (.A(n_8_0_3588), .ZN(n_8_0_7125));
   INV_X1 i_8_0_6204 (.A(n_8_0_6607), .ZN(n_8_0_7126));
   OR2_X1 i_8_0_6207 (.A1(n_8_0_3592), .A2(n_8_0_3685), .ZN(n_8_0_7127));
   INV_X1 i_8_0_6208 (.A(n_8_0_3577), .ZN(n_8_0_7128));
   NAND2_X1 i_8_0_6211 (.A1(n_8_0_4058), .A2(n_8_0_3578), .ZN(n_8_0_3577));
   INV_X1 i_8_0_6212 (.A(n_8_0_3594), .ZN(n_8_0_7129));
   OAI211_X1 i_8_0_6213 (.A(n_8_0_3597), .B(n_8_0_3803), .C1(n_8_0_3595), 
      .C2(n_8_0_554), .ZN(n_8_0_3594));
   NOR2_X1 i_8_0_6214 (.A1(n_8_0_3576), .A2(n_8_0_3575), .ZN(n_8_0_3574));
   AOI21_X1 i_8_0_6215 (.A(n_8_0_7130), .B1(n_8_0_6729), .B2(n_8_0_7133), 
      .ZN(n_8_0_3580));
   AOI22_X1 i_8_0_6216 (.A1(n_8_0_6730), .A2(n_8_0_7132), .B1(n_8_0_4424), 
      .B2(n_8_0_7131), .ZN(n_8_0_7130));
   NAND3_X1 i_8_0_6225 (.A1(\out_bs[7] [4]), .A2(\out_bs[7] [3]), .A3(n_8_0_6542), 
      .ZN(n_8_0_7131));
   INV_X1 i_8_0_6233 (.A(n_8_0_7133), .ZN(n_8_0_7132));
   NOR2_X1 i_8_0_6283 (.A1(n_8_0_3658), .A2(n_8_0_546), .ZN(n_8_0_7133));
   AOI21_X1 i_8_0_6284 (.A(n_8_0_6853), .B1(n_8_0_3601), .B2(n_8_0_7134), 
      .ZN(n_229));
   INV_X1 i_8_0_6296 (.A(n_8_0_7135), .ZN(n_8_0_7134));
   OR4_X1 i_8_0_6323 (.A1(n_8_0_7140), .A2(n_8_0_7139), .A3(n_8_0_3615), 
      .A4(n_8_0_7136), .ZN(n_8_0_7135));
   NAND4_X1 i_8_0_6345 (.A1(n_8_0_3625), .A2(n_8_0_3612), .A3(n_8_0_3607), 
      .A4(n_8_0_7137), .ZN(n_8_0_7136));
   INV_X1 i_8_0_6346 (.A(n_8_0_7138), .ZN(n_8_0_7137));
   OAI211_X1 i_8_0_6347 (.A(n_8_0_3610), .B(n_8_0_4132), .C1(n_8_0_6811), 
      .C2(n_8_0_6593), .ZN(n_8_0_7138));
   OAI221_X1 i_8_0_6348 (.A(n_8_0_3803), .B1(n_8_0_3621), .B2(n_8_0_6681), 
      .C1(n_8_0_3616), .C2(n_8_0_517), .ZN(n_8_0_3615));
   INV_X1 i_8_0_6349 (.A(n_8_0_3628), .ZN(n_8_0_7139));
   INV_X1 i_8_0_6354 (.A(n_8_0_3631), .ZN(n_8_0_7140));
   AOI21_X1 i_8_0_6359 (.A(n_8_0_7141), .B1(n_8_0_6729), .B2(n_8_0_7143), 
      .ZN(n_8_0_3601));
   AOI22_X1 i_8_0_6360 (.A1(n_8_0_6730), .A2(n_8_0_7142), .B1(n_8_0_7432), 
      .B2(n_8_0_4424), .ZN(n_8_0_7141));
   INV_X1 i_8_0_6361 (.A(n_8_0_7143), .ZN(n_8_0_7142));
   NOR2_X1 i_8_0_6362 (.A1(n_8_0_507), .A2(n_8_0_3658), .ZN(n_8_0_7143));
   INV_X1 i_8_0_6363 (.A(n_8_0_3659), .ZN(n_8_0_3658));
   NOR2_X1 i_8_0_6368 (.A1(\out_as[7] [6]), .A2(\out_as[7] [5]), .ZN(n_8_0_3659));
   AOI21_X1 i_8_0_6373 (.A(n_8_0_6853), .B1(n_8_0_3689), .B2(n_8_0_7144), 
      .ZN(n_230));
   INV_X1 i_8_0_6381 (.A(n_8_0_7145), .ZN(n_8_0_7144));
   NAND2_X1 i_8_0_6402 (.A1(n_8_0_3687), .A2(n_8_0_7146), .ZN(n_8_0_7145));
   NOR4_X1 i_8_0_6421 (.A1(n_8_0_3688), .A2(n_8_0_3681), .A3(n_8_0_3682), 
      .A4(n_8_0_7147), .ZN(n_8_0_7146));
   OR4_X1 i_8_0_6422 (.A1(n_8_0_3693), .A2(n_8_0_3694), .A3(n_8_0_4133), 
      .A4(n_8_0_3695), .ZN(n_8_0_7147));
   OAI21_X1 i_8_0_6423 (.A(n_8_0_4364), .B1(n_8_0_957), .B2(n_8_0_4125), 
      .ZN(n_8_0_3694));
   OAI21_X1 i_8_0_6424 (.A(n_8_0_3683), .B1(n_8_0_4472), .B2(n_8_0_956), 
      .ZN(n_8_0_3682));
   OAI21_X1 i_8_0_6425 (.A(n_8_0_4058), .B1(n_8_0_955), .B2(n_8_0_4383), 
      .ZN(n_8_0_3681));
   AOI21_X1 i_8_0_6432 (.A(n_8_0_4346), .B1(n_8_0_4559), .B2(n_8_0_6891), 
      .ZN(n_8_0_3687));
   AOI21_X1 i_8_0_6439 (.A(n_8_0_7149), .B1(n_8_0_3691), .B2(n_8_0_7148), 
      .ZN(n_8_0_3689));
   NOR2_X1 i_8_0_6445 (.A1(n_8_0_952), .A2(\out_as[7] [6]), .ZN(n_8_0_7148));
   NAND2_X1 i_8_0_6446 (.A1(n_8_0_6730), .A2(n_8_0_4424), .ZN(n_8_0_3691));
   NOR2_X1 i_8_0_6447 (.A1(n_8_0_6730), .A2(n_8_0_4424), .ZN(n_8_0_7149));
   NOR2_X1 i_8_0_6448 (.A1(\out_bs[7] [6]), .A2(\out_bs[7] [5]), .ZN(n_8_0_4424));
   AOI21_X1 i_8_0_6449 (.A(n_8_0_6853), .B1(n_8_0_7153), .B2(n_8_0_7150), 
      .ZN(n_231));
   INV_X1 i_8_0_6453 (.A(n_8_0_7151), .ZN(n_8_0_7150));
   OR4_X1 i_8_0_6458 (.A1(n_8_0_3721), .A2(n_8_0_3699), .A3(n_8_0_3702), 
      .A4(n_8_0_7152), .ZN(n_8_0_7151));
   OR4_X1 i_8_0_6479 (.A1(n_8_0_3718), .A2(n_8_0_3705), .A3(n_8_0_6250), 
      .A4(n_8_0_3712), .ZN(n_8_0_7152));
   OAI21_X1 i_8_0_6480 (.A(n_8_0_3706), .B1(n_8_0_948), .B2(n_8_0_4590), 
      .ZN(n_8_0_3705));
   OAI21_X1 i_8_0_6484 (.A(n_8_0_3703), .B1(n_8_0_946), .B2(n_8_0_4571), 
      .ZN(n_8_0_3702));
   OAI21_X1 i_8_0_6485 (.A(n_8_0_3701), .B1(n_8_0_945), .B2(n_8_0_3700), 
      .ZN(n_8_0_3699));
   AOI21_X1 i_8_0_6494 (.A(n_8_0_4409), .B1(n_8_0_7154), .B2(n_8_0_7155), 
      .ZN(n_8_0_7153));
   OAI21_X1 i_8_0_6496 (.A(n_8_0_4503), .B1(n_8_0_6041), .B2(n_8_0_4599), 
      .ZN(n_8_0_7154));
   INV_X1 i_8_0_6504 (.A(n_8_0_7221), .ZN(n_8_0_4503));
   INV_X1 i_8_0_6505 (.A(n_8_0_6042), .ZN(n_8_0_6041));
   NAND2_X1 i_8_0_6506 (.A1(n_8_0_7199), .A2(n_8_0_944), .ZN(n_8_0_7155));
   NAND2_X1 i_8_0_6507 (.A1(n_8_0_6467), .A2(n_8_0_6465), .ZN(n_8_0_4409));
   INV_X1 i_8_0_6508 (.A(n_8_0_7156), .ZN(n_232));
   OAI21_X1 i_8_0_6520 (.A(n_8_0_6854), .B1(n_8_0_7163), .B2(n_8_0_7157), 
      .ZN(n_8_0_7156));
   NAND2_X1 i_8_0_6524 (.A1(n_8_0_3813), .A2(n_8_0_7158), .ZN(n_8_0_7157));
   NOR3_X1 i_8_0_6525 (.A1(n_8_0_3822), .A2(n_8_0_3835), .A3(n_8_0_7159), 
      .ZN(n_8_0_7158));
   OR3_X1 i_8_0_6526 (.A1(n_8_0_3816), .A2(n_8_0_7162), .A3(n_8_0_7160), 
      .ZN(n_8_0_7159));
   NAND3_X1 i_8_0_6527 (.A1(n_8_0_6606), .A2(n_8_0_3830), .A3(n_8_0_7161), 
      .ZN(n_8_0_7160));
   NOR2_X1 i_8_0_6528 (.A1(n_8_0_3831), .A2(n_8_0_3825), .ZN(n_8_0_7161));
   INV_X1 i_8_0_6537 (.A(n_8_0_3828), .ZN(n_8_0_7162));
   OAI211_X1 i_8_0_6544 (.A(n_8_0_3836), .B(n_8_0_3896), .C1(n_8_0_3898), 
      .C2(n_8_0_3838), .ZN(n_8_0_3835));
   NAND2_X1 i_8_0_6550 (.A1(n_8_0_7164), .A2(n_8_0_7165), .ZN(n_8_0_7163));
   AOI21_X1 i_8_0_6611 (.A(n_8_0_6466), .B1(n_8_0_7201), .B2(n_8_0_7167), 
      .ZN(n_8_0_7164));
   OAI211_X1 i_8_0_6612 (.A(n_8_0_4598), .B(n_8_0_7166), .C1(n_8_0_7234), 
      .C2(n_8_0_7167), .ZN(n_8_0_7165));
   OR2_X1 i_8_0_6627 (.A1(n_8_0_5975), .A2(n_8_0_6542), .ZN(n_8_0_7166));
   INV_X1 i_8_0_6628 (.A(n_8_0_912), .ZN(n_8_0_7167));
   INV_X1 i_8_0_6629 (.A(n_8_0_7168), .ZN(n_233));
   OAI21_X1 i_8_0_6634 (.A(n_8_0_6854), .B1(n_8_0_7172), .B2(n_8_0_7169), 
      .ZN(n_8_0_7168));
   OR3_X1 i_8_0_6639 (.A1(n_8_0_7171), .A2(n_8_0_3855), .A3(n_8_0_7170), 
      .ZN(n_8_0_7169));
   NAND4_X1 i_8_0_6640 (.A1(n_8_0_3841), .A2(n_8_0_3860), .A3(n_8_0_3849), 
      .A4(n_8_0_3847), .ZN(n_8_0_7170));
   OAI21_X1 i_8_0_6647 (.A(n_8_0_3865), .B1(n_8_0_905), .B2(n_8_0_3864), 
      .ZN(n_8_0_7171));
   INV_X1 i_8_0_6652 (.A(n_8_0_3856), .ZN(n_8_0_3855));
   OAI211_X1 i_8_0_6653 (.A(n_8_0_7173), .B(n_8_0_6465), .C1(n_8_0_904), 
      .C2(n_8_0_4595), .ZN(n_8_0_7172));
   OAI211_X1 i_8_0_6654 (.A(n_8_0_4598), .B(n_8_0_5674), .C1(n_8_0_7234), 
      .C2(n_8_0_7174), .ZN(n_8_0_7173));
   NAND2_X1 i_8_0_6655 (.A1(n_8_0_5976), .A2(n_8_0_6724), .ZN(n_8_0_5674));
   INV_X1 i_8_0_6657 (.A(n_8_0_904), .ZN(n_8_0_7174));
   INV_X1 i_8_0_6661 (.A(n_8_0_7175), .ZN(n_234));
   OAI21_X1 i_8_0_6666 (.A(n_8_0_6854), .B1(n_8_0_7177), .B2(n_8_0_7176), 
      .ZN(n_8_0_7175));
   OR4_X1 i_8_0_6717 (.A1(n_8_0_3915), .A2(n_8_0_3899), .A3(n_8_0_3895), 
      .A4(n_8_0_3002), .ZN(n_8_0_7176));
   NAND2_X1 i_8_0_6718 (.A1(n_8_0_7178), .A2(n_8_0_7179), .ZN(n_8_0_7177));
   AOI21_X1 i_8_0_6719 (.A(n_8_0_6466), .B1(n_8_0_7201), .B2(n_8_0_7180), 
      .ZN(n_8_0_7178));
   OAI211_X1 i_8_0_6720 (.A(n_8_0_5975), .B(n_8_0_4598), .C1(n_8_0_7234), 
      .C2(n_8_0_7180), .ZN(n_8_0_7179));
   INV_X1 i_8_0_6721 (.A(n_8_0_5976), .ZN(n_8_0_5975));
   INV_X1 i_8_0_6722 (.A(n_8_0_888), .ZN(n_8_0_7180));
   INV_X1 i_8_0_6723 (.A(n_8_0_7181), .ZN(n_235));
   OAI21_X1 i_8_0_6774 (.A(n_8_0_6854), .B1(n_8_0_4001), .B2(n_8_0_7182), 
      .ZN(n_8_0_7181));
   OR4_X1 i_8_0_6794 (.A1(n_8_0_4004), .A2(n_8_0_4013), .A3(n_8_0_4009), 
      .A4(n_8_0_3100), .ZN(n_8_0_7182));
   OAI211_X1 i_8_0_6795 (.A(n_8_0_7183), .B(n_8_0_6465), .C1(n_8_0_856), 
      .C2(n_8_0_4595), .ZN(n_8_0_4001));
   OAI211_X1 i_8_0_6821 (.A(n_8_0_4598), .B(n_8_0_7184), .C1(n_8_0_7234), 
      .C2(n_8_0_7185), .ZN(n_8_0_7183));
   INV_X1 i_8_0_6822 (.A(n_8_0_5954), .ZN(n_8_0_7184));
   NOR2_X1 i_8_0_6823 (.A1(\out_bs[7] [4]), .A2(n_8_0_7433), .ZN(n_8_0_5954));
   INV_X1 i_8_0_6837 (.A(n_8_0_856), .ZN(n_8_0_7185));
   INV_X1 i_8_0_6848 (.A(n_8_0_7186), .ZN(n_236));
   OAI21_X1 i_8_0_6850 (.A(n_8_0_6854), .B1(n_8_0_7191), .B2(n_8_0_7187), 
      .ZN(n_8_0_7186));
   OR3_X1 i_8_0_6852 (.A1(n_8_0_4083), .A2(n_8_0_4101), .A3(n_8_0_7188), 
      .ZN(n_8_0_7187));
   NAND3_X1 i_8_0_6857 (.A1(n_8_0_4096), .A2(n_8_0_7190), .A3(n_8_0_7189), 
      .ZN(n_8_0_7188));
   AOI211_X1 i_8_0_6869 (.A(n_8_0_4078), .B(n_8_0_4093), .C1(n_8_0_6597), 
      .C2(n_8_0_6664), .ZN(n_8_0_7189));
   INV_X1 i_8_0_6870 (.A(n_8_0_4090), .ZN(n_8_0_7190));
   OAI211_X1 i_8_0_6871 (.A(n_8_0_6577), .B(n_8_0_4091), .C1(n_8_0_836), 
      .C2(n_8_0_4590), .ZN(n_8_0_4090));
   AOI21_X1 i_8_0_6970 (.A(n_8_0_4097), .B1(n_8_0_4543), .B2(n_8_0_6911), 
      .ZN(n_8_0_4096));
   OAI21_X1 i_8_0_6971 (.A(n_8_0_4084), .B1(n_8_0_833), .B2(n_8_0_4085), 
      .ZN(n_8_0_4083));
   OAI211_X1 i_8_0_6975 (.A(n_8_0_7192), .B(n_8_0_6465), .C1(n_8_0_832), 
      .C2(n_8_0_4595), .ZN(n_8_0_7191));
   OAI211_X1 i_8_0_6976 (.A(n_8_0_5973), .B(n_8_0_4598), .C1(n_8_0_7234), 
      .C2(n_8_0_7193), .ZN(n_8_0_7192));
   INV_X1 i_8_0_6977 (.A(n_8_0_4599), .ZN(n_8_0_4598));
   NAND2_X1 i_8_0_6980 (.A1(n_8_0_3710), .A2(\out_bs[7] [5]), .ZN(n_8_0_4599));
   INV_X1 i_8_0_6983 (.A(n_8_0_832), .ZN(n_8_0_7193));
   AOI21_X1 i_8_0_6985 (.A(n_8_0_6853), .B1(n_8_0_7197), .B2(n_8_0_7194), 
      .ZN(n_237));
   AND2_X1 i_8_0_6986 (.A1(n_8_0_7196), .A2(n_8_0_7195), .ZN(n_8_0_7194));
   NOR4_X1 i_8_0_6987 (.A1(n_8_0_4150), .A2(n_8_0_4153), .A3(n_8_0_4148), 
      .A4(n_8_0_4138), .ZN(n_8_0_7195));
   INV_X1 i_8_0_6988 (.A(n_8_0_4157), .ZN(n_8_0_7196));
   INV_X1 i_8_0_6989 (.A(n_8_0_7198), .ZN(n_8_0_7197));
   OAI211_X1 i_8_0_6990 (.A(n_8_0_7200), .B(n_8_0_6465), .C1(n_8_0_6998), 
      .C2(n_8_0_7199), .ZN(n_8_0_7198));
   NAND2_X1 i_8_0_6991 (.A1(n_8_0_7234), .A2(n_8_0_6042), .ZN(n_8_0_7199));
   OAI211_X1 i_8_0_6992 (.A(n_8_0_7221), .B(n_8_0_7202), .C1(n_8_0_7201), 
      .C2(n_8_0_6042), .ZN(n_8_0_7200));
   INV_X1 i_8_0_6993 (.A(n_8_0_4595), .ZN(n_8_0_7201));
   INV_X1 i_8_0_6994 (.A(n_8_0_801), .ZN(n_8_0_7202));
   INV_X1 i_8_0_7008 (.A(n_8_0_7203), .ZN(n_238));
   OAI21_X1 i_8_0_7011 (.A(n_8_0_6854), .B1(n_8_0_7205), .B2(n_8_0_7204), 
      .ZN(n_8_0_7203));
   OR4_X1 i_8_0_7067 (.A1(n_8_0_4204), .A2(n_8_0_4191), .A3(n_8_0_4214), 
      .A4(n_8_0_4209), .ZN(n_8_0_7204));
   OAI211_X1 i_8_0_7109 (.A(n_8_0_7206), .B(n_8_0_6465), .C1(n_8_0_769), 
      .C2(n_8_0_4595), .ZN(n_8_0_7205));
   OAI21_X1 i_8_0_7110 (.A(n_8_0_6118), .B1(n_8_0_6468), .B2(n_8_0_7207), 
      .ZN(n_8_0_7206));
   INV_X1 i_8_0_7115 (.A(n_8_0_7208), .ZN(n_8_0_7207));
   OR2_X1 i_8_0_7122 (.A1(n_8_0_4532), .A2(n_8_0_769), .ZN(n_8_0_7208));
   INV_X1 i_8_0_7124 (.A(n_8_0_6117), .ZN(n_8_0_6118));
   INV_X1 i_8_0_7126 (.A(n_8_0_7209), .ZN(n_239));
   OAI21_X1 i_8_0_7127 (.A(n_8_0_6854), .B1(n_8_0_4370), .B2(n_8_0_7210), 
      .ZN(n_8_0_7209));
   NAND4_X1 i_8_0_7128 (.A1(n_8_0_4373), .A2(n_8_0_4376), .A3(n_8_0_7213), 
      .A4(n_8_0_7211), .ZN(n_8_0_7210));
   NOR4_X1 i_8_0_7243 (.A1(n_8_0_4380), .A2(n_8_0_4386), .A3(n_8_0_7212), 
      .A4(n_8_0_4363), .ZN(n_8_0_7211));
   OAI221_X1 i_8_0_7244 (.A(n_8_0_6606), .B1(n_8_0_6282), .B2(n_8_0_6333), 
      .C1(n_8_0_4368), .C2(n_8_0_673), .ZN(n_8_0_4363));
   INV_X1 i_8_0_7245 (.A(n_8_0_4357), .ZN(n_8_0_7212));
   OR2_X1 i_8_0_7252 (.A1(n_8_0_4571), .A2(n_8_0_664), .ZN(n_8_0_7213));
   OAI211_X1 i_8_0_7253 (.A(n_8_0_7214), .B(n_8_0_6465), .C1(n_8_0_658), 
      .C2(n_8_0_4595), .ZN(n_8_0_4370));
   NAND3_X1 i_8_0_7254 (.A1(n_8_0_7215), .A2(\out_bs[7] [3]), .A3(n_8_0_6363), 
      .ZN(n_8_0_7214));
   OAI21_X1 i_8_0_7255 (.A(n_8_0_6467), .B1(n_8_0_658), .B2(n_8_0_4532), 
      .ZN(n_8_0_7215));
   INV_X1 i_8_0_7256 (.A(n_8_0_7216), .ZN(n_240));
   OAI21_X1 i_8_0_7257 (.A(n_8_0_6854), .B1(n_8_0_7218), .B2(n_8_0_7217), 
      .ZN(n_8_0_7216));
   OR4_X1 i_8_0_7259 (.A1(n_8_0_4405), .A2(n_8_0_4398), .A3(n_8_0_4397), 
      .A4(n_8_0_4389), .ZN(n_8_0_7217));
   OAI21_X1 i_8_0_7260 (.A(n_8_0_7219), .B1(n_8_0_6467), .B2(n_8_0_7222), 
      .ZN(n_8_0_7218));
   AOI21_X1 i_8_0_7261 (.A(n_8_0_6466), .B1(n_8_0_7220), .B2(n_8_0_7221), 
      .ZN(n_8_0_7219));
   AOI21_X1 i_8_0_7346 (.A(n_8_0_634), .B1(n_8_0_4595), .B2(n_8_0_6403), 
      .ZN(n_8_0_7220));
   NAND2_X1 i_8_0_7347 (.A1(n_8_0_4595), .A2(n_8_0_4532), .ZN(n_8_0_7221));
   NAND2_X1 i_8_0_7348 (.A1(n_8_0_4600), .A2(\out_bs[7] [4]), .ZN(n_8_0_4532));
   NAND2_X1 i_8_0_7349 (.A1(\out_bs[7] [3]), .A2(n_8_0_7223), .ZN(n_8_0_7222));
   INV_X1 i_8_0_7350 (.A(n_8_0_6405), .ZN(n_8_0_7223));
   INV_X1 i_8_0_7351 (.A(n_8_0_7224), .ZN(n_241));
   OAI21_X1 i_8_0_7352 (.A(n_8_0_6854), .B1(n_8_0_4468), .B2(n_8_0_7225), 
      .ZN(n_8_0_7224));
   OR4_X1 i_8_0_7353 (.A1(n_8_0_4455), .A2(n_8_0_4445), .A3(n_8_0_4448), 
      .A4(n_8_0_7226), .ZN(n_8_0_7225));
   OR2_X1 i_8_0_7354 (.A1(n_8_0_4471), .A2(n_8_0_7227), .ZN(n_8_0_7226));
   OR4_X1 i_8_0_7355 (.A1(n_8_0_7229), .A2(n_8_0_4452), .A3(n_8_0_4465), 
      .A4(n_8_0_7228), .ZN(n_8_0_7227));
   OAI21_X1 i_8_0_7356 (.A(n_8_0_6249), .B1(n_8_0_4514), .B2(n_8_0_607), 
      .ZN(n_8_0_7228));
   OAI221_X1 i_8_0_7357 (.A(n_8_0_6526), .B1(n_8_0_6689), .B2(n_8_0_6321), 
      .C1(n_8_0_4466), .C2(n_8_0_603), .ZN(n_8_0_4465));
   INV_X1 i_8_0_7358 (.A(n_8_0_4461), .ZN(n_8_0_7229));
   OAI221_X1 i_8_0_7359 (.A(n_8_0_6577), .B1(n_8_0_4473), .B2(n_8_0_595), 
      .C1(n_8_0_6325), .C2(n_8_0_5467), .ZN(n_8_0_4471));
   OAI211_X1 i_8_0_7360 (.A(n_8_0_7233), .B(n_8_0_6465), .C1(n_8_0_579), 
      .C2(n_8_0_4595), .ZN(n_8_0_4468));
   NAND2_X1 i_8_0_7361 (.A1(n_8_0_7230), .A2(n_8_0_7232), .ZN(n_8_0_4595));
   OR2_X1 i_8_0_7362 (.A1(n_8_0_7422), .A2(n_8_0_7231), .ZN(n_8_0_7230));
   NAND2_X1 i_8_0_7363 (.A1(n_8_0_7000), .A2(n_8_0_6854), .ZN(n_8_0_7231));
   INV_X1 i_8_0_7364 (.A(\out_as[7] [6]), .ZN(n_8_0_7232));
   INV_X1 i_8_0_7365 (.A(n_8_0_6466), .ZN(n_8_0_6465));
   NOR2_X1 i_8_0_7366 (.A1(n_8_0_7251), .A2(n_8_0_7000), .ZN(n_8_0_6466));
   OAI21_X1 i_8_0_7367 (.A(n_8_0_7433), .B1(n_8_0_6468), .B2(n_8_0_7235), 
      .ZN(n_8_0_7233));
   INV_X1 i_8_0_7368 (.A(n_8_0_6467), .ZN(n_8_0_6468));
   NAND2_X1 i_8_0_7369 (.A1(n_8_0_7234), .A2(\out_bs[7] [4]), .ZN(n_8_0_6467));
   AOI21_X1 i_8_0_7370 (.A(n_8_0_6999), .B1(n_8_0_7421), .B2(n_8_0_6854), 
      .ZN(n_8_0_7234));
   INV_X1 i_8_0_7371 (.A(n_8_0_7236), .ZN(n_8_0_7235));
   NAND3_X1 i_8_0_7372 (.A1(n_8_0_4600), .A2(\out_bs[7] [4]), .A3(n_8_0_7237), 
      .ZN(n_8_0_7236));
   INV_X1 i_8_0_7373 (.A(n_8_0_579), .ZN(n_8_0_7237));
   AOI21_X1 i_8_0_7374 (.A(n_8_0_6853), .B1(n_8_0_7243), .B2(n_8_0_7238), 
      .ZN(n_242));
   AOI21_X1 i_8_0_7375 (.A(n_8_0_7239), .B1(\out_bs[7] [6]), .B2(n_8_0_7244), 
      .ZN(n_8_0_7238));
   OR4_X1 i_8_0_7376 (.A1(n_8_0_4625), .A2(n_8_0_4623), .A3(n_8_0_4624), 
      .A4(n_8_0_7240), .ZN(n_8_0_7239));
   NAND2_X1 i_8_0_7377 (.A1(n_8_0_4619), .A2(n_8_0_7241), .ZN(n_8_0_7240));
   NOR3_X1 i_8_0_7378 (.A1(n_8_0_4617), .A2(n_8_0_4618), .A3(n_8_0_7242), 
      .ZN(n_8_0_7241));
   OAI21_X1 i_8_0_7379 (.A(n_8_0_6249), .B1(n_8_0_5274), .B2(n_8_0_5), .ZN(
      n_8_0_7242));
   AOI21_X1 i_8_0_7380 (.A(n_8_0_5395), .B1(n_8_0_6526), .B2(n_8_0_63), .ZN(
      n_8_0_4618));
   AOI21_X1 i_8_0_7381 (.A(n_8_0_5428), .B1(n_8_0_6606), .B2(n_8_0_126), 
      .ZN(n_8_0_4617));
   NOR2_X1 i_8_0_7382 (.A1(n_8_0_6578), .A2(n_8_0_4620), .ZN(n_8_0_4619));
   OAI21_X1 i_8_0_7383 (.A(n_8_0_6556), .B1(n_8_0_252), .B2(n_8_0_5460), 
      .ZN(n_8_0_4624));
   AOI21_X1 i_8_0_7384 (.A(n_8_0_5302), .B1(n_8_0_6513), .B2(n_8_0_315), 
      .ZN(n_8_0_4623));
   OAI21_X1 i_8_0_7385 (.A(n_8_0_6590), .B1(n_8_0_378), .B2(n_8_0_5456), 
      .ZN(n_8_0_4625));
   OAI21_X1 i_8_0_7386 (.A(n_8_0_6731), .B1(\out_bs[7] [6]), .B2(n_8_0_7244), 
      .ZN(n_8_0_7243));
   INV_X1 i_8_0_7387 (.A(n_8_0_441), .ZN(n_8_0_7244));
   AOI21_X1 i_8_0_7388 (.A(n_8_0_6853), .B1(n_8_0_4820), .B2(n_8_0_7245), 
      .ZN(n_243));
   INV_X1 i_8_0_7389 (.A(n_8_0_7246), .ZN(n_8_0_7245));
   NAND3_X1 i_8_0_7390 (.A1(n_8_0_7249), .A2(n_8_0_4816), .A3(n_8_0_7247), 
      .ZN(n_8_0_7246));
   NOR3_X1 i_8_0_7391 (.A1(n_8_0_4842), .A2(n_8_0_4827), .A3(n_8_0_7248), 
      .ZN(n_8_0_7247));
   OR3_X1 i_8_0_7392 (.A1(n_8_0_4831), .A2(n_8_0_4837), .A3(n_8_0_4841), 
      .ZN(n_8_0_7248));
   OAI21_X1 i_8_0_7393 (.A(n_8_0_4828), .B1(n_8_0_6837), .B2(n_8_0_197), 
      .ZN(n_8_0_4827));
   OAI21_X1 i_8_0_7394 (.A(n_8_0_4817), .B1(n_8_0_6825), .B2(n_8_0_4819), 
      .ZN(n_8_0_4816));
   INV_X1 i_8_0_7395 (.A(n_8_0_4824), .ZN(n_8_0_7249));
   OAI21_X1 i_8_0_7396 (.A(n_8_0_4825), .B1(n_8_0_386), .B2(n_8_0_6755), 
      .ZN(n_8_0_4824));
   OAI21_X1 i_8_0_7397 (.A(n_8_0_7250), .B1(n_8_0_6729), .B2(n_8_0_7253), 
      .ZN(n_8_0_4820));
   OAI21_X1 i_8_0_7398 (.A(n_8_0_449), .B1(n_8_0_7251), .B2(n_8_0_7254), 
      .ZN(n_8_0_7250));
   INV_X1 i_8_0_7399 (.A(n_8_0_7252), .ZN(n_8_0_7251));
   NAND2_X1 i_8_0_7400 (.A1(n_8_0_3882), .A2(n_8_0_6854), .ZN(n_8_0_7252));
   INV_X1 i_8_0_7401 (.A(n_8_0_7254), .ZN(n_8_0_7253));
   NAND2_X1 i_8_0_7402 (.A1(\out_bs[7] [6]), .A2(n_8_0_4823), .ZN(n_8_0_7254));
   NAND2_X1 i_8_0_7403 (.A1(n_8_0_5976), .A2(n_8_0_6999), .ZN(n_8_0_4823));
   AOI21_X1 i_8_0_7404 (.A(n_8_0_6853), .B1(n_8_0_7262), .B2(n_8_0_7255), 
      .ZN(n_244));
   NOR3_X1 i_8_0_7405 (.A1(n_8_0_4857), .A2(n_8_0_4867), .A3(n_8_0_7256), 
      .ZN(n_8_0_7255));
   NAND2_X1 i_8_0_7406 (.A1(n_8_0_4864), .A2(n_8_0_7257), .ZN(n_8_0_7256));
   INV_X1 i_8_0_7407 (.A(n_8_0_7258), .ZN(n_8_0_7257));
   OR4_X1 i_8_0_7408 (.A1(n_8_0_4854), .A2(n_8_0_4861), .A3(n_8_0_4870), 
      .A4(n_8_0_4851), .ZN(n_8_0_7258));
   INV_X1 i_8_0_7409 (.A(n_8_0_7259), .ZN(n_8_0_4851));
   NAND2_X1 i_8_0_7410 (.A1(n_8_0_7260), .A2(n_8_0_7261), .ZN(n_8_0_7259));
   AOI21_X1 i_8_0_7411 (.A(n_8_0_5428), .B1(n_8_0_4852), .B2(n_8_0_7059), 
      .ZN(n_8_0_7260));
   NAND2_X1 i_8_0_7412 (.A1(n_8_0_6606), .A2(n_8_0_135), .ZN(n_8_0_7261));
   OAI21_X1 i_8_0_7413 (.A(n_8_0_4862), .B1(n_8_0_6837), .B2(n_8_0_198), 
      .ZN(n_8_0_4861));
   OAI21_X1 i_8_0_7414 (.A(n_8_0_4866), .B1(n_8_0_4865), .B2(n_8_0_5223), 
      .ZN(n_8_0_4864));
   OAI21_X1 i_8_0_7415 (.A(n_8_0_4868), .B1(n_8_0_6824), .B2(n_8_0_324), 
      .ZN(n_8_0_4867));
   INV_X1 i_8_0_7416 (.A(n_8_0_4848), .ZN(n_8_0_7262));
   AND2_X1 i_8_0_7417 (.A1(n_8_0_7264), .A2(n_8_0_7263), .ZN(n_8_0_4848));
   NAND2_X1 i_8_0_7418 (.A1(n_8_0_7265), .A2(n_8_0_450), .ZN(n_8_0_7263));
   OAI21_X1 i_8_0_7419 (.A(n_8_0_6730), .B1(n_8_0_450), .B2(n_8_0_7265), 
      .ZN(n_8_0_7264));
   OAI21_X1 i_8_0_7420 (.A(\out_bs[7] [6]), .B1(n_8_0_5056), .B2(n_8_0_6362), 
      .ZN(n_8_0_7265));
   NAND2_X1 i_8_0_7421 (.A1(n_8_0_6999), .A2(n_8_0_6998), .ZN(n_8_0_5056));
   INV_X1 i_8_0_7422 (.A(n_8_0_7266), .ZN(n_8_0_6362));
   OAI21_X1 i_8_0_7423 (.A(\out_bs[7] [3]), .B1(\out_bs[7] [2]), .B2(n_8_0_7381), 
      .ZN(n_8_0_7266));
   AOI21_X1 i_8_0_7424 (.A(n_8_0_6853), .B1(n_8_0_7267), .B2(n_8_0_7280), 
      .ZN(n_245));
   INV_X1 i_8_0_7425 (.A(n_8_0_7268), .ZN(n_8_0_7267));
   OAI211_X1 i_8_0_7426 (.A(n_8_0_7278), .B(n_8_0_7269), .C1(n_8_0_6232), 
      .C2(n_8_0_5081), .ZN(n_8_0_7268));
   NOR4_X1 i_8_0_7427 (.A1(n_8_0_5069), .A2(n_8_0_5065), .A3(n_8_0_5082), 
      .A4(n_8_0_7270), .ZN(n_8_0_7269));
   NAND3_X1 i_8_0_7428 (.A1(n_8_0_5077), .A2(n_8_0_5074), .A3(n_8_0_7271), 
      .ZN(n_8_0_7270));
   NOR2_X1 i_8_0_7429 (.A1(n_8_0_7276), .A2(n_8_0_7272), .ZN(n_8_0_7271));
   OAI21_X1 i_8_0_7430 (.A(n_8_0_6247), .B1(n_8_0_6249), .B2(n_8_0_6054), 
      .ZN(n_8_0_7272));
   INV_X1 i_8_0_7431 (.A(n_8_0_7273), .ZN(n_8_0_6054));
   NAND2_X1 i_8_0_7432 (.A1(n_8_0_7275), .A2(n_8_0_7274), .ZN(n_8_0_7273));
   NAND2_X1 i_8_0_7433 (.A1(\out_bs[0] [4]), .A2(\out_bs[0] [0]), .ZN(n_8_0_7274));
   INV_X1 i_8_0_7434 (.A(n_8_0_6082), .ZN(n_8_0_7275));
   AOI21_X1 i_8_0_7435 (.A(n_8_0_17), .B1(n_8_0_6595), .B2(n_8_0_6052), .ZN(
      n_8_0_7276));
   NAND2_X1 i_8_0_7436 (.A1(n_8_0_5076), .A2(n_8_0_5075), .ZN(n_8_0_5074));
   OAI21_X1 i_8_0_7437 (.A(n_8_0_5078), .B1(n_8_0_5079), .B2(n_8_0_6605), 
      .ZN(n_8_0_5077));
   OR2_X1 i_8_0_7438 (.A1(n_8_0_5084), .A2(n_8_0_5083), .ZN(n_8_0_5082));
   OAI22_X1 i_8_0_7439 (.A1(n_8_0_7277), .A2(n_8_0_5066), .B1(n_8_0_5067), 
      .B2(n_8_0_7294), .ZN(n_8_0_5065));
   OR2_X1 i_8_0_7440 (.A1(n_8_0_5221), .A2(n_8_0_269), .ZN(n_8_0_7277));
   INV_X1 i_8_0_7441 (.A(n_8_0_5071), .ZN(n_8_0_7278));
   NAND2_X1 i_8_0_7442 (.A1(n_8_0_7279), .A2(n_8_0_5072), .ZN(n_8_0_5071));
   OR2_X1 i_8_0_7443 (.A1(n_8_0_6755), .A2(n_8_0_395), .ZN(n_8_0_7279));
   OAI21_X1 i_8_0_7444 (.A(n_8_0_7282), .B1(n_8_0_6233), .B2(n_8_0_7281), 
      .ZN(n_8_0_7280));
   INV_X1 i_8_0_7445 (.A(n_8_0_5081), .ZN(n_8_0_7281));
   AOI21_X1 i_8_0_7446 (.A(n_8_0_6728), .B1(n_8_0_6717), .B2(n_8_0_6042), 
      .ZN(n_8_0_5081));
   NAND2_X1 i_8_0_7447 (.A1(n_8_0_6157), .A2(n_8_0_6544), .ZN(n_8_0_6042));
   NOR2_X1 i_8_0_7448 (.A1(\out_bs[7] [3]), .A2(\out_bs[7] [2]), .ZN(n_8_0_6157));
   INV_X1 i_8_0_7449 (.A(n_8_0_458), .ZN(n_8_0_7282));
   AOI21_X1 i_8_0_7450 (.A(n_8_0_6853), .B1(n_8_0_7296), .B2(n_8_0_7283), 
      .ZN(n_246));
   NOR3_X1 i_8_0_7451 (.A1(n_8_0_5192), .A2(n_8_0_7295), .A3(n_8_0_7284), 
      .ZN(n_8_0_7283));
   OR4_X1 i_8_0_7452 (.A1(n_8_0_5176), .A2(n_8_0_5195), .A3(n_8_0_5178), 
      .A4(n_8_0_7285), .ZN(n_8_0_7284));
   NAND3_X1 i_8_0_7453 (.A1(n_8_0_7289), .A2(n_8_0_5188), .A3(n_8_0_7286), 
      .ZN(n_8_0_7285));
   AOI21_X1 i_8_0_7454 (.A(n_8_0_7287), .B1(n_8_0_7288), .B2(n_8_0_7393), 
      .ZN(n_8_0_7286));
   AOI211_X1 i_8_0_7455 (.A(n_8_0_7085), .B(n_8_0_5191), .C1(n_8_0_6812), 
      .C2(n_8_0_21), .ZN(n_8_0_7287));
   INV_X1 i_8_0_7456 (.A(n_8_0_21), .ZN(n_8_0_7288));
   OAI21_X1 i_8_0_7457 (.A(n_8_0_5189), .B1(n_8_0_5190), .B2(\out_bs[1] [5]), 
      .ZN(n_8_0_5188));
   OAI221_X1 i_8_0_7458 (.A(n_8_0_7341), .B1(n_8_0_7291), .B2(n_8_0_7340), 
      .C1(n_8_0_7290), .C2(n_8_0_7292), .ZN(n_8_0_7289));
   INV_X1 i_8_0_7459 (.A(n_8_0_5187), .ZN(n_8_0_7290));
   INV_X1 i_8_0_7460 (.A(n_8_0_6182), .ZN(n_8_0_7291));
   INV_X1 i_8_0_7461 (.A(n_8_0_147), .ZN(n_8_0_7292));
   OAI21_X1 i_8_0_7462 (.A(n_8_0_5179), .B1(n_8_0_6837), .B2(n_8_0_210), 
      .ZN(n_8_0_5178));
   OAI22_X1 i_8_0_7463 (.A1(n_8_0_7293), .A2(n_8_0_5196), .B1(n_8_0_5197), 
      .B2(n_8_0_7294), .ZN(n_8_0_5195));
   OR2_X1 i_8_0_7464 (.A1(n_8_0_5221), .A2(n_8_0_273), .ZN(n_8_0_7293));
   OR2_X1 i_8_0_7465 (.A1(n_8_0_6556), .A2(n_8_0_5224), .ZN(n_8_0_7294));
   OAI221_X1 i_8_0_7466 (.A(n_8_0_6511), .B1(n_8_0_5470), .B2(n_8_0_6211), 
      .C1(n_8_0_5177), .C2(n_8_0_336), .ZN(n_8_0_5176));
   INV_X1 i_8_0_7467 (.A(n_8_0_5182), .ZN(n_8_0_7295));
   OAI21_X1 i_8_0_7468 (.A(n_8_0_5184), .B1(n_8_0_6754), .B2(n_8_0_5183), 
      .ZN(n_8_0_5182));
   NOR2_X1 i_8_0_7469 (.A1(n_8_0_5194), .A2(n_8_0_462), .ZN(n_8_0_5192));
   NAND2_X1 i_8_0_7470 (.A1(n_8_0_6233), .A2(n_8_0_5193), .ZN(n_8_0_7296));
   NAND2_X1 i_8_0_7471 (.A1(n_8_0_5194), .A2(n_8_0_462), .ZN(n_8_0_5193));
   INV_X1 i_8_0_7472 (.A(n_8_0_7297), .ZN(n_247));
   OAI21_X1 i_8_0_7473 (.A(n_8_0_6854), .B1(n_8_0_7298), .B2(n_8_0_7307), 
      .ZN(n_8_0_7297));
   OAI211_X1 i_8_0_7474 (.A(n_8_0_5368), .B(n_8_0_7299), .C1(n_8_0_6232), 
      .C2(n_8_0_469), .ZN(n_8_0_7298));
   INV_X1 i_8_0_7475 (.A(n_8_0_7300), .ZN(n_8_0_7299));
   OR3_X1 i_8_0_7476 (.A1(n_8_0_5377), .A2(n_8_0_5371), .A3(n_8_0_7301), 
      .ZN(n_8_0_7300));
   OAI211_X1 i_8_0_7477 (.A(n_8_0_5375), .B(n_8_0_7302), .C1(n_8_0_6837), 
      .C2(n_8_0_217), .ZN(n_8_0_7301));
   AOI221_X1 i_8_0_7478 (.A(n_8_0_5365), .B1(n_8_0_7304), .B2(n_8_0_7303), 
      .C1(n_8_0_7305), .C2(n_8_0_5363), .ZN(n_8_0_7302));
   OAI211_X1 i_8_0_7479 (.A(n_8_0_6525), .B(n_8_0_5366), .C1(n_8_0_6265), 
      .C2(n_8_0_91), .ZN(n_8_0_5365));
   OAI21_X1 i_8_0_7480 (.A(n_8_0_5360), .B1(n_8_0_28), .B2(n_8_0_6595), .ZN(
      n_8_0_7303));
   NAND2_X1 i_8_0_7481 (.A1(n_8_0_6812), .A2(n_8_0_28), .ZN(n_8_0_7304));
   AND2_X1 i_8_0_7482 (.A1(n_8_0_7306), .A2(n_8_0_5427), .ZN(n_8_0_7305));
   OR2_X1 i_8_0_7483 (.A1(n_8_0_5425), .A2(n_8_0_6707), .ZN(n_8_0_7306));
   AOI21_X1 i_8_0_7484 (.A(n_8_0_5372), .B1(n_8_0_280), .B2(n_8_0_5373), 
      .ZN(n_8_0_5371));
   OAI211_X1 i_8_0_7485 (.A(n_8_0_6511), .B(n_8_0_5378), .C1(n_8_0_343), 
      .C2(n_8_0_6376), .ZN(n_8_0_5377));
   AOI21_X1 i_8_0_7486 (.A(n_8_0_5480), .B1(n_8_0_6232), .B2(n_8_0_469), 
      .ZN(n_8_0_7307));
   AOI21_X1 i_8_0_7487 (.A(n_8_0_6728), .B1(n_8_0_6717), .B2(n_8_0_7433), 
      .ZN(n_8_0_5480));
   INV_X1 i_8_0_7488 (.A(n_8_0_7308), .ZN(n_248));
   OAI21_X1 i_8_0_7489 (.A(n_8_0_6854), .B1(n_8_0_7309), .B2(n_8_0_7325), 
      .ZN(n_8_0_7308));
   OAI211_X1 i_8_0_7490 (.A(n_8_0_5382), .B(n_8_0_7310), .C1(n_8_0_6232), 
      .C2(n_8_0_5403), .ZN(n_8_0_7309));
   INV_X1 i_8_0_7491 (.A(n_8_0_7311), .ZN(n_8_0_7310));
   OAI211_X1 i_8_0_7492 (.A(n_8_0_7323), .B(n_8_0_7312), .C1(n_8_0_5406), 
      .C2(n_8_0_344), .ZN(n_8_0_7311));
   NOR4_X1 i_8_0_7493 (.A1(n_8_0_5407), .A2(n_8_0_5388), .A3(n_8_0_5398), 
      .A4(n_8_0_7313), .ZN(n_8_0_7312));
   OAI21_X1 i_8_0_7494 (.A(n_8_0_7314), .B1(n_8_0_29), .B2(n_8_0_6595), .ZN(
      n_8_0_7313));
   OAI221_X1 i_8_0_7495 (.A(n_8_0_7316), .B1(n_8_0_7319), .B2(n_8_0_7317), 
      .C1(n_8_0_7315), .C2(n_8_0_7318), .ZN(n_8_0_7314));
   INV_X1 i_8_0_7496 (.A(n_8_0_5393), .ZN(n_8_0_7315));
   INV_X1 i_8_0_7497 (.A(n_8_0_5395), .ZN(n_8_0_7316));
   INV_X1 i_8_0_7498 (.A(n_8_0_6526), .ZN(n_8_0_7317));
   INV_X1 i_8_0_7499 (.A(n_8_0_6530), .ZN(n_8_0_7318));
   INV_X1 i_8_0_7500 (.A(n_8_0_92), .ZN(n_8_0_7319));
   INV_X1 i_8_0_7501 (.A(n_8_0_7320), .ZN(n_8_0_5398));
   OAI21_X1 i_8_0_7502 (.A(n_8_0_7321), .B1(n_8_0_7322), .B2(n_8_0_7370), 
      .ZN(n_8_0_7320));
   INV_X1 i_8_0_7503 (.A(n_8_0_5399), .ZN(n_8_0_7321));
   INV_X1 i_8_0_7504 (.A(n_8_0_155), .ZN(n_8_0_7322));
   OAI211_X1 i_8_0_7505 (.A(n_8_0_6575), .B(n_8_0_5389), .C1(n_8_0_6572), 
      .C2(n_8_0_218), .ZN(n_8_0_5388));
   AOI221_X1 i_8_0_7506 (.A(n_8_0_5460), .B1(n_8_0_281), .B2(n_8_0_5408), 
      .C1(n_8_0_6795), .C2(n_8_0_5409), .ZN(n_8_0_5407));
   INV_X1 i_8_0_7507 (.A(n_8_0_7324), .ZN(n_8_0_7323));
   OAI21_X1 i_8_0_7508 (.A(n_8_0_6511), .B1(n_8_0_6515), .B2(n_8_0_5470), 
      .ZN(n_8_0_7324));
   AOI21_X1 i_8_0_7509 (.A(n_8_0_470), .B1(n_8_0_6232), .B2(n_8_0_5403), 
      .ZN(n_8_0_7325));
   INV_X1 i_8_0_7510 (.A(n_8_0_5404), .ZN(n_8_0_5403));
   OAI21_X1 i_8_0_7511 (.A(n_8_0_6727), .B1(n_8_0_6716), .B2(n_8_0_6540), 
      .ZN(n_8_0_5404));
   NAND2_X1 i_8_0_7512 (.A1(n_8_0_6542), .A2(\out_bs[7] [3]), .ZN(n_8_0_6540));
   INV_X1 i_8_0_7513 (.A(n_8_0_7326), .ZN(n_249));
   NAND2_X1 i_8_0_7514 (.A1(n_8_0_7327), .A2(n_8_0_6854), .ZN(n_8_0_7326));
   NAND4_X1 i_8_0_7515 (.A1(n_8_0_7343), .A2(n_8_0_5433), .A3(n_8_0_5420), 
      .A4(n_8_0_7328), .ZN(n_8_0_7327));
   INV_X1 i_8_0_7516 (.A(n_8_0_7329), .ZN(n_8_0_7328));
   OR3_X1 i_8_0_7517 (.A1(n_8_0_5416), .A2(n_8_0_5438), .A3(n_8_0_7330), 
      .ZN(n_8_0_7329));
   NAND3_X1 i_8_0_7518 (.A1(n_8_0_5414), .A2(n_8_0_7337), .A3(n_8_0_7331), 
      .ZN(n_8_0_7330));
   INV_X1 i_8_0_7519 (.A(n_8_0_7332), .ZN(n_8_0_7331));
   OR3_X1 i_8_0_7520 (.A1(n_8_0_5430), .A2(n_8_0_7334), .A3(n_8_0_7333), 
      .ZN(n_8_0_7332));
   OAI21_X1 i_8_0_7521 (.A(n_8_0_6247), .B1(n_8_0_6249), .B2(n_8_0_6593), 
      .ZN(n_8_0_7333));
   NAND2_X1 i_8_0_7522 (.A1(n_8_0_6813), .A2(\out_bs[0] [6]), .ZN(n_8_0_6249));
   NAND2_X1 i_8_0_7523 (.A1(n_8_0_6663), .A2(n_8_0_6668), .ZN(n_8_0_6593));
   NAND2_X1 i_8_0_7524 (.A1(n_8_0_6813), .A2(n_8_0_6671), .ZN(n_8_0_6247));
   AOI21_X1 i_8_0_7525 (.A(n_8_0_30), .B1(n_8_0_7336), .B2(n_8_0_7335), .ZN(
      n_8_0_7334));
   NAND2_X1 i_8_0_7526 (.A1(n_8_0_6438), .A2(n_8_0_6668), .ZN(n_8_0_7335));
   INV_X1 i_8_0_7527 (.A(n_8_0_6594), .ZN(n_8_0_7336));
   OAI211_X1 i_8_0_7528 (.A(n_8_0_6525), .B(n_8_0_5431), .C1(n_8_0_6265), 
      .C2(n_8_0_93), .ZN(n_8_0_5430));
   OAI221_X1 i_8_0_7529 (.A(n_8_0_7341), .B1(n_8_0_7340), .B2(n_8_0_7339), 
      .C1(n_8_0_7338), .C2(n_8_0_7342), .ZN(n_8_0_7337));
   INV_X1 i_8_0_7530 (.A(n_8_0_5424), .ZN(n_8_0_7338));
   INV_X1 i_8_0_7531 (.A(n_8_0_6610), .ZN(n_8_0_7339));
   INV_X1 i_8_0_7532 (.A(n_8_0_5426), .ZN(n_8_0_7340));
   INV_X1 i_8_0_7533 (.A(n_8_0_5428), .ZN(n_8_0_7341));
   INV_X1 i_8_0_7534 (.A(n_8_0_156), .ZN(n_8_0_7342));
   AOI21_X1 i_8_0_7535 (.A(n_8_0_5415), .B1(n_8_0_6838), .B2(n_8_0_6926), 
      .ZN(n_8_0_5414));
   AOI21_X1 i_8_0_7536 (.A(n_8_0_5440), .B1(n_8_0_282), .B2(n_8_0_5439), 
      .ZN(n_8_0_5438));
   NAND2_X1 i_8_0_7537 (.A1(n_8_0_5417), .A2(n_8_0_6511), .ZN(n_8_0_5416));
   OAI21_X1 i_8_0_7538 (.A(n_8_0_5455), .B1(n_8_0_5421), .B2(n_8_0_5422), 
      .ZN(n_8_0_5420));
   NAND2_X1 i_8_0_7539 (.A1(n_8_0_6233), .A2(n_8_0_5436), .ZN(n_8_0_7343));
   OAI211_X1 i_8_0_7540 (.A(n_8_0_471), .B(n_8_0_6727), .C1(n_8_0_6543), 
      .C2(n_8_0_6724), .ZN(n_8_0_5436));
   NAND2_X1 i_8_0_7541 (.A1(\out_bs[7] [2]), .A2(\out_bs[7] [1]), .ZN(n_8_0_6724));
   NAND2_X1 i_8_0_7542 (.A1(\out_bs[7] [6]), .A2(\out_bs[7] [5]), .ZN(n_8_0_6727));
   INV_X1 i_8_0_7543 (.A(n_8_0_6232), .ZN(n_8_0_6233));
   NAND2_X1 i_8_0_7544 (.A1(n_8_0_6731), .A2(n_8_0_6854), .ZN(n_8_0_6232));
   INV_X1 i_8_0_7545 (.A(n_8_0_7344), .ZN(n_250));
   OAI21_X1 i_8_0_7546 (.A(n_8_0_6854), .B1(n_8_0_7350), .B2(n_8_0_7345), 
      .ZN(n_8_0_7344));
   NAND4_X1 i_8_0_7547 (.A1(n_8_0_7349), .A2(n_8_0_6002), .A3(n_8_0_7348), 
      .A4(n_8_0_7346), .ZN(n_8_0_7345));
   NOR2_X1 i_8_0_7548 (.A1(n_8_0_5985), .A2(n_8_0_7347), .ZN(n_8_0_7346));
   NAND2_X1 i_8_0_7549 (.A1(n_8_0_5977), .A2(n_8_0_5997), .ZN(n_8_0_7347));
   AOI21_X1 i_8_0_7550 (.A(n_8_0_5986), .B1(n_8_0_173), .B2(n_8_0_6772), 
      .ZN(n_8_0_5985));
   INV_X1 i_8_0_7551 (.A(n_8_0_5993), .ZN(n_8_0_7348));
   OAI21_X1 i_8_0_7552 (.A(n_8_0_5994), .B1(n_8_0_299), .B2(n_8_0_6795), 
      .ZN(n_8_0_5993));
   OAI21_X1 i_8_0_7553 (.A(n_8_0_5965), .B1(\out_bs[5] [4]), .B2(n_8_0_5966), 
      .ZN(n_8_0_7349));
   OR2_X1 i_8_0_7554 (.A1(n_8_0_7354), .A2(n_8_0_7351), .ZN(n_8_0_7350));
   OAI21_X1 i_8_0_7555 (.A(n_8_0_7352), .B1(n_8_0_425), .B2(n_8_0_6755), 
      .ZN(n_8_0_7351));
   OAI211_X1 i_8_0_7556 (.A(n_8_0_5969), .B(n_8_0_7353), .C1(n_8_0_6759), 
      .C2(n_8_0_6879), .ZN(n_8_0_7352));
   INV_X1 i_8_0_7557 (.A(n_8_0_6752), .ZN(n_8_0_7353));
   NAND2_X1 i_8_0_7558 (.A1(\out_bs[6] [6]), .A2(\out_bs[6] [5]), .ZN(n_8_0_6752));
   OAI21_X1 i_8_0_7559 (.A(n_8_0_7357), .B1(n_8_0_6730), .B2(n_8_0_7355), 
      .ZN(n_8_0_7354));
   INV_X1 i_8_0_7560 (.A(n_8_0_7356), .ZN(n_8_0_7355));
   NAND2_X1 i_8_0_7561 (.A1(n_8_0_7358), .A2(n_8_0_488), .ZN(n_8_0_7356));
   OR2_X1 i_8_0_7562 (.A1(n_8_0_7358), .A2(n_8_0_488), .ZN(n_8_0_7357));
   NAND3_X1 i_8_0_7563 (.A1(\out_bs[7] [6]), .A2(\out_bs[7] [5]), .A3(n_8_0_5973), 
      .ZN(n_8_0_7358));
   INV_X1 i_8_0_7564 (.A(n_8_0_7359), .ZN(n_8_0_5973));
   AOI21_X1 i_8_0_7565 (.A(\out_bs[7] [4]), .B1(n_8_0_6726), .B2(n_8_0_7433), 
      .ZN(n_8_0_7359));
   AOI21_X1 i_8_0_7566 (.A(n_8_0_6853), .B1(n_8_0_6115), .B2(n_8_0_7360), 
      .ZN(n_251));
   INV_X1 i_8_0_7567 (.A(n_8_0_7361), .ZN(n_8_0_7360));
   NAND4_X1 i_8_0_7568 (.A1(n_8_0_6120), .A2(n_8_0_6132), .A3(n_8_0_6110), 
      .A4(n_8_0_7362), .ZN(n_8_0_7361));
   INV_X1 i_8_0_7569 (.A(n_8_0_7363), .ZN(n_8_0_7362));
   OR4_X1 i_8_0_7570 (.A1(n_8_0_6105), .A2(n_8_0_6129), .A3(n_8_0_7367), 
      .A4(n_8_0_7364), .ZN(n_8_0_7363));
   AOI21_X1 i_8_0_7571 (.A(n_8_0_6595), .B1(n_8_0_7366), .B2(n_8_0_7365), 
      .ZN(n_8_0_7364));
   NAND2_X1 i_8_0_7572 (.A1(n_8_0_6248), .A2(n_8_0_6140), .ZN(n_8_0_7365));
   NOR2_X1 i_8_0_7573 (.A1(n_8_0_6810), .A2(n_8_0_6671), .ZN(n_8_0_6595));
   INV_X1 i_8_0_7574 (.A(n_8_0_6138), .ZN(n_8_0_7366));
   INV_X1 i_8_0_7575 (.A(n_8_0_6124), .ZN(n_8_0_7367));
   OAI21_X1 i_8_0_7576 (.A(n_8_0_6125), .B1(n_8_0_6783), .B2(n_8_0_6966), 
      .ZN(n_8_0_6124));
   INV_X1 i_8_0_7577 (.A(n_8_0_7368), .ZN(n_8_0_6129));
   OAI21_X1 i_8_0_7578 (.A(n_8_0_7369), .B1(n_8_0_7371), .B2(n_8_0_7370), 
      .ZN(n_8_0_7368));
   INV_X1 i_8_0_7579 (.A(n_8_0_6130), .ZN(n_8_0_7369));
   INV_X1 i_8_0_7580 (.A(n_8_0_6772), .ZN(n_8_0_7370));
   INV_X1 i_8_0_7581 (.A(n_8_0_177), .ZN(n_8_0_7371));
   OAI21_X1 i_8_0_7582 (.A(n_8_0_6106), .B1(n_8_0_6837), .B2(n_8_0_240), 
      .ZN(n_8_0_6105));
   NAND2_X1 i_8_0_7583 (.A1(n_8_0_6111), .A2(n_8_0_6112), .ZN(n_8_0_6110));
   AOI21_X1 i_8_0_7584 (.A(n_8_0_7372), .B1(n_8_0_7373), .B2(n_8_0_6729), 
      .ZN(n_8_0_6115));
   AOI211_X1 i_8_0_7585 (.A(n_8_0_6715), .B(n_8_0_6117), .C1(n_8_0_6730), 
      .C2(n_8_0_492), .ZN(n_8_0_7372));
   NOR2_X1 i_8_0_7586 (.A1(\out_bs[7] [3]), .A2(n_8_0_6475), .ZN(n_8_0_6117));
   INV_X1 i_8_0_7587 (.A(n_8_0_492), .ZN(n_8_0_7373));
   AOI21_X1 i_8_0_7588 (.A(n_8_0_6853), .B1(n_8_0_6199), .B2(n_8_0_7374), 
      .ZN(n_252));
   INV_X1 i_8_0_7589 (.A(n_8_0_7375), .ZN(n_8_0_7374));
   OR4_X1 i_8_0_7590 (.A1(n_8_0_6193), .A2(n_8_0_6207), .A3(n_8_0_6186), 
      .A4(n_8_0_7376), .ZN(n_8_0_7375));
   NAND4_X1 i_8_0_7591 (.A1(n_8_0_6212), .A2(n_8_0_6179), .A3(n_8_0_6203), 
      .A4(n_8_0_7377), .ZN(n_8_0_7376));
   AOI21_X1 i_8_0_7592 (.A(n_8_0_6183), .B1(n_8_0_6185), .B2(n_8_0_6248), 
      .ZN(n_8_0_7377));
   NAND2_X1 i_8_0_7593 (.A1(n_8_0_6204), .A2(n_8_0_6205), .ZN(n_8_0_6203));
   OAI21_X1 i_8_0_7594 (.A(n_8_0_6180), .B1(n_8_0_6773), .B2(n_8_0_6943), 
      .ZN(n_8_0_6179));
   NAND2_X1 i_8_0_7595 (.A1(n_8_0_6213), .A2(n_8_0_6214), .ZN(n_8_0_6212));
   INV_X1 i_8_0_7596 (.A(n_8_0_7378), .ZN(n_8_0_6186));
   NAND2_X1 i_8_0_7597 (.A1(n_8_0_6187), .A2(n_8_0_6188), .ZN(n_8_0_7378));
   OAI21_X1 i_8_0_7598 (.A(n_8_0_6208), .B1(n_8_0_6824), .B2(n_8_0_368), 
      .ZN(n_8_0_6207));
   OAI21_X1 i_8_0_7599 (.A(n_8_0_6194), .B1(n_8_0_431), .B2(n_8_0_6755), 
      .ZN(n_8_0_6193));
   AOI21_X1 i_8_0_7600 (.A(n_8_0_7379), .B1(n_8_0_7382), .B2(n_8_0_6729), 
      .ZN(n_8_0_6199));
   AOI211_X1 i_8_0_7601 (.A(n_8_0_6715), .B(n_8_0_7380), .C1(n_8_0_6730), 
      .C2(n_8_0_494), .ZN(n_8_0_7379));
   AOI21_X1 i_8_0_7602 (.A(\out_bs[7] [3]), .B1(\out_bs[7] [2]), .B2(n_8_0_7381), 
      .ZN(n_8_0_7380));
   INV_X1 i_8_0_7603 (.A(n_8_0_6544), .ZN(n_8_0_7381));
   INV_X1 i_8_0_7604 (.A(n_8_0_6730), .ZN(n_8_0_6729));
   INV_X1 i_8_0_7605 (.A(n_8_0_494), .ZN(n_8_0_7382));
   INV_X1 i_8_0_7606 (.A(n_8_0_7383), .ZN(n_253));
   OAI21_X1 i_8_0_7607 (.A(n_8_0_6854), .B1(n_8_0_7396), .B2(n_8_0_7384), 
      .ZN(n_8_0_7383));
   NAND2_X1 i_8_0_7608 (.A1(n_8_0_6289), .A2(n_8_0_7385), .ZN(n_8_0_7384));
   INV_X1 i_8_0_7609 (.A(n_8_0_7386), .ZN(n_8_0_7385));
   OR2_X1 i_8_0_7610 (.A1(n_8_0_6296), .A2(n_8_0_7387), .ZN(n_8_0_7386));
   NAND4_X1 i_8_0_7611 (.A1(n_8_0_6272), .A2(n_8_0_6302), .A3(n_8_0_6280), 
      .A4(n_8_0_7388), .ZN(n_8_0_7387));
   INV_X1 i_8_0_7612 (.A(n_8_0_7389), .ZN(n_8_0_7388));
   OAI211_X1 i_8_0_7613 (.A(n_8_0_6263), .B(n_8_0_7390), .C1(n_8_0_55), .C2(
      n_8_0_6811), .ZN(n_8_0_7389));
   NAND2_X1 i_8_0_7614 (.A1(n_8_0_7392), .A2(n_8_0_7391), .ZN(n_8_0_7390));
   NOR2_X1 i_8_0_7615 (.A1(n_8_0_6261), .A2(n_8_0_6670), .ZN(n_8_0_7391));
   NAND2_X1 i_8_0_7616 (.A1(n_8_0_6812), .A2(n_8_0_55), .ZN(n_8_0_7392));
   INV_X1 i_8_0_7617 (.A(n_8_0_7393), .ZN(n_8_0_6811));
   NAND2_X1 i_8_0_7618 (.A1(n_8_0_7394), .A2(n_8_0_7395), .ZN(n_8_0_7393));
   INV_X1 i_8_0_7619 (.A(n_8_0_6813), .ZN(n_8_0_7394));
   INV_X1 i_8_0_7620 (.A(n_8_0_6814), .ZN(n_8_0_7395));
   NAND2_X1 i_8_0_7621 (.A1(n_8_0_6281), .A2(n_8_0_6284), .ZN(n_8_0_6280));
   AOI22_X1 i_8_0_7622 (.A1(n_8_0_6303), .A2(n_8_0_6304), .B1(n_8_0_6648), 
      .B2(n_8_0_6576), .ZN(n_8_0_6302));
   AOI22_X1 i_8_0_7623 (.A1(n_8_0_6794), .A2(n_8_0_6909), .B1(n_8_0_6636), 
      .B2(n_8_0_6273), .ZN(n_8_0_6272));
   OAI22_X1 i_8_0_7624 (.A1(n_8_0_6297), .A2(n_8_0_370), .B1(n_8_0_6298), 
      .B2(n_8_0_6509), .ZN(n_8_0_6296));
   AOI22_X1 i_8_0_7625 (.A1(n_8_0_6754), .A2(n_8_0_6877), .B1(n_8_0_6753), 
      .B2(n_8_0_6290), .ZN(n_8_0_6289));
   OAI21_X1 i_8_0_7626 (.A(n_8_0_7399), .B1(n_8_0_6730), .B2(n_8_0_7397), 
      .ZN(n_8_0_7396));
   INV_X1 i_8_0_7627 (.A(n_8_0_7398), .ZN(n_8_0_7397));
   NAND2_X1 i_8_0_7628 (.A1(n_8_0_7400), .A2(n_8_0_496), .ZN(n_8_0_7398));
   OR2_X1 i_8_0_7629 (.A1(n_8_0_7400), .A2(n_8_0_496), .ZN(n_8_0_7399));
   OR2_X1 i_8_0_7630 (.A1(n_8_0_6715), .A2(n_8_0_6279), .ZN(n_8_0_7400));
   NOR2_X1 i_8_0_7631 (.A1(n_8_0_6723), .A2(\out_bs[7] [3]), .ZN(n_8_0_6279));
   AOI21_X1 i_8_0_7632 (.A(n_8_0_6853), .B1(n_8_0_6401), .B2(n_8_0_7401), 
      .ZN(n_254));
   NOR4_X1 i_8_0_7633 (.A1(n_8_0_6383), .A2(n_8_0_7413), .A3(n_8_0_6378), 
      .A4(n_8_0_7402), .ZN(n_8_0_7401));
   NAND4_X1 i_8_0_7634 (.A1(n_8_0_7407), .A2(n_8_0_6396), .A3(n_8_0_7406), 
      .A4(n_8_0_6389), .ZN(n_8_0_7402));
   INV_X1 i_8_0_7635 (.A(n_8_0_7403), .ZN(n_8_0_6389));
   NAND2_X1 i_8_0_7636 (.A1(n_8_0_7404), .A2(n_8_0_7405), .ZN(n_8_0_7403));
   NAND2_X1 i_8_0_7637 (.A1(n_8_0_6391), .A2(n_8_0_6691), .ZN(n_8_0_7404));
   INV_X1 i_8_0_7638 (.A(n_8_0_6390), .ZN(n_8_0_7405));
   NAND2_X1 i_8_0_7639 (.A1(n_8_0_6416), .A2(n_8_0_6418), .ZN(n_8_0_7406));
   OAI21_X1 i_8_0_7640 (.A(n_8_0_6397), .B1(n_8_0_6773), .B2(n_8_0_6940), 
      .ZN(n_8_0_6396));
   OR2_X1 i_8_0_7641 (.A1(n_8_0_7408), .A2(n_8_0_6411), .ZN(n_8_0_7407));
   INV_X1 i_8_0_7642 (.A(n_8_0_7409), .ZN(n_8_0_7408));
   NAND2_X1 i_8_0_7643 (.A1(n_8_0_6837), .A2(n_8_0_247), .ZN(n_8_0_7409));
   INV_X1 i_8_0_7644 (.A(n_8_0_7410), .ZN(n_8_0_6378));
   NAND2_X1 i_8_0_7645 (.A1(n_8_0_7411), .A2(n_8_0_7412), .ZN(n_8_0_7410));
   NAND2_X1 i_8_0_7646 (.A1(n_8_0_6795), .A2(n_8_0_310), .ZN(n_8_0_7411));
   INV_X1 i_8_0_7647 (.A(n_8_0_6379), .ZN(n_8_0_7412));
   INV_X1 i_8_0_7648 (.A(n_8_0_6406), .ZN(n_8_0_7413));
   OAI21_X1 i_8_0_7649 (.A(n_8_0_6407), .B1(n_8_0_6825), .B2(n_8_0_6896), 
      .ZN(n_8_0_6406));
   AOI221_X1 i_8_0_7650 (.A(n_8_0_6584), .B1(n_8_0_436), .B2(n_8_0_6384), 
      .C1(n_8_0_6387), .C2(n_8_0_6755), .ZN(n_8_0_6383));
   NAND2_X1 i_8_0_7651 (.A1(n_8_0_7415), .A2(n_8_0_7414), .ZN(n_8_0_6401));
   NAND2_X1 i_8_0_7652 (.A1(n_8_0_7416), .A2(n_8_0_499), .ZN(n_8_0_7414));
   OAI21_X1 i_8_0_7653 (.A(n_8_0_6730), .B1(n_8_0_499), .B2(n_8_0_7416), 
      .ZN(n_8_0_7415));
   OR2_X1 i_8_0_7654 (.A1(n_8_0_6715), .A2(n_8_0_6403), .ZN(n_8_0_7416));
   OAI21_X1 i_8_0_7655 (.A(\out_bs[7] [3]), .B1(\out_bs[7] [2]), .B2(
      \out_bs[7] [1]), .ZN(n_8_0_6403));
   NAND2_X1 i_8_0_7656 (.A1(n_8_0_6728), .A2(\out_bs[7] [4]), .ZN(n_8_0_6715));
   INV_X1 i_8_0_7657 (.A(n_8_0_7417), .ZN(n_255));
   OAI21_X1 i_8_0_7658 (.A(n_8_0_6854), .B1(n_8_0_6614), .B2(n_8_0_7418), 
      .ZN(n_8_0_7417));
   OR4_X1 i_8_0_7659 (.A1(n_8_0_6620), .A2(n_8_0_6582), .A3(n_8_0_6569), 
      .A4(n_8_0_7419), .ZN(n_8_0_7418));
   OR2_X1 i_8_0_7660 (.A1(n_8_0_6602), .A2(n_8_0_6592), .ZN(n_8_0_7419));
   OAI22_X1 i_8_0_7661 (.A1(n_8_0_6603), .A2(n_8_0_188), .B1(n_8_0_6604), 
      .B2(n_8_0_6610), .ZN(n_8_0_6602));
   AOI221_X1 i_8_0_7662 (.A(n_8_0_6584), .B1(n_8_0_440), .B2(n_8_0_6585), 
      .C1(n_8_0_6743), .C2(n_8_0_6755), .ZN(n_8_0_6582));
   NOR2_X1 i_8_0_7663 (.A1(n_8_0_6759), .A2(n_8_0_6757), .ZN(n_8_0_6755));
   OAI21_X1 i_8_0_7664 (.A(n_8_0_7430), .B1(n_8_0_6730), .B2(n_8_0_7420), 
      .ZN(n_8_0_6614));
   AOI21_X1 i_8_0_7665 (.A(n_8_0_7435), .B1(n_8_0_6728), .B2(n_8_0_7431), 
      .ZN(n_8_0_7420));
   NOR2_X1 i_8_0_7666 (.A1(n_8_0_6731), .A2(n_8_0_6853), .ZN(n_8_0_6730));
   INV_X1 i_8_0_7667 (.A(n_8_0_7421), .ZN(n_8_0_6731));
   OAI21_X1 i_8_0_7668 (.A(n_8_0_7422), .B1(\out_as[7] [6]), .B2(n_8_0_7000), 
      .ZN(n_8_0_7421));
   NAND2_X1 i_8_0_7669 (.A1(n_8_0_7424), .A2(n_8_0_7423), .ZN(n_8_0_7422));
   AOI22_X1 i_8_0_7670 (.A1(n_8_0_7000), .A2(\out_as[7] [6]), .B1(\out_as[7] [5]), 
      .B2(n_8_0_6999), .ZN(n_8_0_7423));
   OAI221_X1 i_8_0_7671 (.A(n_8_0_7425), .B1(\out_as[7] [5]), .B2(n_8_0_6999), 
      .C1(\out_as[7] [4]), .C2(n_8_0_6998), .ZN(n_8_0_7424));
   OAI221_X1 i_8_0_7672 (.A(n_8_0_7426), .B1(n_8_0_7004), .B2(\out_bs[7] [4]), 
      .C1(n_8_0_7003), .C2(\out_bs[7] [3]), .ZN(n_8_0_7425));
   OAI21_X1 i_8_0_7673 (.A(n_8_0_7427), .B1(\out_as[7] [3]), .B2(n_8_0_6997), 
      .ZN(n_8_0_7426));
   AOI21_X1 i_8_0_7674 (.A(n_8_0_7428), .B1(n_8_0_7429), .B2(\out_bs[7] [2]), 
      .ZN(n_8_0_7427));
   AOI221_X1 i_8_0_7675 (.A(n_8_0_3711), .B1(\out_as[7] [1]), .B2(n_8_0_3756), 
      .C1(n_8_0_6996), .C2(\out_as[7] [2]), .ZN(n_8_0_7428));
   INV_X1 i_8_0_7676 (.A(\out_bs[7] [2]), .ZN(n_8_0_6996));
   INV_X1 i_8_0_7677 (.A(\out_as[7] [2]), .ZN(n_8_0_7429));
   INV_X1 i_8_0_7678 (.A(\out_bs[7] [3]), .ZN(n_8_0_6997));
   INV_X1 i_8_0_7679 (.A(\out_as[7] [3]), .ZN(n_8_0_7003));
   INV_X1 i_8_0_7680 (.A(\out_as[7] [4]), .ZN(n_8_0_7004));
   INV_X1 i_8_0_7681 (.A(\out_bs[7] [4]), .ZN(n_8_0_6998));
   INV_X1 i_8_0_7682 (.A(\out_bs[7] [5]), .ZN(n_8_0_6999));
   INV_X1 i_8_0_7683 (.A(\out_bs[7] [6]), .ZN(n_8_0_7000));
   NAND3_X1 i_8_0_7684 (.A1(n_8_0_6728), .A2(n_8_0_7435), .A3(n_8_0_7431), 
      .ZN(n_8_0_7430));
   INV_X1 i_8_0_7685 (.A(n_8_0_7432), .ZN(n_8_0_7431));
   NAND3_X1 i_8_0_7686 (.A1(\out_bs[7] [4]), .A2(\out_bs[7] [1]), .A3(n_8_0_7433), 
      .ZN(n_8_0_7432));
   INV_X1 i_8_0_7687 (.A(n_8_0_7434), .ZN(n_8_0_7433));
   NAND2_X1 i_8_0_7688 (.A1(\out_bs[7] [3]), .A2(\out_bs[7] [2]), .ZN(n_8_0_7434));
   INV_X1 i_8_0_7689 (.A(n_8_0_503), .ZN(n_8_0_7435));
   INV_X1 i_8_0_7690 (.A(n_8_0_6853), .ZN(n_8_0_6854));
   NAND2_X1 i_8_0_7691 (.A1(enbl_in), .A2(n_8_0_7436), .ZN(n_8_0_6853));
   INV_X1 i_8_0_7692 (.A(rst), .ZN(n_8_0_7436));
   DFFS_X1 error_success_reg (.D(n_0_164), .SN(n_0_169), .CK(clk), .Q(
      error_success), .QN());
   CLKGATETST_X1 clk_gate_out_data_reg (.CK(clk), .E(n_0_40), .SE(1'b0), 
      .GCK(n_0_39));
   DFF_X1 \out_data_reg[31]  (.D(n_0_38), .CK(n_0_39), .Q(out_data[31]), .QN());
   DFF_X1 \out_data_reg[30]  (.D(n_0_37), .CK(n_0_39), .Q(out_data[30]), .QN());
   DFF_X1 \out_data_reg[29]  (.D(n_0_36), .CK(n_0_39), .Q(out_data[29]), .QN());
   DFF_X1 \out_data_reg[28]  (.D(n_0_35), .CK(n_0_39), .Q(out_data[28]), .QN());
   DFF_X1 \out_data_reg[27]  (.D(n_0_34), .CK(n_0_39), .Q(out_data[27]), .QN());
   DFF_X1 \out_data_reg[26]  (.D(n_0_33), .CK(n_0_39), .Q(out_data[26]), .QN());
   DFF_X1 \out_data_reg[25]  (.D(n_0_32), .CK(n_0_39), .Q(out_data[25]), .QN());
   DFF_X1 \out_data_reg[24]  (.D(n_0_31), .CK(n_0_39), .Q(out_data[24]), .QN());
   DFF_X1 \out_data_reg[23]  (.D(n_0_30), .CK(n_0_39), .Q(out_data[23]), .QN());
   DFF_X1 \out_data_reg[22]  (.D(n_0_29), .CK(n_0_39), .Q(out_data[22]), .QN());
   DFF_X1 \out_data_reg[21]  (.D(n_0_28), .CK(n_0_39), .Q(out_data[21]), .QN());
   DFF_X1 \out_data_reg[20]  (.D(n_0_27), .CK(n_0_39), .Q(out_data[20]), .QN());
   DFF_X1 \out_data_reg[19]  (.D(n_0_26), .CK(n_0_39), .Q(out_data[19]), .QN());
   DFF_X1 \out_data_reg[18]  (.D(n_0_25), .CK(n_0_39), .Q(out_data[18]), .QN());
   DFF_X1 \out_data_reg[17]  (.D(n_0_24), .CK(n_0_39), .Q(out_data[17]), .QN());
   DFF_X1 \out_data_reg[16]  (.D(n_0_23), .CK(n_0_39), .Q(out_data[16]), .QN());
   DFF_X1 \out_data_reg[15]  (.D(n_0_22), .CK(n_0_39), .Q(out_data[15]), .QN());
   DFF_X1 \out_data_reg[14]  (.D(n_0_21), .CK(n_0_39), .Q(out_data[14]), .QN());
   DFF_X1 \out_data_reg[13]  (.D(n_0_20), .CK(n_0_39), .Q(out_data[13]), .QN());
   DFF_X1 \out_data_reg[12]  (.D(n_0_19), .CK(n_0_39), .Q(out_data[12]), .QN());
   DFF_X1 \out_data_reg[11]  (.D(n_0_18), .CK(n_0_39), .Q(out_data[11]), .QN());
   DFF_X1 \out_data_reg[10]  (.D(n_0_17), .CK(n_0_39), .Q(out_data[10]), .QN());
   DFF_X1 \out_data_reg[9]  (.D(n_0_16), .CK(n_0_39), .Q(out_data[9]), .QN());
   DFF_X1 \out_data_reg[8]  (.D(n_0_15), .CK(n_0_39), .Q(out_data[8]), .QN());
   DFF_X1 \out_data_reg[7]  (.D(n_0_14), .CK(n_0_39), .Q(out_data[7]), .QN());
   DFF_X1 \out_data_reg[6]  (.D(n_0_13), .CK(n_0_39), .Q(out_data[6]), .QN());
   DFF_X1 \out_data_reg[5]  (.D(n_0_12), .CK(n_0_39), .Q(out_data[5]), .QN());
   DFF_X1 \out_data_reg[4]  (.D(n_0_11), .CK(n_0_39), .Q(out_data[4]), .QN());
   DFF_X1 \out_data_reg[3]  (.D(n_0_10), .CK(n_0_39), .Q(out_data[3]), .QN());
   DFF_X1 \out_data_reg[2]  (.D(n_0_9), .CK(n_0_39), .Q(out_data[2]), .QN());
   DFF_X1 \out_data_reg[1]  (.D(n_0_8), .CK(n_0_39), .Q(out_data[1]), .QN());
   DFF_X1 \out_data_reg[0]  (.D(n_0_7), .CK(n_0_39), .Q(out_data[0]), .QN());
   DFF_X1 \buf_reg[127]  (.D(n_0_295), .CK(clk), .Q(n_0_0), .QN());
   DFF_X1 \buf_reg[126]  (.D(n_0_294), .CK(clk), .Q(n_0_1), .QN());
   DFF_X1 \buf_reg[125]  (.D(n_0_293), .CK(clk), .Q(n_0_2), .QN());
   DFF_X1 \buf_reg[124]  (.D(n_0_292), .CK(clk), .Q(n_0_3), .QN());
   DFF_X1 \buf_reg[123]  (.D(n_0_291), .CK(clk), .Q(n_0_4), .QN());
   DFF_X1 \buf_reg[122]  (.D(n_0_290), .CK(clk), .Q(n_0_6), .QN());
   DFF_X1 \buf_reg[121]  (.D(n_0_289), .CK(clk), .Q(n_0_41), .QN());
   DFF_X1 \buf_reg[120]  (.D(n_0_288), .CK(clk), .Q(n_0_42), .QN());
   DFF_X1 \buf_reg[119]  (.D(n_0_287), .CK(clk), .Q(n_0_43), .QN());
   DFF_X1 \buf_reg[118]  (.D(n_0_286), .CK(clk), .Q(n_0_44), .QN());
   DFF_X1 \buf_reg[117]  (.D(n_0_285), .CK(clk), .Q(n_0_45), .QN());
   DFF_X1 \buf_reg[116]  (.D(n_0_284), .CK(clk), .Q(n_0_46), .QN());
   DFF_X1 \buf_reg[115]  (.D(n_0_283), .CK(clk), .Q(n_0_47), .QN());
   DFF_X1 \buf_reg[114]  (.D(n_0_282), .CK(clk), .Q(n_0_48), .QN());
   DFF_X1 \buf_reg[113]  (.D(n_0_281), .CK(clk), .Q(n_0_49), .QN());
   DFF_X1 \buf_reg[112]  (.D(n_0_280), .CK(clk), .Q(n_0_50), .QN());
   DFF_X1 \buf_reg[111]  (.D(n_0_279), .CK(clk), .Q(n_0_51), .QN());
   DFF_X1 \buf_reg[110]  (.D(n_0_278), .CK(clk), .Q(n_0_52), .QN());
   DFF_X1 \buf_reg[109]  (.D(n_0_277), .CK(clk), .Q(n_0_53), .QN());
   DFF_X1 \buf_reg[108]  (.D(n_0_276), .CK(clk), .Q(n_0_54), .QN());
   DFF_X1 \buf_reg[107]  (.D(n_0_275), .CK(clk), .Q(n_0_55), .QN());
   DFF_X1 \buf_reg[106]  (.D(n_0_274), .CK(clk), .Q(n_0_56), .QN());
   DFF_X1 \buf_reg[105]  (.D(n_0_273), .CK(clk), .Q(n_0_57), .QN());
   DFF_X1 \buf_reg[104]  (.D(n_0_272), .CK(clk), .Q(n_0_58), .QN());
   DFF_X1 \buf_reg[103]  (.D(n_0_271), .CK(clk), .Q(n_0_59), .QN());
   DFF_X1 \buf_reg[102]  (.D(n_0_270), .CK(clk), .Q(n_0_60), .QN());
   DFF_X1 \buf_reg[101]  (.D(n_0_269), .CK(clk), .Q(n_0_61), .QN());
   DFF_X1 \buf_reg[100]  (.D(n_0_268), .CK(clk), .Q(n_0_62), .QN());
   DFF_X1 \buf_reg[99]  (.D(n_0_267), .CK(clk), .Q(n_0_63), .QN());
   DFF_X1 \buf_reg[98]  (.D(n_0_266), .CK(clk), .Q(n_0_64), .QN());
   DFF_X1 \buf_reg[97]  (.D(n_0_265), .CK(clk), .Q(n_0_65), .QN());
   DFF_X1 \buf_reg[96]  (.D(n_0_264), .CK(clk), .Q(n_0_66), .QN());
   DFF_X1 \buf_reg[95]  (.D(n_0_263), .CK(clk), .Q(n_0_67), .QN());
   DFF_X1 \buf_reg[94]  (.D(n_0_262), .CK(clk), .Q(n_0_68), .QN());
   DFF_X1 \buf_reg[93]  (.D(n_0_261), .CK(clk), .Q(n_0_69), .QN());
   DFF_X1 \buf_reg[92]  (.D(n_0_260), .CK(clk), .Q(n_0_70), .QN());
   DFF_X1 \buf_reg[91]  (.D(n_0_259), .CK(clk), .Q(n_0_71), .QN());
   DFF_X1 \buf_reg[90]  (.D(n_0_258), .CK(clk), .Q(n_0_72), .QN());
   DFF_X1 \buf_reg[89]  (.D(n_0_257), .CK(clk), .Q(n_0_73), .QN());
   DFF_X1 \buf_reg[88]  (.D(n_0_256), .CK(clk), .Q(n_0_74), .QN());
   DFF_X1 \buf_reg[87]  (.D(n_0_255), .CK(clk), .Q(n_0_75), .QN());
   DFF_X1 \buf_reg[86]  (.D(n_0_254), .CK(clk), .Q(n_0_76), .QN());
   DFF_X1 \buf_reg[85]  (.D(n_0_253), .CK(clk), .Q(n_0_77), .QN());
   DFF_X1 \buf_reg[84]  (.D(n_0_252), .CK(clk), .Q(n_0_78), .QN());
   DFF_X1 \buf_reg[83]  (.D(n_0_251), .CK(clk), .Q(n_0_79), .QN());
   DFF_X1 \buf_reg[82]  (.D(n_0_250), .CK(clk), .Q(n_0_80), .QN());
   DFF_X1 \buf_reg[81]  (.D(n_0_249), .CK(clk), .Q(n_0_81), .QN());
   DFF_X1 \buf_reg[80]  (.D(n_0_248), .CK(clk), .Q(n_0_82), .QN());
   DFF_X1 \buf_reg[79]  (.D(n_0_247), .CK(clk), .Q(n_0_83), .QN());
   DFF_X1 \buf_reg[78]  (.D(n_0_246), .CK(clk), .Q(n_0_84), .QN());
   DFF_X1 \buf_reg[77]  (.D(n_0_245), .CK(clk), .Q(n_0_85), .QN());
   DFF_X1 \buf_reg[76]  (.D(n_0_244), .CK(clk), .Q(n_0_86), .QN());
   DFF_X1 \buf_reg[75]  (.D(n_0_243), .CK(clk), .Q(n_0_87), .QN());
   DFF_X1 \buf_reg[74]  (.D(n_0_242), .CK(clk), .Q(n_0_88), .QN());
   DFF_X1 \buf_reg[73]  (.D(n_0_241), .CK(clk), .Q(n_0_89), .QN());
   DFF_X1 \buf_reg[72]  (.D(n_0_240), .CK(clk), .Q(n_0_90), .QN());
   DFF_X1 \buf_reg[71]  (.D(n_0_239), .CK(clk), .Q(n_0_91), .QN());
   DFF_X1 \buf_reg[70]  (.D(n_0_238), .CK(clk), .Q(n_0_92), .QN());
   DFF_X1 \buf_reg[69]  (.D(n_0_237), .CK(clk), .Q(n_0_93), .QN());
   DFF_X1 \buf_reg[68]  (.D(n_0_236), .CK(clk), .Q(n_0_94), .QN());
   DFF_X1 \buf_reg[67]  (.D(n_0_235), .CK(clk), .Q(n_0_95), .QN());
   DFF_X1 \buf_reg[66]  (.D(n_0_234), .CK(clk), .Q(n_0_96), .QN());
   DFF_X1 \buf_reg[65]  (.D(n_0_233), .CK(clk), .Q(n_0_97), .QN());
   DFF_X1 \buf_reg[64]  (.D(n_0_232), .CK(clk), .Q(n_0_98), .QN());
   DFF_X1 \buf_reg[63]  (.D(n_0_231), .CK(clk), .Q(n_0_99), .QN());
   DFF_X1 \buf_reg[62]  (.D(n_0_230), .CK(clk), .Q(n_0_100), .QN());
   DFF_X1 \buf_reg[61]  (.D(n_0_229), .CK(clk), .Q(n_0_101), .QN());
   DFF_X1 \buf_reg[60]  (.D(n_0_228), .CK(clk), .Q(n_0_102), .QN());
   DFF_X1 \buf_reg[59]  (.D(n_0_227), .CK(clk), .Q(n_0_103), .QN());
   DFF_X1 \buf_reg[58]  (.D(n_0_226), .CK(clk), .Q(n_0_104), .QN());
   DFF_X1 \buf_reg[57]  (.D(n_0_225), .CK(clk), .Q(n_0_105), .QN());
   DFF_X1 \buf_reg[56]  (.D(n_0_224), .CK(clk), .Q(n_0_106), .QN());
   DFF_X1 \buf_reg[55]  (.D(n_0_223), .CK(clk), .Q(n_0_107), .QN());
   DFF_X1 \buf_reg[54]  (.D(n_0_222), .CK(clk), .Q(n_0_108), .QN());
   DFF_X1 \buf_reg[53]  (.D(n_0_221), .CK(clk), .Q(n_0_109), .QN());
   DFF_X1 \buf_reg[52]  (.D(n_0_220), .CK(clk), .Q(n_0_110), .QN());
   DFF_X1 \buf_reg[51]  (.D(n_0_219), .CK(clk), .Q(n_0_111), .QN());
   DFF_X1 \buf_reg[50]  (.D(n_0_218), .CK(clk), .Q(n_0_112), .QN());
   DFF_X1 \buf_reg[49]  (.D(n_0_217), .CK(clk), .Q(n_0_113), .QN());
   DFF_X1 \buf_reg[48]  (.D(n_0_216), .CK(clk), .Q(n_0_114), .QN());
   DFF_X1 \buf_reg[47]  (.D(n_0_215), .CK(clk), .Q(n_0_115), .QN());
   DFF_X1 \buf_reg[46]  (.D(n_0_214), .CK(clk), .Q(n_0_116), .QN());
   DFF_X1 \buf_reg[45]  (.D(n_0_213), .CK(clk), .Q(n_0_117), .QN());
   DFF_X1 \buf_reg[44]  (.D(n_0_212), .CK(clk), .Q(n_0_118), .QN());
   DFF_X1 \buf_reg[43]  (.D(n_0_211), .CK(clk), .Q(n_0_119), .QN());
   DFF_X1 \buf_reg[42]  (.D(n_0_210), .CK(clk), .Q(n_0_120), .QN());
   DFF_X1 \buf_reg[41]  (.D(n_0_209), .CK(clk), .Q(n_0_121), .QN());
   DFF_X1 \buf_reg[40]  (.D(n_0_208), .CK(clk), .Q(n_0_122), .QN());
   DFF_X1 \buf_reg[39]  (.D(n_0_207), .CK(clk), .Q(n_0_123), .QN());
   DFF_X1 \buf_reg[38]  (.D(n_0_206), .CK(clk), .Q(n_0_124), .QN());
   DFF_X1 \buf_reg[37]  (.D(n_0_205), .CK(clk), .Q(n_0_125), .QN());
   DFF_X1 \buf_reg[36]  (.D(n_0_204), .CK(clk), .Q(n_0_126), .QN());
   DFF_X1 \buf_reg[35]  (.D(n_0_203), .CK(clk), .Q(n_0_127), .QN());
   DFF_X1 \buf_reg[34]  (.D(n_0_202), .CK(clk), .Q(n_0_128), .QN());
   DFF_X1 \buf_reg[33]  (.D(n_0_201), .CK(clk), .Q(n_0_129), .QN());
   DFF_X1 \buf_reg[32]  (.D(n_0_200), .CK(clk), .Q(n_0_130), .QN());
   DFF_X1 \buf_reg[31]  (.D(n_0_199), .CK(clk), .Q(n_0_131), .QN());
   DFF_X1 \buf_reg[30]  (.D(n_0_198), .CK(clk), .Q(n_0_132), .QN());
   DFF_X1 \buf_reg[29]  (.D(n_0_197), .CK(clk), .Q(n_0_133), .QN());
   DFF_X1 \buf_reg[28]  (.D(n_0_196), .CK(clk), .Q(n_0_134), .QN());
   DFF_X1 \buf_reg[27]  (.D(n_0_195), .CK(clk), .Q(n_0_135), .QN());
   DFF_X1 \buf_reg[26]  (.D(n_0_194), .CK(clk), .Q(n_0_136), .QN());
   DFF_X1 \buf_reg[25]  (.D(n_0_193), .CK(clk), .Q(n_0_137), .QN());
   DFF_X1 \buf_reg[24]  (.D(n_0_192), .CK(clk), .Q(n_0_138), .QN());
   DFF_X1 \buf_reg[23]  (.D(n_0_191), .CK(clk), .Q(n_0_139), .QN());
   DFF_X1 \buf_reg[22]  (.D(n_0_190), .CK(clk), .Q(n_0_140), .QN());
   DFF_X1 \buf_reg[21]  (.D(n_0_189), .CK(clk), .Q(n_0_141), .QN());
   DFF_X1 \buf_reg[20]  (.D(n_0_188), .CK(clk), .Q(n_0_142), .QN());
   DFF_X1 \buf_reg[19]  (.D(n_0_187), .CK(clk), .Q(n_0_143), .QN());
   DFF_X1 \buf_reg[18]  (.D(n_0_186), .CK(clk), .Q(n_0_144), .QN());
   DFF_X1 \buf_reg[17]  (.D(n_0_185), .CK(clk), .Q(n_0_145), .QN());
   DFF_X1 \buf_reg[16]  (.D(n_0_184), .CK(clk), .Q(n_0_146), .QN());
   DFF_X1 \buf_reg[15]  (.D(n_0_183), .CK(clk), .Q(n_0_147), .QN());
   DFF_X1 \buf_reg[14]  (.D(n_0_182), .CK(clk), .Q(n_0_148), .QN());
   DFF_X1 \buf_reg[13]  (.D(n_0_181), .CK(clk), .Q(n_0_149), .QN());
   DFF_X1 \buf_reg[12]  (.D(n_0_180), .CK(clk), .Q(n_0_150), .QN());
   DFF_X1 \buf_reg[11]  (.D(n_0_179), .CK(clk), .Q(n_0_151), .QN());
   DFF_X1 \buf_reg[10]  (.D(n_0_178), .CK(clk), .Q(n_0_152), .QN());
   DFF_X1 \buf_reg[9]  (.D(n_0_177), .CK(clk), .Q(n_0_153), .QN());
   DFF_X1 \buf_reg[8]  (.D(n_0_176), .CK(clk), .Q(n_0_154), .QN());
   DFF_X1 \buf_reg[7]  (.D(n_0_175), .CK(clk), .Q(n_0_155), .QN());
   DFF_X1 \buf_reg[6]  (.D(n_0_174), .CK(clk), .Q(n_0_156), .QN());
   DFF_X1 \buf_reg[5]  (.D(n_0_173), .CK(clk), .Q(n_0_157), .QN());
   DFF_X1 \buf_reg[4]  (.D(n_0_172), .CK(clk), .Q(n_0_158), .QN());
   DFF_X1 \buf_reg[3]  (.D(n_0_168), .CK(clk), .Q(n_0_159), .QN());
   DFF_X1 \buf_reg[2]  (.D(n_0_167), .CK(clk), .Q(n_0_160), .QN());
   DFF_X1 \buf_reg[1]  (.D(n_0_166), .CK(clk), .Q(n_0_161), .QN());
   DFF_X1 \buf_reg[0]  (.D(n_0_165), .CK(clk), .Q(n_0_162), .QN());
   DFFR_X1 out_ready_reg (.D(n_0_5), .RN(n_0_169), .CK(clk), .Q(out_ready), 
      .QN());
   DFFR_X1 \buf_flush_i_reg[5]  (.D(n_0_170), .RN(n_0_169), .CK(clk), .Q(
      buf_flush_i[5]), .QN());
   MUX2_X1 \buf_flush_i_reg[5]_enable_mux_0  (.A(buf_flush_i[5]), .B(
      buf_flush_i_inc[5]), .S(n_0_5), .Z(n_0_170));
   DFFR_X1 \buf_flush_i_reg[6]  (.D(n_0_296), .RN(n_0_169), .CK(clk), .Q(
      buf_flush_i[6]), .QN());
   MUX2_X1 \buf_flush_i_reg[6]_enable_mux_0  (.A(buf_flush_i[6]), .B(
      buf_flush_i_inc[6]), .S(n_0_5), .Z(n_0_296));
   DFFS_X1 \buf_fill_i_reg[6]  (.D(\out_bs[7] [6]), .SN(n_0_169), .CK(n_0_171), 
      .Q(buf_fill_i[6]), .QN());
   DFFS_X1 \buf_fill_i_reg[5]  (.D(\out_bs[7] [5]), .SN(n_0_169), .CK(n_0_171), 
      .Q(buf_fill_i[5]), .QN());
   DFFS_X1 \buf_fill_i_reg[4]  (.D(\out_bs[7] [4]), .SN(n_0_169), .CK(n_0_171), 
      .Q(buf_fill_i[4]), .QN());
   DFFS_X1 \buf_fill_i_reg[3]  (.D(\out_bs[7] [3]), .SN(n_0_169), .CK(n_0_171), 
      .Q(buf_fill_i[3]), .QN());
   DFFS_X1 \buf_fill_i_reg[2]  (.D(\out_bs[7] [2]), .SN(n_0_169), .CK(n_0_171), 
      .Q(buf_fill_i[2]), .QN());
   DFFS_X1 \buf_fill_i_reg[1]  (.D(\out_bs[7] [1]), .SN(n_0_169), .CK(n_0_171), 
      .Q(buf_fill_i[1]), .QN());
   DFFS_X1 \buf_fill_i_reg[0]  (.D(\out_bs[7] [0]), .SN(n_0_169), .CK(n_0_171), 
      .Q(buf_fill_i[0]), .QN());
   DFFS_X1 buf_is_empty_reg (.D(1'b0), .SN(n_0_169), .CK(n_0_171), .Q(
      buf_is_empty), .QN());
   CLKGATETST_X1 clk_gate_buf_fill_i_reg (.CK(clk), .E(enbl_in), .SE(1'b0), 
      .GCK(n_0_171));
   NOR3_X1 i_0_1_0 (.A1(buf_is_empty), .A2(rst), .A3(n_0_1_68), .ZN(n_0_40));
   NOR2_X1 i_0_1_1 (.A1(n_0_1_1), .A2(n_0_1_0), .ZN(n_0_7));
   OAI22_X1 i_0_1_2 (.A1(n_0_99), .A2(n_0_1_64), .B1(n_0_1_63), .B2(n_0_67), 
      .ZN(n_0_1_0));
   OAI22_X1 i_0_1_3 (.A1(n_0_1_66), .A2(n_0_131), .B1(n_0_1_69), .B2(n_0_0), 
      .ZN(n_0_1_1));
   NOR2_X1 i_0_1_4 (.A1(n_0_1_3), .A2(n_0_1_2), .ZN(n_0_8));
   OAI22_X1 i_0_1_5 (.A1(n_0_100), .A2(n_0_1_64), .B1(n_0_1_63), .B2(n_0_68), 
      .ZN(n_0_1_2));
   OAI22_X1 i_0_1_6 (.A1(n_0_1_66), .A2(n_0_132), .B1(n_0_1_69), .B2(n_0_1), 
      .ZN(n_0_1_3));
   NOR2_X1 i_0_1_7 (.A1(n_0_1_5), .A2(n_0_1_4), .ZN(n_0_9));
   OAI22_X1 i_0_1_8 (.A1(n_0_101), .A2(n_0_1_64), .B1(n_0_1_63), .B2(n_0_69), 
      .ZN(n_0_1_4));
   OAI22_X1 i_0_1_9 (.A1(n_0_1_66), .A2(n_0_133), .B1(n_0_1_69), .B2(n_0_2), 
      .ZN(n_0_1_5));
   NOR2_X1 i_0_1_10 (.A1(n_0_1_7), .A2(n_0_1_6), .ZN(n_0_10));
   OAI22_X1 i_0_1_11 (.A1(n_0_102), .A2(n_0_1_64), .B1(n_0_1_63), .B2(n_0_70), 
      .ZN(n_0_1_6));
   OAI22_X1 i_0_1_12 (.A1(n_0_1_66), .A2(n_0_134), .B1(n_0_1_69), .B2(n_0_3), 
      .ZN(n_0_1_7));
   NOR2_X1 i_0_1_13 (.A1(n_0_1_9), .A2(n_0_1_8), .ZN(n_0_11));
   OAI22_X1 i_0_1_14 (.A1(n_0_103), .A2(n_0_1_64), .B1(n_0_1_63), .B2(n_0_71), 
      .ZN(n_0_1_8));
   OAI22_X1 i_0_1_15 (.A1(n_0_1_66), .A2(n_0_135), .B1(n_0_1_69), .B2(n_0_4), 
      .ZN(n_0_1_9));
   NOR2_X1 i_0_1_16 (.A1(n_0_1_11), .A2(n_0_1_10), .ZN(n_0_12));
   OAI22_X1 i_0_1_17 (.A1(n_0_104), .A2(n_0_1_64), .B1(n_0_1_63), .B2(n_0_72), 
      .ZN(n_0_1_10));
   OAI22_X1 i_0_1_18 (.A1(n_0_1_66), .A2(n_0_136), .B1(n_0_1_69), .B2(n_0_6), 
      .ZN(n_0_1_11));
   NOR2_X1 i_0_1_19 (.A1(n_0_1_13), .A2(n_0_1_12), .ZN(n_0_13));
   OAI22_X1 i_0_1_20 (.A1(n_0_105), .A2(n_0_1_64), .B1(n_0_1_63), .B2(n_0_73), 
      .ZN(n_0_1_12));
   OAI22_X1 i_0_1_21 (.A1(n_0_1_66), .A2(n_0_137), .B1(n_0_1_69), .B2(n_0_41), 
      .ZN(n_0_1_13));
   NOR2_X1 i_0_1_22 (.A1(n_0_1_15), .A2(n_0_1_14), .ZN(n_0_14));
   OAI22_X1 i_0_1_23 (.A1(n_0_106), .A2(n_0_1_64), .B1(n_0_1_63), .B2(n_0_74), 
      .ZN(n_0_1_14));
   OAI22_X1 i_0_1_24 (.A1(n_0_1_66), .A2(n_0_138), .B1(n_0_1_69), .B2(n_0_42), 
      .ZN(n_0_1_15));
   NOR2_X1 i_0_1_25 (.A1(n_0_1_17), .A2(n_0_1_16), .ZN(n_0_15));
   OAI22_X1 i_0_1_26 (.A1(n_0_107), .A2(n_0_1_64), .B1(n_0_1_63), .B2(n_0_75), 
      .ZN(n_0_1_16));
   OAI22_X1 i_0_1_27 (.A1(n_0_1_66), .A2(n_0_139), .B1(n_0_1_69), .B2(n_0_43), 
      .ZN(n_0_1_17));
   NOR2_X1 i_0_1_28 (.A1(n_0_1_19), .A2(n_0_1_18), .ZN(n_0_16));
   OAI22_X1 i_0_1_29 (.A1(n_0_108), .A2(n_0_1_64), .B1(n_0_1_63), .B2(n_0_76), 
      .ZN(n_0_1_18));
   OAI22_X1 i_0_1_30 (.A1(n_0_1_66), .A2(n_0_140), .B1(n_0_1_69), .B2(n_0_44), 
      .ZN(n_0_1_19));
   NOR2_X1 i_0_1_31 (.A1(n_0_1_21), .A2(n_0_1_20), .ZN(n_0_17));
   OAI22_X1 i_0_1_32 (.A1(n_0_109), .A2(n_0_1_64), .B1(n_0_1_63), .B2(n_0_77), 
      .ZN(n_0_1_20));
   OAI22_X1 i_0_1_33 (.A1(n_0_1_66), .A2(n_0_141), .B1(n_0_1_69), .B2(n_0_45), 
      .ZN(n_0_1_21));
   NOR2_X1 i_0_1_34 (.A1(n_0_1_23), .A2(n_0_1_22), .ZN(n_0_18));
   OAI22_X1 i_0_1_35 (.A1(n_0_110), .A2(n_0_1_64), .B1(n_0_1_63), .B2(n_0_78), 
      .ZN(n_0_1_22));
   OAI22_X1 i_0_1_36 (.A1(n_0_1_66), .A2(n_0_142), .B1(n_0_1_69), .B2(n_0_46), 
      .ZN(n_0_1_23));
   NOR2_X1 i_0_1_37 (.A1(n_0_1_25), .A2(n_0_1_24), .ZN(n_0_19));
   OAI22_X1 i_0_1_38 (.A1(n_0_111), .A2(n_0_1_64), .B1(n_0_1_63), .B2(n_0_79), 
      .ZN(n_0_1_24));
   OAI22_X1 i_0_1_39 (.A1(n_0_1_66), .A2(n_0_143), .B1(n_0_1_69), .B2(n_0_47), 
      .ZN(n_0_1_25));
   NOR2_X1 i_0_1_40 (.A1(n_0_1_27), .A2(n_0_1_26), .ZN(n_0_20));
   OAI22_X1 i_0_1_41 (.A1(n_0_112), .A2(n_0_1_64), .B1(n_0_1_63), .B2(n_0_80), 
      .ZN(n_0_1_26));
   OAI22_X1 i_0_1_42 (.A1(n_0_1_66), .A2(n_0_144), .B1(n_0_1_69), .B2(n_0_48), 
      .ZN(n_0_1_27));
   NOR2_X1 i_0_1_43 (.A1(n_0_1_29), .A2(n_0_1_28), .ZN(n_0_21));
   OAI22_X1 i_0_1_44 (.A1(n_0_113), .A2(n_0_1_64), .B1(n_0_1_63), .B2(n_0_81), 
      .ZN(n_0_1_28));
   OAI22_X1 i_0_1_45 (.A1(n_0_1_66), .A2(n_0_145), .B1(n_0_1_69), .B2(n_0_49), 
      .ZN(n_0_1_29));
   NOR2_X1 i_0_1_46 (.A1(n_0_1_31), .A2(n_0_1_30), .ZN(n_0_22));
   OAI22_X1 i_0_1_47 (.A1(n_0_114), .A2(n_0_1_64), .B1(n_0_1_63), .B2(n_0_82), 
      .ZN(n_0_1_30));
   OAI22_X1 i_0_1_48 (.A1(n_0_1_66), .A2(n_0_146), .B1(n_0_1_69), .B2(n_0_50), 
      .ZN(n_0_1_31));
   NOR2_X1 i_0_1_49 (.A1(n_0_1_33), .A2(n_0_1_32), .ZN(n_0_23));
   OAI22_X1 i_0_1_50 (.A1(n_0_115), .A2(n_0_1_64), .B1(n_0_1_63), .B2(n_0_83), 
      .ZN(n_0_1_32));
   OAI22_X1 i_0_1_51 (.A1(n_0_1_66), .A2(n_0_147), .B1(n_0_1_69), .B2(n_0_51), 
      .ZN(n_0_1_33));
   NOR2_X1 i_0_1_52 (.A1(n_0_1_35), .A2(n_0_1_34), .ZN(n_0_24));
   OAI22_X1 i_0_1_53 (.A1(n_0_116), .A2(n_0_1_64), .B1(n_0_1_63), .B2(n_0_84), 
      .ZN(n_0_1_34));
   OAI22_X1 i_0_1_54 (.A1(n_0_1_66), .A2(n_0_148), .B1(n_0_1_69), .B2(n_0_52), 
      .ZN(n_0_1_35));
   NOR2_X1 i_0_1_55 (.A1(n_0_1_37), .A2(n_0_1_36), .ZN(n_0_25));
   OAI22_X1 i_0_1_56 (.A1(n_0_117), .A2(n_0_1_64), .B1(n_0_1_63), .B2(n_0_85), 
      .ZN(n_0_1_36));
   OAI22_X1 i_0_1_57 (.A1(n_0_1_66), .A2(n_0_149), .B1(n_0_1_69), .B2(n_0_53), 
      .ZN(n_0_1_37));
   NOR2_X1 i_0_1_58 (.A1(n_0_1_39), .A2(n_0_1_38), .ZN(n_0_26));
   OAI22_X1 i_0_1_59 (.A1(n_0_118), .A2(n_0_1_64), .B1(n_0_1_63), .B2(n_0_86), 
      .ZN(n_0_1_38));
   OAI22_X1 i_0_1_60 (.A1(n_0_1_66), .A2(n_0_150), .B1(n_0_1_69), .B2(n_0_54), 
      .ZN(n_0_1_39));
   NOR2_X1 i_0_1_61 (.A1(n_0_1_41), .A2(n_0_1_40), .ZN(n_0_27));
   OAI22_X1 i_0_1_62 (.A1(n_0_119), .A2(n_0_1_64), .B1(n_0_1_63), .B2(n_0_87), 
      .ZN(n_0_1_40));
   OAI22_X1 i_0_1_63 (.A1(n_0_1_66), .A2(n_0_151), .B1(n_0_1_69), .B2(n_0_55), 
      .ZN(n_0_1_41));
   NOR2_X1 i_0_1_64 (.A1(n_0_1_43), .A2(n_0_1_42), .ZN(n_0_28));
   OAI22_X1 i_0_1_65 (.A1(n_0_120), .A2(n_0_1_64), .B1(n_0_1_63), .B2(n_0_88), 
      .ZN(n_0_1_42));
   OAI22_X1 i_0_1_66 (.A1(n_0_1_66), .A2(n_0_152), .B1(n_0_1_69), .B2(n_0_56), 
      .ZN(n_0_1_43));
   NOR2_X1 i_0_1_67 (.A1(n_0_1_45), .A2(n_0_1_44), .ZN(n_0_29));
   OAI22_X1 i_0_1_68 (.A1(n_0_121), .A2(n_0_1_64), .B1(n_0_1_63), .B2(n_0_89), 
      .ZN(n_0_1_44));
   OAI22_X1 i_0_1_69 (.A1(n_0_1_66), .A2(n_0_153), .B1(n_0_1_69), .B2(n_0_57), 
      .ZN(n_0_1_45));
   NOR2_X1 i_0_1_70 (.A1(n_0_1_47), .A2(n_0_1_46), .ZN(n_0_30));
   OAI22_X1 i_0_1_71 (.A1(n_0_122), .A2(n_0_1_64), .B1(n_0_1_63), .B2(n_0_90), 
      .ZN(n_0_1_46));
   OAI22_X1 i_0_1_72 (.A1(n_0_1_66), .A2(n_0_154), .B1(n_0_1_69), .B2(n_0_58), 
      .ZN(n_0_1_47));
   NOR2_X1 i_0_1_73 (.A1(n_0_1_49), .A2(n_0_1_48), .ZN(n_0_31));
   OAI22_X1 i_0_1_74 (.A1(n_0_123), .A2(n_0_1_64), .B1(n_0_1_63), .B2(n_0_91), 
      .ZN(n_0_1_48));
   OAI22_X1 i_0_1_75 (.A1(n_0_1_66), .A2(n_0_155), .B1(n_0_1_69), .B2(n_0_59), 
      .ZN(n_0_1_49));
   NOR2_X1 i_0_1_76 (.A1(n_0_1_51), .A2(n_0_1_50), .ZN(n_0_32));
   OAI22_X1 i_0_1_77 (.A1(n_0_124), .A2(n_0_1_64), .B1(n_0_1_63), .B2(n_0_92), 
      .ZN(n_0_1_50));
   OAI22_X1 i_0_1_78 (.A1(n_0_1_66), .A2(n_0_156), .B1(n_0_1_69), .B2(n_0_60), 
      .ZN(n_0_1_51));
   NOR2_X1 i_0_1_79 (.A1(n_0_1_53), .A2(n_0_1_52), .ZN(n_0_33));
   OAI22_X1 i_0_1_80 (.A1(n_0_125), .A2(n_0_1_64), .B1(n_0_1_63), .B2(n_0_93), 
      .ZN(n_0_1_52));
   OAI22_X1 i_0_1_81 (.A1(n_0_1_66), .A2(n_0_157), .B1(n_0_1_69), .B2(n_0_61), 
      .ZN(n_0_1_53));
   NOR2_X1 i_0_1_82 (.A1(n_0_1_55), .A2(n_0_1_54), .ZN(n_0_34));
   OAI22_X1 i_0_1_83 (.A1(n_0_126), .A2(n_0_1_64), .B1(n_0_1_63), .B2(n_0_94), 
      .ZN(n_0_1_54));
   OAI22_X1 i_0_1_84 (.A1(n_0_1_66), .A2(n_0_158), .B1(n_0_1_69), .B2(n_0_62), 
      .ZN(n_0_1_55));
   NOR2_X1 i_0_1_85 (.A1(n_0_1_57), .A2(n_0_1_56), .ZN(n_0_35));
   OAI22_X1 i_0_1_86 (.A1(n_0_127), .A2(n_0_1_64), .B1(n_0_1_63), .B2(n_0_95), 
      .ZN(n_0_1_56));
   OAI22_X1 i_0_1_87 (.A1(n_0_1_66), .A2(n_0_159), .B1(n_0_1_69), .B2(n_0_63), 
      .ZN(n_0_1_57));
   NOR2_X1 i_0_1_88 (.A1(n_0_1_59), .A2(n_0_1_58), .ZN(n_0_36));
   OAI22_X1 i_0_1_89 (.A1(n_0_128), .A2(n_0_1_64), .B1(n_0_1_63), .B2(n_0_96), 
      .ZN(n_0_1_58));
   OAI22_X1 i_0_1_90 (.A1(n_0_1_66), .A2(n_0_160), .B1(n_0_1_69), .B2(n_0_64), 
      .ZN(n_0_1_59));
   NOR2_X1 i_0_1_91 (.A1(n_0_1_61), .A2(n_0_1_60), .ZN(n_0_37));
   OAI22_X1 i_0_1_92 (.A1(n_0_129), .A2(n_0_1_64), .B1(n_0_1_63), .B2(n_0_97), 
      .ZN(n_0_1_60));
   OAI22_X1 i_0_1_93 (.A1(n_0_1_66), .A2(n_0_161), .B1(n_0_1_69), .B2(n_0_65), 
      .ZN(n_0_1_61));
   NOR2_X1 i_0_1_94 (.A1(n_0_1_65), .A2(n_0_1_62), .ZN(n_0_38));
   OAI22_X1 i_0_1_95 (.A1(n_0_130), .A2(n_0_1_64), .B1(n_0_1_63), .B2(n_0_98), 
      .ZN(n_0_1_62));
   NAND2_X1 i_0_1_96 (.A1(n_0_1_78), .A2(buf_flush_i[6]), .ZN(n_0_1_63));
   NAND2_X1 i_0_1_97 (.A1(n_0_1_79), .A2(buf_flush_i[5]), .ZN(n_0_1_64));
   OAI22_X1 i_0_1_98 (.A1(n_0_1_66), .A2(n_0_162), .B1(n_0_1_69), .B2(n_0_66), 
      .ZN(n_0_1_65));
   NAND2_X1 i_0_1_99 (.A1(n_0_1_79), .A2(n_0_1_78), .ZN(n_0_1_66));
   NOR2_X1 i_0_1_100 (.A1(n_0_5), .A2(n_0_1_67), .ZN(n_0_163));
   OAI21_X1 i_0_1_101 (.A(state_wait), .B1(n_0_1_74), .B2(n_0_1_70), .ZN(
      n_0_1_67));
   NOR2_X1 i_0_1_102 (.A1(buf_is_empty), .A2(n_0_1_68), .ZN(n_0_5));
   AOI22_X1 i_0_1_103 (.A1(n_0_1_74), .A2(n_0_1_71), .B1(n_0_1_70), .B2(n_0_1_76), 
      .ZN(n_0_1_68));
   NAND2_X1 i_0_1_104 (.A1(buf_flush_i[6]), .A2(buf_flush_i[5]), .ZN(n_0_1_69));
   OAI22_X1 i_0_1_105 (.A1(n_0_1_79), .A2(\out_as[0] [6]), .B1(n_0_1_78), 
      .B2(\out_as[0] [5]), .ZN(n_0_1_70));
   INV_X1 i_0_1_106 (.A(n_0_1_72), .ZN(n_0_1_71));
   AOI211_X1 i_0_1_107 (.A(buf_fill_flush_diff[6]), .B(buf_fill_flush_diff[5]), 
      .C1(\out_as[0] [1]), .C2(n_0_1_73), .ZN(n_0_1_72));
   AND4_X1 i_0_1_108 (.A1(\out_as[0] [4]), .A2(\out_as[0] [3]), .A3(
      \out_as[0] [2]), .A4(\out_as[0] [0]), .ZN(n_0_1_73));
   NAND3_X1 i_0_1_109 (.A1(n_0_1_77), .A2(n_0_1_75), .A3(n_0_1_76), .ZN(n_0_1_74));
   AOI211_X1 i_0_1_110 (.A(\out_as[0] [4]), .B(\out_as[0] [3]), .C1(n_0_1_78), 
      .C2(\out_as[0] [5]), .ZN(n_0_1_75));
   NAND2_X1 i_0_1_111 (.A1(n_0_1_79), .A2(\out_as[0] [6]), .ZN(n_0_1_76));
   NOR3_X1 i_0_1_112 (.A1(\out_as[0] [2]), .A2(\out_as[0] [1]), .A3(
      \out_as[0] [0]), .ZN(n_0_1_77));
   INV_X1 i_0_1_113 (.A(rst), .ZN(n_0_169));
   INV_X1 i_0_1_114 (.A(buf_flush_i[5]), .ZN(n_0_1_78));
   INV_X1 i_0_1_115 (.A(buf_flush_i[6]), .ZN(n_0_1_79));
   INV_X1 error_success_reg_enable_mux_0 (.A(error_success), .ZN(
      error_success_reg_enable_mux_n_0));
   NOR2_X1 error_success_reg_enable_mux_1 (.A1(error_success_reg_enable_mux_n_0), 
      .A2(n_0_163), .ZN(n_0_164));
   MUX2_X1 i_0_0_0 (.A(n_0_0), .B(n_110), .S(n_186), .Z(n_0_295));
   MUX2_X1 i_0_0_1 (.A(n_0_1), .B(n_109), .S(n_255), .Z(n_0_294));
   MUX2_X1 i_0_0_2 (.A(n_0_2), .B(n_108), .S(n_185), .Z(n_0_293));
   MUX2_X1 i_0_0_3 (.A(n_0_3), .B(n_107), .S(n_184), .Z(n_0_292));
   MUX2_X1 i_0_0_4 (.A(n_0_4), .B(n_106), .S(n_183), .Z(n_0_291));
   MUX2_X1 i_0_0_5 (.A(n_0_6), .B(n_105), .S(n_254), .Z(n_0_290));
   MUX2_X1 i_0_0_6 (.A(n_0_41), .B(n_104), .S(n_182), .Z(n_0_289));
   MUX2_X1 i_0_0_7 (.A(n_0_42), .B(n_103), .S(n_181), .Z(n_0_288));
   MUX2_X1 i_0_0_8 (.A(n_0_43), .B(n_102), .S(n_253), .Z(n_0_287));
   MUX2_X1 i_0_0_9 (.A(n_0_44), .B(n_101), .S(n_180), .Z(n_0_286));
   MUX2_X1 i_0_0_10 (.A(n_0_45), .B(n_100), .S(n_252), .Z(n_0_285));
   MUX2_X1 i_0_0_11 (.A(n_0_46), .B(n_99), .S(n_179), .Z(n_0_284));
   MUX2_X1 i_0_0_12 (.A(n_0_47), .B(n_98), .S(n_251), .Z(n_0_283));
   MUX2_X1 i_0_0_13 (.A(n_0_48), .B(n_97), .S(n_178), .Z(n_0_282));
   MUX2_X1 i_0_0_14 (.A(n_0_49), .B(n_96), .S(n_177), .Z(n_0_281));
   MUX2_X1 i_0_0_15 (.A(n_0_50), .B(n_95), .S(n_176), .Z(n_0_280));
   MUX2_X1 i_0_0_16 (.A(n_0_51), .B(n_215), .S(n_250), .Z(n_0_279));
   MUX2_X1 i_0_0_17 (.A(n_0_52), .B(n_94), .S(n_175), .Z(n_0_278));
   MUX2_X1 i_0_0_18 (.A(n_0_53), .B(n_93), .S(n_174), .Z(n_0_277));
   MUX2_X1 i_0_0_19 (.A(n_0_54), .B(n_92), .S(n_173), .Z(n_0_276));
   MUX2_X1 i_0_0_20 (.A(n_0_55), .B(n_91), .S(n_172), .Z(n_0_275));
   MUX2_X1 i_0_0_21 (.A(n_0_56), .B(n_90), .S(n_171), .Z(n_0_274));
   MUX2_X1 i_0_0_22 (.A(n_0_57), .B(n_89), .S(n_170), .Z(n_0_273));
   MUX2_X1 i_0_0_23 (.A(n_0_58), .B(n_88), .S(n_169), .Z(n_0_272));
   MUX2_X1 i_0_0_24 (.A(n_0_59), .B(n_87), .S(n_168), .Z(n_0_271));
   MUX2_X1 i_0_0_25 (.A(n_0_60), .B(n_86), .S(n_167), .Z(n_0_270));
   MUX2_X1 i_0_0_26 (.A(n_0_61), .B(n_85), .S(n_166), .Z(n_0_269));
   MUX2_X1 i_0_0_27 (.A(n_0_62), .B(n_84), .S(n_165), .Z(n_0_268));
   MUX2_X1 i_0_0_28 (.A(n_0_63), .B(n_83), .S(n_164), .Z(n_0_267));
   MUX2_X1 i_0_0_29 (.A(n_0_64), .B(n_82), .S(n_163), .Z(n_0_266));
   MUX2_X1 i_0_0_30 (.A(n_0_65), .B(n_81), .S(n_162), .Z(n_0_265));
   MUX2_X1 i_0_0_31 (.A(n_0_66), .B(n_80), .S(n_161), .Z(n_0_264));
   MUX2_X1 i_0_0_32 (.A(n_0_67), .B(n_79), .S(n_160), .Z(n_0_263));
   MUX2_X1 i_0_0_33 (.A(n_0_68), .B(n_78), .S(n_249), .Z(n_0_262));
   MUX2_X1 i_0_0_34 (.A(n_0_69), .B(n_77), .S(n_248), .Z(n_0_261));
   MUX2_X1 i_0_0_35 (.A(n_0_70), .B(n_76), .S(n_247), .Z(n_0_260));
   MUX2_X1 i_0_0_36 (.A(n_0_71), .B(n_75), .S(n_159), .Z(n_0_259));
   MUX2_X1 i_0_0_37 (.A(n_0_72), .B(n_74), .S(n_158), .Z(n_0_258));
   MUX2_X1 i_0_0_38 (.A(n_0_73), .B(n_73), .S(n_157), .Z(n_0_257));
   MUX2_X1 i_0_0_39 (.A(n_0_74), .B(n_72), .S(n_156), .Z(n_0_256));
   MUX2_X1 i_0_0_40 (.A(n_0_75), .B(n_71), .S(n_155), .Z(n_0_255));
   MUX2_X1 i_0_0_41 (.A(n_0_76), .B(n_70), .S(n_154), .Z(n_0_254));
   MUX2_X1 i_0_0_42 (.A(n_0_77), .B(n_69), .S(n_246), .Z(n_0_253));
   MUX2_X1 i_0_0_43 (.A(n_0_78), .B(n_68), .S(n_153), .Z(n_0_252));
   MUX2_X1 i_0_0_44 (.A(n_0_79), .B(n_67), .S(n_152), .Z(n_0_251));
   MUX2_X1 i_0_0_45 (.A(n_0_80), .B(n_66), .S(n_151), .Z(n_0_250));
   MUX2_X1 i_0_0_46 (.A(n_0_81), .B(n_65), .S(n_245), .Z(n_0_249));
   MUX2_X1 i_0_0_47 (.A(n_0_82), .B(n_64), .S(n_150), .Z(n_0_248));
   MUX2_X1 i_0_0_48 (.A(n_0_83), .B(n_63), .S(n_149), .Z(n_0_247));
   MUX2_X1 i_0_0_49 (.A(n_0_84), .B(n_62), .S(n_148), .Z(n_0_246));
   MUX2_X1 i_0_0_50 (.A(n_0_85), .B(n_61), .S(n_147), .Z(n_0_245));
   MUX2_X1 i_0_0_51 (.A(n_0_86), .B(n_60), .S(n_146), .Z(n_0_244));
   MUX2_X1 i_0_0_52 (.A(n_0_87), .B(n_59), .S(n_145), .Z(n_0_243));
   MUX2_X1 i_0_0_53 (.A(n_0_88), .B(n_58), .S(n_144), .Z(n_0_242));
   MUX2_X1 i_0_0_54 (.A(n_0_89), .B(n_57), .S(n_244), .Z(n_0_241));
   MUX2_X1 i_0_0_55 (.A(n_0_90), .B(n_56), .S(n_243), .Z(n_0_240));
   MUX2_X1 i_0_0_56 (.A(n_0_91), .B(n_55), .S(n_143), .Z(n_0_239));
   MUX2_X1 i_0_0_57 (.A(n_0_92), .B(n_54), .S(n_142), .Z(n_0_238));
   MUX2_X1 i_0_0_58 (.A(n_0_93), .B(n_53), .S(n_141), .Z(n_0_237));
   MUX2_X1 i_0_0_59 (.A(n_0_94), .B(n_52), .S(n_140), .Z(n_0_236));
   MUX2_X1 i_0_0_60 (.A(n_0_95), .B(n_51), .S(n_139), .Z(n_0_235));
   MUX2_X1 i_0_0_61 (.A(n_0_96), .B(n_50), .S(n_138), .Z(n_0_234));
   MUX2_X1 i_0_0_62 (.A(n_0_97), .B(n_49), .S(n_137), .Z(n_0_233));
   MUX2_X1 i_0_0_63 (.A(n_0_98), .B(n_48), .S(n_242), .Z(n_0_232));
   MUX2_X1 i_0_0_64 (.A(n_0_99), .B(n_47), .S(n_199), .Z(n_0_231));
   MUX2_X1 i_0_0_65 (.A(n_0_100), .B(n_46), .S(n_136), .Z(n_0_230));
   MUX2_X1 i_0_0_66 (.A(n_0_101), .B(n_45), .S(n_198), .Z(n_0_229));
   MUX2_X1 i_0_0_67 (.A(n_0_102), .B(n_44), .S(n_241), .Z(n_0_228));
   MUX2_X1 i_0_0_68 (.A(n_0_103), .B(n_43), .S(n_135), .Z(n_0_227));
   MUX2_X1 i_0_0_69 (.A(n_0_104), .B(n_214), .S(n_240), .Z(n_0_226));
   MUX2_X1 i_0_0_70 (.A(n_0_105), .B(n_42), .S(n_239), .Z(n_0_225));
   MUX2_X1 i_0_0_71 (.A(n_0_106), .B(n_41), .S(n_134), .Z(n_0_224));
   MUX2_X1 i_0_0_73 (.A(n_0_108), .B(n_40), .S(n_197), .Z(n_0_222));
   MUX2_X1 i_0_0_74 (.A(n_0_109), .B(n_39), .S(n_196), .Z(n_0_221));
   MUX2_X1 i_0_0_75 (.A(n_0_110), .B(n_38), .S(n_133), .Z(n_0_220));
   MUX2_X1 i_0_0_76 (.A(n_0_111), .B(n_213), .S(n_238), .Z(n_0_219));
   MUX2_X1 i_0_0_77 (.A(n_0_112), .B(n_37), .S(n_201), .Z(n_0_218));
   MUX2_X1 i_0_0_78 (.A(n_0_113), .B(n_212), .S(n_237), .Z(n_0_217));
   MUX2_X1 i_0_0_79 (.A(n_0_114), .B(n_211), .S(n_132), .Z(n_0_216));
   MUX2_X1 i_0_0_80 (.A(n_0_115), .B(n_36), .S(n_236), .Z(n_0_215));
   MUX2_X1 i_0_0_81 (.A(n_0_116), .B(n_35), .S(n_195), .Z(n_0_214));
   MUX2_X1 i_0_0_82 (.A(n_0_117), .B(n_34), .S(n_194), .Z(n_0_213));
   MUX2_X1 i_0_0_83 (.A(n_0_118), .B(n_33), .S(n_235), .Z(n_0_212));
   MUX2_X1 i_0_0_84 (.A(n_0_119), .B(n_32), .S(n_131), .Z(n_0_211));
   MUX2_X1 i_0_0_85 (.A(n_0_120), .B(n_31), .S(n_130), .Z(n_0_210));
   MUX2_X1 i_0_0_86 (.A(n_0_121), .B(n_30), .S(n_193), .Z(n_0_209));
   MUX2_X1 i_0_0_87 (.A(n_0_122), .B(n_29), .S(n_234), .Z(n_0_208));
   MUX2_X1 i_0_0_88 (.A(n_0_123), .B(n_28), .S(n_192), .Z(n_0_207));
   MUX2_X1 i_0_0_89 (.A(n_0_124), .B(n_210), .S(n_233), .Z(n_0_206));
   MUX2_X1 i_0_0_90 (.A(n_0_125), .B(n_209), .S(n_232), .Z(n_0_205));
   MUX2_X1 i_0_0_91 (.A(n_0_126), .B(n_27), .S(n_129), .Z(n_0_204));
   MUX2_X1 i_0_0_92 (.A(n_0_127), .B(n_188), .S(n_191), .Z(n_0_203));
   MUX2_X1 i_0_0_93 (.A(n_0_128), .B(n_26), .S(n_128), .Z(n_0_202));
   MUX2_X1 i_0_0_94 (.A(n_0_129), .B(n_200), .S(n_231), .Z(n_0_201));
   MUX2_X1 i_0_0_95 (.A(n_0_130), .B(n_25), .S(n_230), .Z(n_0_200));
   MUX2_X1 i_0_0_96 (.A(n_0_131), .B(n_24), .S(n_127), .Z(n_0_199));
   MUX2_X1 i_0_0_97 (.A(n_0_132), .B(n_23), .S(n_229), .Z(n_0_198));
   MUX2_X1 i_0_0_98 (.A(n_0_133), .B(n_22), .S(n_228), .Z(n_0_197));
   MUX2_X1 i_0_0_99 (.A(n_0_134), .B(n_21), .S(n_227), .Z(n_0_196));
   MUX2_X1 i_0_0_100 (.A(n_0_135), .B(n_20), .S(n_126), .Z(n_0_195));
   MUX2_X1 i_0_0_101 (.A(n_0_136), .B(n_19), .S(n_125), .Z(n_0_194));
   MUX2_X1 i_0_0_102 (.A(n_0_137), .B(n_208), .S(n_226), .Z(n_0_193));
   MUX2_X1 i_0_0_103 (.A(n_0_138), .B(n_18), .S(n_124), .Z(n_0_192));
   MUX2_X1 i_0_0_104 (.A(n_0_139), .B(n_17), .S(n_123), .Z(n_0_191));
   MUX2_X1 i_0_0_105 (.A(n_0_140), .B(n_16), .S(n_122), .Z(n_0_190));
   MUX2_X1 i_0_0_106 (.A(n_0_141), .B(n_207), .S(n_225), .Z(n_0_189));
   MUX2_X1 i_0_0_107 (.A(n_0_142), .B(n_206), .S(n_224), .Z(n_0_188));
   MUX2_X1 i_0_0_108 (.A(n_0_143), .B(n_205), .S(n_121), .Z(n_0_187));
   MUX2_X1 i_0_0_109 (.A(n_0_144), .B(n_204), .S(n_223), .Z(n_0_186));
   MUX2_X1 i_0_0_110 (.A(n_0_145), .B(n_15), .S(n_120), .Z(n_0_185));
   MUX2_X1 i_0_0_111 (.A(n_0_146), .B(n_14), .S(n_222), .Z(n_0_184));
   MUX2_X1 i_0_0_112 (.A(n_0_147), .B(n_13), .S(n_221), .Z(n_0_183));
   MUX2_X1 i_0_0_113 (.A(n_0_148), .B(n_12), .S(n_119), .Z(n_0_182));
   MUX2_X1 i_0_0_114 (.A(n_0_149), .B(n_11), .S(n_220), .Z(n_0_181));
   MUX2_X1 i_0_0_115 (.A(n_0_150), .B(n_10), .S(n_219), .Z(n_0_180));
   MUX2_X1 i_0_0_116 (.A(n_0_151), .B(n_203), .S(n_218), .Z(n_0_179));
   MUX2_X1 i_0_0_117 (.A(n_0_152), .B(n_9), .S(n_118), .Z(n_0_178));
   MUX2_X1 i_0_0_118 (.A(n_0_153), .B(n_8), .S(n_117), .Z(n_0_177));
   MUX2_X1 i_0_0_119 (.A(n_0_154), .B(n_7), .S(n_190), .Z(n_0_176));
   MUX2_X1 i_0_0_120 (.A(n_0_155), .B(n_202), .S(n_116), .Z(n_0_175));
   MUX2_X1 i_0_0_121 (.A(n_0_156), .B(n_6), .S(n_217), .Z(n_0_174));
   MUX2_X1 i_0_0_122 (.A(n_0_157), .B(n_5), .S(n_115), .Z(n_0_173));
   MUX2_X1 i_0_0_123 (.A(n_0_158), .B(n_4), .S(n_114), .Z(n_0_172));
   MUX2_X1 i_0_0_124 (.A(n_0_159), .B(n_3), .S(n_113), .Z(n_0_168));
   MUX2_X1 i_0_0_125 (.A(n_0_160), .B(n_2), .S(n_112), .Z(n_0_167));
   MUX2_X1 i_0_0_126 (.A(n_0_161), .B(n_1), .S(n_216), .Z(n_0_166));
   MUX2_X1 i_0_0_127 (.A(n_0_162), .B(n_0), .S(n_111), .Z(n_0_165));
   OAI21_X1 i_0_0_72 (.A(n_0_0_0), .B1(n_0_0_1), .B2(n_187), .ZN(n_0_223));
   NAND2_X1 i_0_0_128 (.A1(n_187), .A2(n_189), .ZN(n_0_0_0));
   INV_X1 i_0_0_129 (.A(n_0_107), .ZN(n_0_0_1));
   range_extractor__3_149 range_extr_0 (.in_a(buf_fill_i), .in_size({in_data[31], 
      in_data[30], in_data[29]}), .out_a(\out_as[0] ), .out_b(\out_bs[0] ));
   int_adder__parameterized0 buf_flush_i_adder (.a({buf_flush_i[6], 
      buf_flush_i[5], uc_0, uc_1, uc_2, uc_3, uc_4}), .b(), .cin(), .enbl(), 
      .c({buf_flush_i_inc[6], buf_flush_i_inc[5], uc_5, uc_6, uc_7, uc_8, uc_9}), 
      .cout());
   int_adder__parameterized1 fill_flush_diff_subtractor (.a({\out_as[0] [6], 
      \out_as[0] [5], uc_10, uc_11, uc_12, uc_13, uc_14}), .b({
      buf_flush_i_inv[6], buf_flush_i_inc[5], uc_15, uc_16, uc_17, uc_18, uc_19}), 
      .cin(), .enbl(), .c({buf_fill_flush_diff[6], buf_fill_flush_diff[5], uc_20, 
      uc_21, uc_22, uc_23, uc_24}), .cout());
   range_extractor__3_201 ranges_1_range_extr_i (.in_a(\out_bs[0] ), .in_size({
      in_data[27], in_data[26], in_data[25]}), .out_a(\out_as[1] ), .out_b(
      \out_bs[1] ));
   range_extractor__3_253 ranges_2_range_extr_i (.in_a(\out_bs[1] ), .in_size({
      in_data[23], in_data[22], in_data[21]}), .out_a(\out_as[2] ), .out_b(
      \out_bs[2] ));
   range_extractor__3_305 ranges_3_range_extr_i (.in_a(\out_bs[2] ), .in_size({
      in_data[19], in_data[18], in_data[17]}), .out_a(\out_as[3] ), .out_b(
      \out_bs[3] ));
   range_extractor__3_357 ranges_4_range_extr_i (.in_a(\out_bs[3] ), .in_size({
      in_data[15], in_data[14], in_data[13]}), .out_a(\out_as[4] ), .out_b(
      \out_bs[4] ));
   range_extractor__3_409 ranges_5_range_extr_i (.in_a(\out_bs[4] ), .in_size({
      in_data[11], in_data[10], in_data[9]}), .out_a(\out_as[5] ), .out_b(
      \out_bs[5] ));
   range_extractor__3_461 ranges_6_range_extr_i (.in_a(\out_bs[5] ), .in_size({
      in_data[7], in_data[6], in_data[5]}), .out_a(\out_as[6] ), .out_b(
      \out_bs[6] ));
   range_extractor ranges_7_range_extr_i (.in_a(\out_bs[6] ), .in_size({
      in_data[3], in_data[2], in_data[1]}), .out_a(\out_as[7] ), .out_b(
      \out_bs[7] ));
   INV_X1 i_1_10_6 (.A(buf_flush_i[6]), .ZN(buf_flush_i_inv[6]));
endmodule

module full_adder__4_196(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(f));
   AND2_X1 i_0_1 (.A1(b), .A2(a), .ZN(cout));
endmodule

module full_adder__4_200(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   wire n_0_1;
   wire n_0_0;

   XOR2_X1 i_0_0 (.A(a), .B(b), .Z(n_0_1));
   XOR2_X1 i_0_1 (.A(n_0_1), .B(cin), .Z(f));
   AOI22_X1 i_0_2 (.A1(n_0_1), .A2(cin), .B1(a), .B2(b), .ZN(n_0_0));
   INV_X1 i_0_3 (.A(n_0_0), .ZN(cout));
endmodule

module full_adder__4_204(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__4_208(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__4_212(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__4_216(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__4_220(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__4_224(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__4_228(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__4_232(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__4_236(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__4_240(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__4_244(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__4_248(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__4_252(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(a), .ZN(cout));
endmodule

module full_adder__4_0(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(a), .B(cin), .Z(f));
endmodule

module int_adder__parameterized2(a, b, cin, enbl, c, cout);
   input [15:0]a;
   input [1:0]b;
   input cin;
   input enbl;
   output [15:0]c;
   output cout;

   full_adder__4_196 full_adder_0_0_full_adder_0_i (.a(a[0]), .b(b[0]), .cin(), 
      .f(c[0]), .cout(n_0));
   full_adder__4_200 full_adder_0_1_full_adder_0_i (.a(a[1]), .b(b[1]), .cin(n_0), 
      .f(c[1]), .cout(n_1));
   full_adder__4_204 full_adder_0_2_full_adder_0_i (.a(a[2]), .b(), .cin(n_1), 
      .f(c[2]), .cout(n_2));
   full_adder__4_208 full_adder_0_3_full_adder_0_i (.a(a[3]), .b(), .cin(n_2), 
      .f(c[3]), .cout(n_3));
   full_adder__4_212 full_adder_0_4_full_adder_0_i (.a(a[4]), .b(), .cin(n_3), 
      .f(c[4]), .cout(n_4));
   full_adder__4_216 full_adder_0_5_full_adder_0_i (.a(a[5]), .b(), .cin(n_4), 
      .f(c[5]), .cout(n_5));
   full_adder__4_220 full_adder_0_6_full_adder_0_i (.a(a[6]), .b(), .cin(n_5), 
      .f(c[6]), .cout(n_6));
   full_adder__4_224 full_adder_0_7_full_adder_0_i (.a(a[7]), .b(), .cin(n_6), 
      .f(c[7]), .cout(n_7));
   full_adder__4_228 full_adder_0_8_full_adder_0_i (.a(a[8]), .b(), .cin(n_7), 
      .f(c[8]), .cout(n_8));
   full_adder__4_232 full_adder_0_9_full_adder_0_i (.a(a[9]), .b(), .cin(n_8), 
      .f(c[9]), .cout(n_9));
   full_adder__4_236 full_adder_0_10_full_adder_0_i (.a(a[10]), .b(), .cin(n_9), 
      .f(c[10]), .cout(n_10));
   full_adder__4_240 full_adder_0_11_full_adder_0_i (.a(a[11]), .b(), .cin(n_10), 
      .f(c[11]), .cout(n_11));
   full_adder__4_244 full_adder_0_12_full_adder_0_i (.a(a[12]), .b(), .cin(n_11), 
      .f(c[12]), .cout(n_12));
   full_adder__4_248 full_adder_0_13_full_adder_0_i (.a(a[13]), .b(), .cin(n_12), 
      .f(c[13]), .cout(n_13));
   full_adder__4_252 full_adder_0_14_full_adder_0_i (.a(a[14]), .b(), .cin(n_13), 
      .f(c[14]), .cout(n_14));
   full_adder__4_0 full_adder_0_15_full_adder_0_i (.a(a[15]), .b(), .cin(n_14), 
      .f(c[15]), .cout());
endmodule

module datapath__0_5921(b, a, i);
   input [2:0]b;
   input [15:0]a;
   output [15:0]i;

   FA_X1 i_147 (.A(n_11), .B(n_10), .CI(n_27), .CO(n_39), .S(i[3]));
   FA_X1 i_148 (.A(n_9), .B(n_8), .CI(n_39), .CO(n_40), .S(i[4]));
   FA_X1 i_149 (.A(n_7), .B(n_6), .CI(n_40), .CO(n_0), .S(i[5]));
   FA_X1 i_150 (.A(n_5), .B(n_2), .CI(n_0), .CO(n_1), .S(i[6]));
   FA_X1 i_151 (.A(n_3), .B(n_4), .CI(n_1), .CO(i[8]), .S(i[7]));
   NOR2_X1 i_0 (.A1(n_12), .A2(n_3), .ZN(n_2));
   AND2_X1 i_1 (.A1(n_22), .A2(n_4), .ZN(n_3));
   AND2_X1 i_2 (.A1(b[2]), .A2(a[5]), .ZN(n_4));
   AOI22_X1 i_3 (.A1(b[1]), .A2(a[5]), .B1(b[2]), .B2(a[4]), .ZN(n_12));
   OAI21_X1 i_4 (.A(n_14), .B1(n_17), .B2(n_16), .ZN(n_5));
   XOR2_X1 i_5 (.A(n_17), .B(n_13), .Z(n_6));
   NAND2_X1 i_6 (.A1(n_15), .A2(n_14), .ZN(n_13));
   NAND3_X1 i_7 (.A1(b[0]), .A2(a[5]), .A3(n_22), .ZN(n_14));
   INV_X1 i_8 (.A(n_16), .ZN(n_15));
   AOI21_X1 i_9 (.A(n_22), .B1(b[0]), .B2(a[5]), .ZN(n_16));
   NAND2_X1 i_10 (.A1(b[2]), .A2(a[3]), .ZN(n_17));
   OAI21_X1 i_11 (.A(n_21), .B1(n_23), .B2(n_20), .ZN(n_7));
   XOR2_X1 i_12 (.A(n_23), .B(n_18), .Z(n_8));
   NAND2_X1 i_13 (.A1(n_21), .A2(n_19), .ZN(n_18));
   INV_X1 i_14 (.A(n_20), .ZN(n_19));
   AOI22_X1 i_15 (.A1(b[1]), .A2(a[3]), .B1(b[0]), .B2(a[4]), .ZN(n_20));
   NAND3_X1 i_16 (.A1(b[0]), .A2(a[3]), .A3(n_22), .ZN(n_21));
   AND2_X1 i_17 (.A1(b[1]), .A2(a[4]), .ZN(n_22));
   NAND2_X1 i_18 (.A1(b[2]), .A2(a[2]), .ZN(n_23));
   OAI21_X1 i_19 (.A(n_28), .B1(n_35), .B2(n_29), .ZN(n_9));
   INV_X1 i_20 (.A(n_24), .ZN(n_27));
   AOI22_X1 i_21 (.A1(n_36), .A2(n_32), .B1(n_37), .B2(n_31), .ZN(n_24));
   XOR2_X1 i_22 (.A(n_34), .B(n_25), .Z(n_10));
   NOR2_X1 i_23 (.A1(n_29), .A2(n_26), .ZN(n_25));
   INV_X1 i_24 (.A(n_28), .ZN(n_26));
   NAND3_X1 i_25 (.A1(b[1]), .A2(a[3]), .A3(n_36), .ZN(n_28));
   AOI22_X1 i_26 (.A1(b[0]), .A2(a[3]), .B1(b[1]), .B2(a[2]), .ZN(n_29));
   NOR2_X1 i_27 (.A1(n_37), .A2(n_30), .ZN(i[1]));
   AOI22_X1 i_28 (.A1(b[1]), .A2(a[0]), .B1(b[0]), .B2(a[1]), .ZN(n_30));
   XNOR2_X1 i_29 (.A(n_38), .B(n_31), .ZN(i[2]));
   XOR2_X1 i_30 (.A(n_36), .B(n_32), .Z(n_31));
   NOR2_X1 i_31 (.A1(n_11), .A2(n_33), .ZN(n_32));
   AOI22_X1 i_32 (.A1(b[1]), .A2(a[1]), .B1(b[2]), .B2(a[0]), .ZN(n_33));
   AND3_X1 i_33 (.A1(b[1]), .A2(a[0]), .A3(n_34), .ZN(n_11));
   INV_X1 i_34 (.A(n_35), .ZN(n_34));
   NAND2_X1 i_35 (.A1(b[2]), .A2(a[1]), .ZN(n_35));
   AND2_X1 i_36 (.A1(b[0]), .A2(a[2]), .ZN(n_36));
   INV_X1 i_37 (.A(n_38), .ZN(n_37));
   NAND3_X1 i_38 (.A1(b[1]), .A2(a[1]), .A3(i[0]), .ZN(n_38));
   AND2_X1 i_39 (.A1(b[0]), .A2(a[0]), .ZN(i[0]));
endmodule

module int_multiplier__parameterized0(a, b, enbl, c);
   input [15:0]a;
   input [2:0]b;
   input enbl;
   output [15:0]c;

   datapath__0_5921 i_0 (.b(b), .a({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      uc_0, uc_1, uc_2, a[5], a[4], a[3], a[2], a[1], a[0]}), .i({uc_3, uc_4, 
      uc_5, uc_6, uc_7, uc_8, uc_9, c[8], c[7], c[6], c[5], c[4], c[3], c[2], 
      c[1], c[0]}));
endmodule

module full_adder__4_312(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   INV_X1 i_3 (.A(b), .ZN(f));
endmodule

module full_adder__4_308(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(b), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(b), .ZN(cout));
endmodule

module full_adder__4_304(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XNOR2_X1 i_0_0 (.A(b), .B(cin), .ZN(f));
   OR2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(cout));
endmodule

module full_adder__4_300(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XNOR2_X1 i_0_0 (.A(b), .B(cin), .ZN(f));
   OR2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(cout));
endmodule

module full_adder__4_296(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(b), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(b), .ZN(cout));
endmodule

module full_adder__4_292(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XNOR2_X1 i_0_0 (.A(b), .B(cin), .ZN(f));
   OR2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(cout));
endmodule

module full_adder__4_288(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XNOR2_X1 i_0_0 (.A(b), .B(cin), .ZN(f));
   OR2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(cout));
endmodule

module full_adder__4_284(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XNOR2_X1 i_0_0 (.A(b), .B(cin), .ZN(f));
   OR2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(cout));
endmodule

module full_adder__4_280(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(b), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(b), .ZN(cout));
endmodule

module int_adder__parameterized3__4_317(a, b, cin, enbl, c, cout);
   input [15:0]a;
   input [15:0]b;
   input cin;
   input enbl;
   output [15:0]c;
   output cout;

   full_adder__4_312 full_adder_0_1_full_adder_0_i (.a(), .b(b[1]), .cin(), 
      .f(c[1]), .cout());
   full_adder__4_308 full_adder_0_2_full_adder_0_i (.a(), .b(b[2]), .cin(b[1]), 
      .f(c[2]), .cout(n_2));
   full_adder__4_304 full_adder_0_3_full_adder_0_i (.a(), .b(b[3]), .cin(n_2), 
      .f(c[3]), .cout(n_3));
   full_adder__4_300 full_adder_0_4_full_adder_0_i (.a(), .b(b[4]), .cin(n_3), 
      .f(c[4]), .cout(n_4));
   full_adder__4_296 full_adder_0_5_full_adder_0_i (.a(), .b(b[5]), .cin(n_4), 
      .f(c[5]), .cout(n_5));
   full_adder__4_292 full_adder_0_6_full_adder_0_i (.a(), .b(b[6]), .cin(n_5), 
      .f(c[6]), .cout(n_6));
   full_adder__4_288 full_adder_0_7_full_adder_0_i (.a(), .b(b[7]), .cin(n_6), 
      .f(c[7]), .cout(n_0));
   full_adder__4_284 full_adder_0_8_full_adder_0_i (.a(), .b(b[8]), .cin(n_0), 
      .f(c[8]), .cout(n_1));
   full_adder__4_280 full_adder_0_9_full_adder_0_i (.a(), .b(b[9]), .cin(n_1), 
      .f(c[9]), .cout(c[10]));
endmodule

module full_adder__4_440(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   INV_X1 i_3 (.A(b), .ZN(f));
endmodule

module full_adder__4_436(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XNOR2_X1 i_0_0 (.A(b), .B(cin), .ZN(f));
   OR2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(cout));
endmodule

module full_adder__4_432(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(b), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(b), .ZN(cout));
endmodule

module full_adder__4_428(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XNOR2_X1 i_0_0 (.A(b), .B(cin), .ZN(f));
   OR2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(cout));
endmodule

module full_adder__4_424(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   INV_X1 i_3 (.A(cin), .ZN(f));
endmodule

module int_adder__parameterized4__4_449(a, b, cin, enbl, c, cout);
   input [15:0]a;
   input [5:0]b;
   input cin;
   input enbl;
   output [15:0]c;
   output cout;

   full_adder__4_440 full_adder_0_2_full_adder_0_i (.a(), .b(b[2]), .cin(), 
      .f(c[2]), .cout());
   full_adder__4_436 full_adder_0_3_full_adder_0_i (.a(), .b(b[3]), .cin(b[2]), 
      .f(c[3]), .cout(n_0));
   full_adder__4_432 full_adder_0_4_full_adder_0_i (.a(), .b(b[4]), .cin(n_0), 
      .f(c[4]), .cout(n_1));
   full_adder__4_428 full_adder_0_5_full_adder_0_i (.a(), .b(b[5]), .cin(n_1), 
      .f(c[5]), .cout(c[7]));
   full_adder__4_424 full_adder_0_6_full_adder_0_i (.a(), .b(), .cin(c[7]), 
      .f(c[6]), .cout());
endmodule

module full_adder__4_76(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   INV_X1 i_3 (.A(b), .ZN(f));
endmodule

module full_adder__4_80(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(b), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(b), .ZN(cout));
endmodule

module full_adder__4_84(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XNOR2_X1 i_0_0 (.A(b), .B(cin), .ZN(f));
   OR2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(cout));
endmodule

module full_adder__4_88(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(b), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(b), .ZN(cout));
endmodule

module int_adder__parameterized4(a, b, cin, enbl, c, cout);
   input [15:0]a;
   input [5:0]b;
   input cin;
   input enbl;
   output [15:0]c;
   output cout;

   full_adder__4_76 full_adder_0_2_full_adder_0_i (.a(), .b(b[2]), .cin(), 
      .f(c[2]), .cout());
   full_adder__4_80 full_adder_0_3_full_adder_0_i (.a(), .b(b[3]), .cin(b[2]), 
      .f(c[3]), .cout(n_0));
   full_adder__4_84 full_adder_0_4_full_adder_0_i (.a(), .b(b[4]), .cin(n_0), 
      .f(c[4]), .cout(n_1));
   full_adder__4_88 full_adder_0_5_full_adder_0_i (.a(), .b(b[5]), .cin(n_1), 
      .f(c[5]), .cout(c[6]));
endmodule

module datapath__4_383(to_int6153, to_int, i);
   input [16:0]to_int6153;
   input [16:0]to_int;
   output [31:0]i;

   HA_X1 i_164 (.A(n_60), .B(n_59), .CO(n_1), .S(n_0));
   FA_X1 i_179 (.A(n_58), .B(n_53), .CI(n_52), .CO(n_3), .S(n_2));
   HA_X1 i_180 (.A(n_51), .B(n_1), .CO(n_5), .S(n_4));
   FA_X1 i_203 (.A(n_50), .B(n_47), .CI(n_45), .CO(n_7), .S(n_6));
   HA_X1 i_204 (.A(n_5), .B(n_3), .CO(n_9), .S(n_8));
   FA_X1 i_227 (.A(n_48), .B(n_46), .CI(n_44), .CO(n_11), .S(n_10));
   FA_X1 i_228 (.A(n_43), .B(n_49), .CI(n_9), .CO(n_13), .S(n_12));
   HA_X1 i_229 (.A(n_10), .B(n_7), .CO(n_15), .S(n_14));
   FA_X1 i_253 (.A(n_42), .B(n_11), .CI(n_15), .CO(n_17), .S(n_16));
   HA_X1 i_254 (.A(n_13), .B(n_41), .CO(n_19), .S(n_18));
   FA_X1 i_286 (.A(1'b0), .B(n_38), .CI(n_37), .CO(n_21), .S(n_20));
   HA_X1 i_287 (.A(n_19), .B(n_17), .CO(n_23), .S(n_22));
   FA_X1 i_320 (.A(1'b0), .B(n_40), .CI(n_39), .CO(n_55), .S(n_54));
   HA_X1 i_321 (.A(n_23), .B(n_21), .CO(n_57), .S(n_56));
   HA_X1 i_355 (.A(n_57), .B(n_55), .CO(n_114), .S(n_113));
   FA_X1 i_522 (.A(n_36), .B(n_35), .CI(n_34), .CO(n_24), .S(i[3]));
   FA_X1 i_523 (.A(n_33), .B(n_0), .CI(n_24), .CO(n_25), .S(i[4]));
   FA_X1 i_524 (.A(n_4), .B(n_2), .CI(n_25), .CO(n_26), .S(i[5]));
   FA_X1 i_525 (.A(n_8), .B(n_6), .CI(n_26), .CO(n_27), .S(i[6]));
   FA_X1 i_526 (.A(n_12), .B(n_14), .CI(n_27), .CO(n_28), .S(i[7]));
   FA_X1 i_527 (.A(n_16), .B(n_18), .CI(n_28), .CO(n_29), .S(i[8]));
   FA_X1 i_528 (.A(n_22), .B(n_20), .CI(n_29), .CO(n_30), .S(i[9]));
   FA_X1 i_529 (.A(n_56), .B(n_54), .CI(n_30), .CO(n_31), .S(i[10]));
   FA_X1 i_530 (.A(1'b0), .B(n_113), .CI(n_31), .CO(n_32), .S(i[11]));
   XNOR2_X1 i_0 (.A(n_101), .B(n_61), .ZN(n_33));
   NOR2_X1 i_1 (.A1(n_96), .A2(n_94), .ZN(n_61));
   OAI21_X1 i_2 (.A(n_109), .B1(n_104), .B2(to_int6153[2]), .ZN(n_34));
   XNOR2_X1 i_3 (.A(n_99), .B(n_62), .ZN(n_35));
   NOR2_X1 i_4 (.A1(n_102), .A2(n_100), .ZN(n_62));
   XOR2_X1 i_5 (.A(n_107), .B(n_92), .Z(n_36));
   OAI22_X1 i_6 (.A1(n_65), .A2(n_68), .B1(n_72), .B2(n_67), .ZN(n_37));
   NOR2_X1 i_7 (.A1(n_63), .A2(n_39), .ZN(n_38));
   AND3_X1 i_8 (.A1(to_int6153[4]), .A2(to_int[4]), .A3(n_40), .ZN(n_39));
   AND2_X1 i_9 (.A1(to_int6153[5]), .A2(to_int[5]), .ZN(n_40));
   AOI22_X1 i_10 (.A1(to_int6153[4]), .A2(to_int[5]), .B1(to_int[4]), .B2(
      to_int6153[5]), .ZN(n_63));
   XNOR2_X1 i_11 (.A(n_68), .B(n_64), .ZN(n_41));
   NOR2_X1 i_12 (.A1(n_66), .A2(n_65), .ZN(n_64));
   AOI22_X1 i_13 (.A1(to_int6153[3]), .A2(to_int[5]), .B1(to_int[4]), .B2(
      to_int6153[4]), .ZN(n_65));
   NOR2_X1 i_14 (.A1(n_72), .A2(n_67), .ZN(n_66));
   NAND2_X1 i_15 (.A1(to_int6153[4]), .A2(to_int[5]), .ZN(n_67));
   NAND2_X1 i_16 (.A1(to_int6153[5]), .A2(to_int[3]), .ZN(n_68));
   AND2_X1 i_17 (.A1(n_71), .A2(n_69), .ZN(n_42));
   OAI21_X1 i_18 (.A(n_73), .B1(n_72), .B2(n_81), .ZN(n_69));
   XNOR2_X1 i_19 (.A(n_73), .B(n_70), .ZN(n_43));
   XOR2_X1 i_20 (.A(n_81), .B(n_72), .Z(n_70));
   NAND2_X1 i_21 (.A1(n_81), .A2(n_72), .ZN(n_71));
   NAND2_X1 i_22 (.A1(to_int6153[3]), .A2(to_int[4]), .ZN(n_72));
   NAND2_X1 i_23 (.A1(to_int6153[4]), .A2(to_int[3]), .ZN(n_73));
   OAI22_X1 i_24 (.A1(n_79), .A2(n_82), .B1(n_91), .B2(n_81), .ZN(n_44));
   NOR2_X1 i_25 (.A1(n_46), .A2(n_74), .ZN(n_45));
   NOR2_X1 i_26 (.A1(n_76), .A2(n_75), .ZN(n_74));
   AND2_X1 i_27 (.A1(n_76), .A2(n_75), .ZN(n_46));
   OAI22_X1 i_28 (.A1(n_88), .A2(n_93), .B1(n_98), .B2(n_90), .ZN(n_75));
   OAI22_X1 i_29 (.A1(n_84), .A2(n_86), .B1(n_95), .B2(n_101), .ZN(n_76));
   XOR2_X1 i_30 (.A(n_95), .B(n_77), .Z(n_47));
   NOR2_X1 i_31 (.A1(n_95), .A2(n_77), .ZN(n_48));
   AND2_X1 i_32 (.A1(to_int6153[5]), .A2(to_int[2]), .ZN(n_49));
   NAND2_X1 i_33 (.A1(to_int6153[5]), .A2(to_int[1]), .ZN(n_77));
   XNOR2_X1 i_34 (.A(n_82), .B(n_78), .ZN(n_50));
   NOR2_X1 i_35 (.A1(n_80), .A2(n_79), .ZN(n_78));
   AOI22_X1 i_36 (.A1(to_int6153[1]), .A2(to_int[5]), .B1(to_int[4]), .B2(
      to_int6153[2]), .ZN(n_79));
   NOR2_X1 i_37 (.A1(n_91), .A2(n_81), .ZN(n_80));
   NAND2_X1 i_38 (.A1(to_int6153[2]), .A2(to_int[5]), .ZN(n_81));
   NAND2_X1 i_39 (.A1(to_int6153[3]), .A2(to_int[3]), .ZN(n_82));
   XNOR2_X1 i_40 (.A(n_86), .B(n_83), .ZN(n_51));
   NOR2_X1 i_41 (.A1(n_85), .A2(n_84), .ZN(n_83));
   AOI22_X1 i_42 (.A1(to_int6153[3]), .A2(to_int[2]), .B1(to_int[1]), .B2(
      to_int6153[4]), .ZN(n_84));
   NOR2_X1 i_43 (.A1(n_101), .A2(n_95), .ZN(n_85));
   NAND2_X1 i_44 (.A1(to_int6153[5]), .A2(to_int[0]), .ZN(n_86));
   XNOR2_X1 i_45 (.A(n_93), .B(n_87), .ZN(n_52));
   NOR2_X1 i_46 (.A1(n_89), .A2(n_88), .ZN(n_87));
   AOI22_X1 i_47 (.A1(to_int6153[0]), .A2(to_int[5]), .B1(to_int[4]), .B2(
      to_int6153[1]), .ZN(n_88));
   NOR2_X1 i_48 (.A1(n_98), .A2(n_90), .ZN(n_89));
   NAND2_X1 i_49 (.A1(to_int6153[1]), .A2(to_int[5]), .ZN(n_90));
   AOI21_X1 i_50 (.A(n_92), .B1(n_91), .B2(n_107), .ZN(n_53));
   NAND2_X1 i_51 (.A1(to_int6153[1]), .A2(to_int[4]), .ZN(n_91));
   NAND2_X1 i_52 (.A1(to_int6153[0]), .A2(to_int[3]), .ZN(n_92));
   NAND2_X1 i_53 (.A1(to_int6153[2]), .A2(to_int[3]), .ZN(n_93));
   OAI22_X1 i_54 (.A1(n_96), .A2(n_101), .B1(n_111), .B2(n_95), .ZN(n_58));
   NOR2_X1 i_55 (.A1(n_111), .A2(n_95), .ZN(n_94));
   NAND2_X1 i_56 (.A1(to_int6153[4]), .A2(to_int[2]), .ZN(n_95));
   AOI22_X1 i_57 (.A1(to_int6153[2]), .A2(to_int[2]), .B1(to_int[0]), .B2(
      to_int6153[4]), .ZN(n_96));
   XOR2_X1 i_58 (.A(n_98), .B(n_97), .Z(n_59));
   OAI211_X1 i_59 (.A(to_int6153[1]), .B(to_int[3]), .C1(n_104), .C2(n_119), 
      .ZN(n_97));
   NAND2_X1 i_60 (.A1(to_int6153[0]), .A2(to_int[4]), .ZN(n_98));
   OAI22_X1 i_61 (.A1(n_102), .A2(n_99), .B1(n_101), .B2(n_111), .ZN(n_60));
   NAND2_X1 i_62 (.A1(to_int6153[1]), .A2(to_int[2]), .ZN(n_99));
   NOR2_X1 i_63 (.A1(n_111), .A2(n_101), .ZN(n_100));
   NAND2_X1 i_64 (.A1(to_int6153[3]), .A2(to_int[1]), .ZN(n_101));
   AOI22_X1 i_65 (.A1(to_int6153[2]), .A2(to_int[1]), .B1(to_int[0]), .B2(
      to_int6153[3]), .ZN(n_102));
   NOR2_X1 i_66 (.A1(n_105), .A2(n_103), .ZN(i[1]));
   INV_X1 i_67 (.A(n_104), .ZN(n_103));
   NAND4_X1 i_68 (.A1(to_int6153[1]), .A2(to_int6153[0]), .A3(to_int[1]), 
      .A4(to_int[0]), .ZN(n_104));
   AOI22_X1 i_69 (.A1(to_int6153[0]), .A2(to_int[1]), .B1(to_int[0]), .B2(
      to_int6153[1]), .ZN(n_105));
   NOR3_X1 i_70 (.A1(n_112), .A2(n_108), .A3(n_106), .ZN(i[2]));
   AOI21_X1 i_71 (.A(to_int6153[0]), .B1(n_110), .B2(n_107), .ZN(n_106));
   OR2_X1 i_72 (.A1(n_117), .A2(n_111), .ZN(n_107));
   AOI21_X1 i_73 (.A(n_109), .B1(to_int[0]), .B2(n_119), .ZN(n_108));
   NAND3_X1 i_74 (.A1(n_110), .A2(to_int[2]), .A3(to_int6153[0]), .ZN(n_109));
   NAND2_X1 i_75 (.A1(n_117), .A2(n_111), .ZN(n_110));
   NAND2_X1 i_76 (.A1(to_int6153[2]), .A2(to_int[0]), .ZN(n_111));
   AOI21_X1 i_77 (.A(to_int[2]), .B1(n_116), .B2(n_115), .ZN(n_112));
   NAND2_X1 i_78 (.A1(i[0]), .A2(n_119), .ZN(n_115));
   AND2_X1 i_79 (.A1(to_int6153[0]), .A2(to_int[0]), .ZN(i[0]));
   NAND2_X1 i_80 (.A1(n_118), .A2(n_117), .ZN(n_116));
   NAND2_X1 i_81 (.A1(to_int6153[1]), .A2(to_int[1]), .ZN(n_117));
   INV_X1 i_82 (.A(to_int[0]), .ZN(n_118));
   INV_X1 i_83 (.A(to_int6153[2]), .ZN(n_119));
endmodule

module int_multiplier__4_384(a, b, enbl, c);
   input [15:0]a;
   input [15:0]b;
   input enbl;
   output [15:0]c;

   datapath__4_383 i_0 (.to_int6153({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, uc_0, uc_1, 
      uc_2, uc_3, uc_4, uc_5, b[5], b[4], b[3], b[2], b[1], b[0]}), .to_int({
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, uc_6, uc_7, uc_8, uc_9, uc_10, uc_11, a[5], 
      a[4], a[3], a[2], a[1], a[0]}), .i({uc_12, uc_13, uc_14, uc_15, uc_16, 
      uc_17, uc_18, uc_19, uc_20, uc_21, uc_22, uc_23, uc_24, uc_25, uc_26, 
      uc_27, uc_28, uc_29, uc_30, uc_31, c[11], c[10], c[9], c[8], c[7], c[6], 
      c[5], c[4], c[3], c[2], c[1], c[0]}));
endmodule

module full_adder__4_373(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   INV_X1 i_3 (.A(b), .ZN(f));
endmodule

module full_adder__4_369(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XNOR2_X1 i_0_0 (.A(b), .B(cin), .ZN(f));
   OR2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(cout));
endmodule

module full_adder__4_365(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(b), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(b), .ZN(cout));
endmodule

module full_adder__4_361(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(b), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(b), .ZN(cout));
endmodule

module full_adder__4_357(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(b), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(b), .ZN(cout));
endmodule

module full_adder__4_353(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XNOR2_X1 i_0_0 (.A(b), .B(cin), .ZN(f));
   OR2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(cout));
endmodule

module full_adder__4_349(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XNOR2_X1 i_0_0 (.A(b), .B(cin), .ZN(f));
   OR2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(cout));
endmodule

module full_adder__4_345(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XNOR2_X1 i_0_0 (.A(b), .B(cin), .ZN(f));
   OR2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(cout));
endmodule

module full_adder__4_341(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(b), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(b), .ZN(cout));
endmodule

module full_adder__4_337(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XOR2_X1 i_0_0 (.A(b), .B(cin), .Z(f));
   AND2_X1 i_0_1 (.A1(cin), .A2(b), .ZN(cout));
endmodule

module full_adder__4_333(a, b, cin, f, cout);
   input a;
   input b;
   input cin;
   output f;
   output cout;

   XNOR2_X1 i_0_0 (.A(b), .B(cin), .ZN(f));
   OR2_X1 i_0_1 (.A1(b), .A2(cin), .ZN(cout));
endmodule

module int_adder__parameterized3__4_382(a, b, cin, enbl, c, cout);
   input [15:0]a;
   input [15:0]b;
   input cin;
   input enbl;
   output [15:0]c;
   output cout;

   full_adder__4_373 full_adder_0_2_full_adder_0_i (.a(), .b(b[2]), .cin(), 
      .f(c[2]), .cout());
   full_adder__4_369 full_adder_0_3_full_adder_0_i (.a(), .b(b[3]), .cin(b[2]), 
      .f(c[3]), .cout(n_3));
   full_adder__4_365 full_adder_0_4_full_adder_0_i (.a(), .b(b[4]), .cin(n_3), 
      .f(c[4]), .cout(n_4));
   full_adder__4_361 full_adder_0_5_full_adder_0_i (.a(), .b(b[5]), .cin(n_4), 
      .f(c[5]), .cout(n_5));
   full_adder__4_357 full_adder_0_6_full_adder_0_i (.a(), .b(b[6]), .cin(n_5), 
      .f(c[6]), .cout(n_6));
   full_adder__4_353 full_adder_0_7_full_adder_0_i (.a(), .b(b[7]), .cin(n_6), 
      .f(c[7]), .cout(n_7));
   full_adder__4_349 full_adder_0_8_full_adder_0_i (.a(), .b(b[8]), .cin(n_7), 
      .f(c[8]), .cout(n_8));
   full_adder__4_345 full_adder_0_9_full_adder_0_i (.a(), .b(b[9]), .cin(n_8), 
      .f(c[9]), .cout(n_0));
   full_adder__4_341 full_adder_0_10_full_adder_0_i (.a(), .b(b[10]), .cin(n_0), 
      .f(c[10]), .cout(n_1));
   full_adder__4_337 full_adder_0_11_full_adder_0_i (.a(), .b(b[11]), .cin(n_1), 
      .f(c[11]), .cout(n_2));
   full_adder__4_333 full_adder_0_12_full_adder_0_i (.a(), .b(b[12]), .cin(n_2), 
      .f(c[12]), .cout(c[13]));
endmodule

module datapath__0_5915(to_int6153, to_int, i);
   input [16:0]to_int6153;
   input [16:0]to_int;
   output [31:0]i;

   HA_X1 i_164 (.A(n_46), .B(n_44), .CO(n_1), .S(n_0));
   FA_X1 i_179 (.A(n_43), .B(n_42), .CI(n_41), .CO(n_3), .S(n_2));
   HA_X1 i_180 (.A(n_41), .B(n_1), .CO(n_5), .S(n_4));
   FA_X1 i_203 (.A(n_36), .B(n_37), .CI(1'b0), .CO(n_7), .S(n_6));
   HA_X1 i_204 (.A(n_5), .B(n_3), .CO(n_9), .S(n_8));
   FA_X1 i_227 (.A(n_38), .B(n_35), .CI(n_34), .CO(n_11), .S(n_10));
   HA_X1 i_229 (.A(n_10), .B(n_7), .CO(n_13), .S(n_12));
   FA_X1 i_253 (.A(n_33), .B(n_11), .CI(n_13), .CO(n_15), .S(n_14));
   HA_X1 i_254 (.A(n_39), .B(to_int6153[4]), .CO(n_17), .S(n_16));
   HA_X1 i_287 (.A(n_17), .B(n_15), .CO(n_19), .S(n_18));
   FA_X1 i_320 (.A(1'b0), .B(to_int6153[5]), .CI(n_40), .CO(n_56), .S(n_55));
   FA_X1 i_522 (.A(n_31), .B(n_45), .CI(n_30), .CO(n_20), .S(i[3]));
   FA_X1 i_523 (.A(n_29), .B(n_0), .CI(n_20), .CO(n_21), .S(i[4]));
   FA_X1 i_524 (.A(n_4), .B(n_2), .CI(n_21), .CO(n_22), .S(i[5]));
   FA_X1 i_525 (.A(n_8), .B(n_6), .CI(n_22), .CO(n_23), .S(i[6]));
   FA_X1 i_526 (.A(n_9), .B(n_12), .CI(n_23), .CO(n_24), .S(i[7]));
   FA_X1 i_527 (.A(n_14), .B(n_16), .CI(n_24), .CO(n_25), .S(i[8]));
   FA_X1 i_528 (.A(n_18), .B(n_32), .CI(n_25), .CO(n_26), .S(i[9]));
   FA_X1 i_529 (.A(n_19), .B(n_55), .CI(n_26), .CO(n_27), .S(i[10]));
   FA_X1 i_530 (.A(1'b0), .B(n_56), .CI(n_27), .CO(n_28), .S(i[11]));
   XNOR2_X1 i_0 (.A(n_62), .B(n_57), .ZN(n_29));
   AOI21_X1 i_1 (.A(n_64), .B1(n_65), .B2(n_62), .ZN(n_30));
   OAI33_X1 i_2 (.A1(n_64), .A2(n_63), .A3(n_46), .B1(n_64), .B2(n_61), .B3(n_45), 
      .ZN(n_31));
   AND2_X1 i_3 (.A1(to_int6153[5]), .A2(to_int[3]), .ZN(n_32));
   AND2_X1 i_4 (.A1(to_int6153[4]), .A2(to_int[3]), .ZN(n_33));
   OAI21_X1 i_5 (.A(n_48), .B1(n_63), .B2(n_47), .ZN(n_34));
   OAI21_X1 i_6 (.A(n_50), .B1(n_53), .B2(n_52), .ZN(n_35));
   XNOR2_X1 i_7 (.A(n_63), .B(n_37), .ZN(n_36));
   NOR2_X1 i_8 (.A1(n_38), .A2(n_47), .ZN(n_37));
   AOI22_X1 i_9 (.A1(to_int6153[5]), .A2(to_int6153[1]), .B1(to_int6153[4]), 
      .B2(to_int[2]), .ZN(n_47));
   INV_X1 i_10 (.A(n_48), .ZN(n_38));
   NAND2_X1 i_11 (.A1(n_46), .A2(n_40), .ZN(n_48));
   AND2_X1 i_12 (.A1(to_int6153[5]), .A2(to_int[2]), .ZN(n_39));
   AND2_X1 i_13 (.A1(to_int6153[5]), .A2(to_int6153[4]), .ZN(n_40));
   XOR2_X1 i_14 (.A(n_53), .B(n_49), .Z(n_41));
   NAND2_X1 i_15 (.A1(n_51), .A2(n_50), .ZN(n_49));
   NAND3_X1 i_16 (.A1(to_int6153[5]), .A2(to_int6153[0]), .A3(n_59), .ZN(n_50));
   INV_X1 i_17 (.A(n_52), .ZN(n_51));
   AOI21_X1 i_18 (.A(n_59), .B1(to_int6153[5]), .B2(to_int6153[0]), .ZN(n_52));
   NAND2_X1 i_19 (.A1(to_int[3]), .A2(to_int[2]), .ZN(n_53));
   NAND2_X1 i_20 (.A1(n_58), .A2(n_54), .ZN(n_42));
   AOI21_X1 i_21 (.A(n_60), .B1(n_62), .B2(n_58), .ZN(n_43));
   XNOR2_X1 i_22 (.A(n_57), .B(n_54), .ZN(n_44));
   NAND2_X1 i_23 (.A1(n_46), .A2(n_45), .ZN(n_54));
   AOI21_X1 i_24 (.A(n_60), .B1(n_59), .B2(n_45), .ZN(n_57));
   NAND2_X1 i_25 (.A1(n_59), .A2(n_45), .ZN(n_58));
   NOR2_X1 i_26 (.A1(n_64), .A2(n_63), .ZN(n_45));
   AND2_X1 i_27 (.A1(to_int6153[4]), .A2(to_int6153[1]), .ZN(n_59));
   AOI22_X1 i_28 (.A1(to_int6153[4]), .A2(to_int6153[0]), .B1(to_int6153[1]), 
      .B2(to_int[3]), .ZN(n_60));
   INV_X1 i_29 (.A(n_61), .ZN(n_46));
   NAND2_X1 i_30 (.A1(to_int6153[1]), .A2(to_int[2]), .ZN(n_61));
   NOR2_X1 i_31 (.A1(n_65), .A2(to_int6153[0]), .ZN(i[2]));
   INV_X1 i_32 (.A(to_int[2]), .ZN(n_62));
   INV_X1 i_33 (.A(to_int[3]), .ZN(n_63));
   INV_X1 i_34 (.A(to_int6153[0]), .ZN(n_64));
   INV_X1 i_35 (.A(to_int6153[1]), .ZN(n_65));
endmodule

module int_multiplier(a, b, enbl, c);
   input [15:0]a;
   input [15:0]b;
   input enbl;
   output [15:0]c;

   datapath__0_5915 i_0 (.to_int6153({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, uc_0, uc_1, 
      uc_2, uc_3, uc_4, uc_5, a[5], a[4], uc_6, uc_7, a[1], a[0]}), .to_int({
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, 
      uc_14, uc_15, a[3], a[2], uc_16, uc_17}), .i({uc_18, uc_19, uc_20, uc_21, 
      uc_22, uc_23, uc_24, uc_25, uc_26, uc_27, uc_28, uc_29, uc_30, uc_31, 
      uc_32, uc_33, uc_34, uc_35, uc_36, uc_37, c[11], c[10], c[9], c[8], c[7], 
      c[6], c[5], c[4], c[3], c[2], uc_38, uc_39}));
endmodule

module next_adr(in_data, enbl, clk, rst, out_adr, done, state_test);
   input [31:0]in_data;
   input enbl;
   input clk;
   input rst;
   output [15:0]out_adr;
   output done;
   output [3:0]state_test;

   wire [15:0]new_adr;
   wire [15:0]hdr_tsize_m;
   wire [15:0]max_us_adr;
   wire [15:0]max_u0_adr;
   wire [15:0]max_x_adr;
   wire [15:0]hdr_n_m;
   wire [15:0]max_b_adr;
   wire [15:0]hdr_n_square;
   wire [25:20]i;
   wire [18:17]fpu_mode;
   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_166;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_180;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_190;
   wire n_0_191;
   wire n_0_192;
   wire n_0_193;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_200;
   wire n_0_201;
   wire n_0_202;
   wire n_0_203;
   wire n_0_204;

   int_adder__parameterized2 iterator (.a(out_adr), .b({n_69, fpu_mode[17]}), 
      .cin(), .enbl(), .c(new_adr), .cout());
   int_multiplier__parameterized0 max_us_adr_mul (.a({uc_0, uc_1, uc_2, uc_3, 
      uc_4, uc_5, uc_6, uc_7, uc_8, uc_9, i[25], i[24], i[23], i[22], i[21], 
      i[20]}), .b({n_27, n_28, n_29}), .enbl(), .c({uc_10, uc_11, uc_12, uc_13, 
      uc_14, uc_15, uc_16, hdr_tsize_m[8], hdr_tsize_m[7], hdr_tsize_m[6], 
      hdr_tsize_m[5], hdr_tsize_m[4], hdr_tsize_m[3], hdr_tsize_m[2], 
      hdr_tsize_m[1], hdr_tsize_m[0]}));
   int_adder__parameterized3__4_317 max_us_adr_add (.a(), .b({uc_17, uc_18, 
      uc_19, uc_20, uc_21, uc_22, hdr_tsize_m[8], hdr_tsize_m[7], hdr_tsize_m[6], 
      hdr_tsize_m[5], hdr_tsize_m[4], hdr_tsize_m[3], hdr_tsize_m[2], 
      hdr_tsize_m[1], hdr_tsize_m[0], uc_23}), .cin(), .enbl(), .c({uc_24, uc_25, 
      uc_26, uc_27, uc_28, max_us_adr[10], max_us_adr[9], max_us_adr[8], 
      max_us_adr[7], max_us_adr[6], max_us_adr[5], max_us_adr[4], max_us_adr[3], 
      max_us_adr[2], max_us_adr[1], uc_29}), .cout());
   int_adder__parameterized4__4_449 max_u0_adr_add (.a(), .b({i[24], i[23], 
      i[22], i[21], uc_30, uc_31}), .cin(), .enbl(), .c({uc_32, uc_33, uc_34, 
      uc_35, uc_36, uc_37, uc_38, uc_39, max_u0_adr[7], max_u0_adr[6], 
      max_u0_adr[5], max_u0_adr[4], max_u0_adr[3], max_u0_adr[2], uc_40, uc_41}), 
      .cout());
   int_adder__parameterized4 max_x_adr_add (.a(), .b({n_22, n_23, n_24, n_25, 
      uc_42, uc_43}), .cin(), .enbl(), .c({uc_44, uc_45, uc_46, uc_47, uc_48, 
      uc_49, uc_50, uc_51, uc_52, max_x_adr[6], max_x_adr[5], max_x_adr[4], 
      max_x_adr[3], max_x_adr[2], uc_53, uc_54}), .cout());
   int_multiplier__4_384 max_b_adr_mul (.a({uc_55, uc_56, uc_57, uc_58, uc_59, 
      uc_60, uc_61, uc_62, uc_63, uc_64, n_21, n_22, n_23, n_24, n_25, n_26}), 
      .b({uc_65, uc_66, uc_67, uc_68, uc_69, uc_70, uc_71, uc_72, uc_73, uc_74, 
      i[25], i[24], i[23], i[22], i[21], i[20]}), .enbl(), .c({uc_75, uc_76, 
      uc_77, uc_78, hdr_n_m[11], hdr_n_m[10], hdr_n_m[9], hdr_n_m[8], hdr_n_m[7], 
      hdr_n_m[6], hdr_n_m[5], hdr_n_m[4], hdr_n_m[3], hdr_n_m[2], hdr_n_m[1], 
      hdr_n_m[0]}));
   int_adder__parameterized3__4_382 max_b_adr_add (.a(), .b({uc_79, uc_80, uc_81, 
      hdr_n_m[11], hdr_n_m[10], hdr_n_m[9], hdr_n_m[8], hdr_n_m[7], hdr_n_m[6], 
      hdr_n_m[5], hdr_n_m[4], hdr_n_m[3], hdr_n_m[2], hdr_n_m[1], uc_82, uc_83}), 
      .cin(), .enbl(), .c({uc_84, uc_85, max_b_adr[13], max_b_adr[12], 
      max_b_adr[11], max_b_adr[10], max_b_adr[9], max_b_adr[8], max_b_adr[7], 
      max_b_adr[6], max_b_adr[5], max_b_adr[4], max_b_adr[3], max_b_adr[2], 
      uc_86, uc_87}), .cout());
   int_multiplier max_a_adr_mul (.a({uc_88, uc_89, uc_90, uc_91, uc_92, uc_93, 
      uc_94, uc_95, uc_96, uc_97, n_21, n_22, n_23, n_24, n_25, n_26}), .b(), 
      .enbl(), .c({uc_98, uc_99, uc_100, uc_101, hdr_n_square[11], 
      hdr_n_square[10], hdr_n_square[9], hdr_n_square[8], hdr_n_square[7], 
      hdr_n_square[6], hdr_n_square[5], hdr_n_square[4], hdr_n_square[3], 
      hdr_n_square[2], uc_102, uc_103}));
   DFFR_X1 done_reg (.D(n_68), .RN(n_71), .CK(n_70), .Q(done), .QN());
   DFFS_X1 \cur_adr_reg[15]  (.D(n_67), .SN(n_71), .CK(n_70), .Q(n_0), .QN());
   DFFS_X1 \cur_adr_reg[14]  (.D(n_66), .SN(n_71), .CK(n_70), .Q(n_1), .QN());
   DFFS_X1 \cur_adr_reg[13]  (.D(n_65), .SN(n_71), .CK(n_70), .Q(n_2), .QN());
   DFFS_X1 \cur_adr_reg[12]  (.D(n_64), .SN(n_71), .CK(n_70), .Q(n_3), .QN());
   DFFS_X1 \cur_adr_reg[11]  (.D(n_63), .SN(n_71), .CK(n_70), .Q(n_4), .QN());
   DFFS_X1 \cur_adr_reg[10]  (.D(n_62), .SN(n_71), .CK(n_70), .Q(n_5), .QN());
   DFFS_X1 \cur_adr_reg[9]  (.D(n_61), .SN(n_71), .CK(n_70), .Q(n_6), .QN());
   DFFS_X1 \cur_adr_reg[8]  (.D(n_60), .SN(n_71), .CK(n_70), .Q(n_7), .QN());
   DFFS_X1 \cur_adr_reg[7]  (.D(n_59), .SN(n_71), .CK(n_70), .Q(n_8), .QN());
   DFFS_X1 \cur_adr_reg[6]  (.D(n_58), .SN(n_71), .CK(n_70), .Q(n_9), .QN());
   DFFS_X1 \cur_adr_reg[5]  (.D(n_57), .SN(n_71), .CK(n_70), .Q(n_10), .QN());
   DFFS_X1 \cur_adr_reg[4]  (.D(n_56), .SN(n_71), .CK(n_70), .Q(n_11), .QN());
   DFFS_X1 \cur_adr_reg[3]  (.D(n_55), .SN(n_71), .CK(n_70), .Q(n_12), .QN());
   DFFS_X1 \cur_adr_reg[2]  (.D(n_54), .SN(n_71), .CK(n_70), .Q(n_13), .QN());
   DFFS_X1 \cur_adr_reg[1]  (.D(n_52), .SN(n_71), .CK(n_70), .Q(n_14), .QN());
   DFFS_X1 \cur_adr_reg[0]  (.D(n_51), .SN(n_71), .CK(n_70), .Q(n_15), .QN());
   TBUF_X1 i_5 (.A(n_15), .EN(n_53), .Z(out_adr[0]));
   TBUF_X1 i_7 (.A(n_14), .EN(n_53), .Z(out_adr[1]));
   TBUF_X1 i_9 (.A(n_13), .EN(n_53), .Z(out_adr[2]));
   TBUF_X1 i_11 (.A(n_12), .EN(n_53), .Z(out_adr[3]));
   TBUF_X1 i_13 (.A(n_11), .EN(n_53), .Z(out_adr[4]));
   TBUF_X1 i_15 (.A(n_10), .EN(n_53), .Z(out_adr[5]));
   TBUF_X1 i_17 (.A(n_9), .EN(n_53), .Z(out_adr[6]));
   TBUF_X1 i_19 (.A(n_8), .EN(n_53), .Z(out_adr[7]));
   TBUF_X1 i_21 (.A(n_7), .EN(n_53), .Z(out_adr[8]));
   TBUF_X1 i_23 (.A(n_6), .EN(n_53), .Z(out_adr[9]));
   TBUF_X1 i_25 (.A(n_5), .EN(n_53), .Z(out_adr[10]));
   TBUF_X1 i_27 (.A(n_4), .EN(n_53), .Z(out_adr[11]));
   TBUF_X1 i_29 (.A(n_3), .EN(n_53), .Z(out_adr[12]));
   TBUF_X1 i_31 (.A(n_2), .EN(n_53), .Z(out_adr[13]));
   TBUF_X1 i_33 (.A(n_1), .EN(n_53), .Z(out_adr[14]));
   TBUF_X1 i_35 (.A(n_0), .EN(n_53), .Z(out_adr[15]));
   INV_X1 i_36 (.A(n_16), .ZN(n_53));
   DFFS_X1 i_39 (.D(n_50), .SN(n_71), .CK(n_70), .Q(n_16), .QN());
   DFFR_X1 \state_reg[3]  (.D(n_49), .RN(n_71), .CK(n_70), .Q(n_17), .QN());
   DFFR_X1 \state_reg[2]  (.D(n_48), .RN(n_71), .CK(n_70), .Q(n_18), .QN());
   DFFR_X1 \state_reg[1]  (.D(n_47), .RN(n_71), .CK(n_70), .Q(n_19), .QN());
   DFFR_X1 \state_reg[0]  (.D(n_46), .RN(n_71), .CK(n_70), .Q(n_20), .QN());
   DFF_X1 \header_reg[31]  (.D(n_45), .CK(n_70), .Q(n_21), .QN());
   DFF_X1 \header_reg[30]  (.D(n_44), .CK(n_70), .Q(n_22), .QN());
   DFF_X1 \header_reg[29]  (.D(n_43), .CK(n_70), .Q(n_23), .QN());
   DFF_X1 \header_reg[28]  (.D(n_42), .CK(n_70), .Q(n_24), .QN());
   DFF_X1 \header_reg[27]  (.D(n_41), .CK(n_70), .Q(n_25), .QN());
   DFF_X1 \header_reg[26]  (.D(n_40), .CK(n_70), .Q(n_26), .QN());
   DFF_X1 \header_reg[25]  (.D(n_39), .CK(n_70), .Q(i[25]), .QN());
   DFF_X1 \header_reg[24]  (.D(n_38), .CK(n_70), .Q(i[24]), .QN());
   DFF_X1 \header_reg[23]  (.D(n_37), .CK(n_70), .Q(i[23]), .QN());
   DFF_X1 \header_reg[22]  (.D(n_36), .CK(n_70), .Q(i[22]), .QN());
   DFF_X1 \header_reg[21]  (.D(n_35), .CK(n_70), .Q(i[21]), .QN());
   DFF_X1 \header_reg[20]  (.D(n_34), .CK(n_70), .Q(i[20]), .QN());
   DFF_X1 \header_reg[17]  (.D(n_33), .CK(n_70), .Q(fpu_mode[17]), .QN());
   DFF_X1 \header_reg[16]  (.D(n_32), .CK(n_70), .Q(n_27), .QN());
   DFF_X1 \header_reg[15]  (.D(n_31), .CK(n_70), .Q(n_28), .QN());
   DFF_X1 \header_reg[14]  (.D(n_30), .CK(n_70), .Q(n_29), .QN());
   MUX2_X1 i_0_0 (.A(n_29), .B(in_data[14]), .S(n_0_1), .Z(n_30));
   MUX2_X1 i_0_1 (.A(n_28), .B(in_data[15]), .S(n_0_1), .Z(n_31));
   MUX2_X1 i_0_2 (.A(n_27), .B(in_data[16]), .S(n_0_1), .Z(n_32));
   OAI21_X1 i_0_3 (.A(n_0_0), .B1(n_0_1), .B2(n_69), .ZN(n_33));
   NAND2_X1 i_0_4 (.A1(in_data[17]), .A2(n_0_1), .ZN(n_0_0));
   MUX2_X1 i_0_5 (.A(i[20]), .B(in_data[20]), .S(n_0_1), .Z(n_34));
   MUX2_X1 i_0_6 (.A(i[21]), .B(in_data[21]), .S(n_0_1), .Z(n_35));
   MUX2_X1 i_0_7 (.A(i[22]), .B(in_data[22]), .S(n_0_1), .Z(n_36));
   MUX2_X1 i_0_8 (.A(i[23]), .B(in_data[23]), .S(n_0_1), .Z(n_37));
   MUX2_X1 i_0_9 (.A(i[24]), .B(in_data[24]), .S(n_0_1), .Z(n_38));
   MUX2_X1 i_0_10 (.A(i[25]), .B(in_data[25]), .S(n_0_1), .Z(n_39));
   MUX2_X1 i_0_11 (.A(n_26), .B(in_data[26]), .S(n_0_1), .Z(n_40));
   MUX2_X1 i_0_12 (.A(n_25), .B(in_data[27]), .S(n_0_1), .Z(n_41));
   MUX2_X1 i_0_13 (.A(n_24), .B(in_data[28]), .S(n_0_1), .Z(n_42));
   MUX2_X1 i_0_14 (.A(n_23), .B(in_data[29]), .S(n_0_1), .Z(n_43));
   MUX2_X1 i_0_15 (.A(n_22), .B(in_data[30]), .S(n_0_1), .Z(n_44));
   MUX2_X1 i_0_16 (.A(n_21), .B(in_data[31]), .S(n_0_1), .Z(n_45));
   NOR4_X1 i_0_17 (.A1(n_0_175), .A2(n_0_173), .A3(n_20), .A4(rst), .ZN(n_0_1));
   OAI211_X1 i_0_18 (.A(n_0_10), .B(n_0_8), .C1(n_0_2), .C2(n_20), .ZN(n_46));
   OAI21_X1 i_0_19 (.A(n_0_202), .B1(n_0_75), .B2(n_0_3), .ZN(n_0_2));
   NOR3_X1 i_0_20 (.A1(n_0_5), .A2(n_0_4), .A3(new_adr[13]), .ZN(n_0_3));
   NAND3_X1 i_0_21 (.A1(new_adr[2]), .A2(n_0_164), .A3(n_0_155), .ZN(n_0_4));
   NAND4_X1 i_0_22 (.A1(new_adr[0]), .A2(n_0_196), .A3(n_0_7), .A4(n_0_6), 
      .ZN(n_0_5));
   NOR4_X1 i_0_23 (.A1(new_adr[12]), .A2(new_adr[10]), .A3(new_adr[9]), .A4(
      new_adr[1]), .ZN(n_0_6));
   NOR4_X1 i_0_24 (.A1(new_adr[8]), .A2(new_adr[6]), .A3(new_adr[4]), .A4(n_18), 
      .ZN(n_0_7));
   AOI22_X1 i_0_25 (.A1(n_0_176), .A2(n_0_9), .B1(n_0_76), .B2(n_0_78), .ZN(
      n_0_8));
   OAI22_X1 i_0_26 (.A1(n_0_179), .A2(n_0_174), .B1(n_0_173), .B2(n_20), 
      .ZN(n_0_9));
   OAI21_X1 i_0_27 (.A(n_20), .B1(n_0_11), .B2(n_0_173), .ZN(n_0_10));
   OAI21_X1 i_0_28 (.A(n_0_12), .B1(n_0_143), .B2(n_0_199), .ZN(n_0_11));
   NAND2_X1 i_0_29 (.A1(n_0_24), .A2(n_0_199), .ZN(n_0_12));
   AOI21_X1 i_0_30 (.A(n_0_13), .B1(n_0_16), .B2(n_0_121), .ZN(n_47));
   OAI22_X1 i_0_31 (.A1(n_0_14), .A2(n_0_199), .B1(n_19), .B2(n_0_170), .ZN(
      n_0_13));
   INV_X1 i_0_32 (.A(n_0_15), .ZN(n_0_14));
   OAI21_X1 i_0_33 (.A(n_0_70), .B1(n_0_147), .B2(n_0_203), .ZN(n_0_15));
   NOR3_X1 i_0_34 (.A1(n_0_203), .A2(n_18), .A3(n_0_198), .ZN(n_0_16));
   NAND2_X1 i_0_35 (.A1(n_0_67), .A2(n_0_17), .ZN(n_48));
   OAI21_X1 i_0_36 (.A(n_18), .B1(n_0_148), .B2(n_0_72), .ZN(n_0_17));
   OAI21_X1 i_0_37 (.A(n_0_200), .B1(n_0_147), .B2(n_0_18), .ZN(n_49));
   NAND3_X1 i_0_38 (.A1(n_18), .A2(n_20), .A3(enbl), .ZN(n_0_18));
   AOI21_X1 i_0_39 (.A(n_0_172), .B1(n_0_85), .B2(n_0_197), .ZN(n_50));
   INV_X1 i_0_40 (.A(n_0_19), .ZN(n_51));
   AOI222_X1 i_0_41 (.A1(n_0_23), .A2(n_0_170), .B1(n_15), .B2(n_0_85), .C1(
      n_0_52), .C2(new_adr[0]), .ZN(n_0_19));
   OAI21_X1 i_0_42 (.A(n_0_20), .B1(n_0_147), .B2(n_0_169), .ZN(n_52));
   AOI22_X1 i_0_43 (.A1(n_0_21), .A2(new_adr[1]), .B1(n_14), .B2(n_0_85), 
      .ZN(n_0_20));
   OAI211_X1 i_0_44 (.A(n_0_87), .B(n_0_22), .C1(n_0_23), .C2(n_0_203), .ZN(
      n_0_21));
   AOI21_X1 i_0_45 (.A(n_0_204), .B1(n_0_141), .B2(n_0_131), .ZN(n_0_22));
   OAI21_X1 i_0_46 (.A(n_0_144), .B1(n_0_24), .B2(n_18), .ZN(n_0_23));
   NOR2_X1 i_0_47 (.A1(n_0_121), .A2(n_0_198), .ZN(n_0_24));
   NAND3_X1 i_0_48 (.A1(n_0_53), .A2(n_0_26), .A3(n_0_25), .ZN(n_54));
   AOI21_X1 i_0_49 (.A(n_0_38), .B1(n_0_85), .B2(n_13), .ZN(n_0_25));
   OAI21_X1 i_0_50 (.A(new_adr[2]), .B1(n_0_139), .B2(n_0_27), .ZN(n_0_26));
   OAI211_X1 i_0_51 (.A(n_0_59), .B(n_0_28), .C1(n_19), .C2(n_0_171), .ZN(n_0_27));
   NAND2_X1 i_0_52 (.A1(n_0_90), .A2(n_0_78), .ZN(n_0_28));
   NAND3_X1 i_0_53 (.A1(n_0_50), .A2(n_0_30), .A3(n_0_29), .ZN(n_55));
   NAND2_X1 i_0_54 (.A1(n_12), .A2(n_0_85), .ZN(n_0_29));
   NAND2_X1 i_0_55 (.A1(n_0_31), .A2(new_adr[3]), .ZN(n_0_30));
   NAND3_X1 i_0_56 (.A1(n_0_169), .A2(n_0_88), .A3(n_0_138), .ZN(n_0_31));
   NAND3_X1 i_0_57 (.A1(n_0_74), .A2(n_0_33), .A3(n_0_32), .ZN(n_56));
   AOI21_X1 i_0_58 (.A(n_0_45), .B1(n_0_85), .B2(n_11), .ZN(n_0_32));
   NAND2_X1 i_0_59 (.A1(n_0_34), .A2(new_adr[4]), .ZN(n_0_33));
   NAND3_X1 i_0_60 (.A1(n_0_142), .A2(n_0_36), .A3(n_0_35), .ZN(n_0_34));
   OAI211_X1 i_0_61 (.A(n_19), .B(n_0_202), .C1(n_0_122), .C2(n_18), .ZN(n_0_35));
   NAND3_X1 i_0_62 (.A1(n_0_175), .A2(n_0_37), .A3(n_0_202), .ZN(n_0_36));
   NAND2_X1 i_0_63 (.A1(n_0_49), .A2(n_20), .ZN(n_0_37));
   OAI21_X1 i_0_64 (.A(n_0_39), .B1(n_0_144), .B2(n_0_169), .ZN(n_57));
   NOR2_X1 i_0_65 (.A1(n_0_169), .A2(n_0_144), .ZN(n_0_38));
   AOI22_X1 i_0_66 (.A1(n_0_40), .A2(new_adr[5]), .B1(n_10), .B2(n_0_85), 
      .ZN(n_0_39));
   NAND4_X1 i_0_67 (.A1(n_0_119), .A2(n_0_59), .A3(n_0_42), .A4(n_0_41), 
      .ZN(n_0_40));
   NAND3_X1 i_0_68 (.A1(n_0_90), .A2(n_0_131), .A3(n_19), .ZN(n_0_41));
   OR2_X1 i_0_69 (.A1(n_0_64), .A2(n_19), .ZN(n_0_42));
   NAND3_X1 i_0_70 (.A1(n_0_43), .A2(n_0_62), .A3(n_0_73), .ZN(n_58));
   AOI22_X1 i_0_71 (.A1(n_9), .A2(n_0_85), .B1(n_0_63), .B2(new_adr[6]), 
      .ZN(n_0_43));
   NAND4_X1 i_0_72 (.A1(n_0_67), .A2(n_0_62), .A3(n_0_46), .A4(n_0_44), .ZN(n_59));
   AOI21_X1 i_0_73 (.A(n_0_45), .B1(n_0_85), .B2(n_8), .ZN(n_0_44));
   NOR2_X1 i_0_74 (.A1(n_0_169), .A2(n_0_147), .ZN(n_0_45));
   OAI21_X1 i_0_75 (.A(new_adr[7]), .B1(n_0_47), .B2(n_0_204), .ZN(n_0_46));
   OAI211_X1 i_0_76 (.A(n_0_140), .B(n_0_48), .C1(n_0_49), .C2(n_0_203), 
      .ZN(n_0_47));
   NAND2_X1 i_0_77 (.A1(n_0_94), .A2(n_0_78), .ZN(n_0_48));
   NAND2_X1 i_0_78 (.A1(n_0_151), .A2(n_18), .ZN(n_0_49));
   NAND3_X1 i_0_79 (.A1(n_0_50), .A2(n_0_74), .A3(n_0_51), .ZN(n_60));
   AND2_X1 i_0_80 (.A1(n_0_73), .A2(n_0_67), .ZN(n_0_50));
   AOI22_X1 i_0_81 (.A1(n_0_52), .A2(new_adr[8]), .B1(n_7), .B2(n_0_85), 
      .ZN(n_0_51));
   OAI21_X1 i_0_82 (.A(n_0_142), .B1(n_0_173), .B2(n_0_176), .ZN(n_0_52));
   NAND3_X1 i_0_83 (.A1(n_0_53), .A2(n_0_54), .A3(n_0_55), .ZN(n_61));
   AOI21_X1 i_0_84 (.A(n_0_66), .B1(n_0_75), .B2(n_0_78), .ZN(n_0_53));
   NAND2_X1 i_0_85 (.A1(n_6), .A2(n_0_85), .ZN(n_0_54));
   OAI21_X1 i_0_86 (.A(new_adr[9]), .B1(n_0_71), .B2(n_0_60), .ZN(n_0_55));
   NAND2_X1 i_0_87 (.A1(n_0_57), .A2(n_0_56), .ZN(n_62));
   AOI22_X1 i_0_88 (.A1(n_5), .A2(n_0_85), .B1(n_0_78), .B2(n_0_75), .ZN(n_0_56));
   OAI21_X1 i_0_89 (.A(new_adr[10]), .B1(n_0_60), .B2(n_0_58), .ZN(n_0_57));
   OAI21_X1 i_0_90 (.A(n_0_119), .B1(n_0_59), .B2(n_0_198), .ZN(n_0_58));
   NAND3_X1 i_0_91 (.A1(n_0_148), .A2(n_0_170), .A3(n_18), .ZN(n_0_59));
   OAI22_X1 i_0_92 (.A1(n_0_76), .A2(n_0_77), .B1(n_0_171), .B2(n_0_70), 
      .ZN(n_0_60));
   NAND3_X1 i_0_93 (.A1(n_0_61), .A2(n_0_62), .A3(n_0_73), .ZN(n_63));
   AOI22_X1 i_0_94 (.A1(n_4), .A2(n_0_85), .B1(n_0_63), .B2(new_adr[11]), 
      .ZN(n_0_61));
   NAND2_X1 i_0_95 (.A1(n_0_78), .A2(n_0_76), .ZN(n_0_62));
   NAND3_X1 i_0_96 (.A1(n_0_142), .A2(n_0_82), .A3(n_0_64), .ZN(n_0_63));
   OAI211_X1 i_0_97 (.A(n_18), .B(n_0_202), .C1(n_0_94), .C2(n_20), .ZN(n_0_64));
   NAND2_X1 i_0_98 (.A1(n_0_68), .A2(n_0_65), .ZN(n_64));
   AOI21_X1 i_0_99 (.A(n_0_66), .B1(n_0_85), .B2(n_3), .ZN(n_0_65));
   INV_X1 i_0_100 (.A(n_0_67), .ZN(n_0_66));
   NAND4_X1 i_0_101 (.A1(n_19), .A2(n_0_170), .A3(n_0_121), .A4(n_0_199), 
      .ZN(n_0_67));
   OAI21_X1 i_0_102 (.A(new_adr[12]), .B1(n_0_71), .B2(n_0_69), .ZN(n_0_68));
   OAI21_X1 i_0_103 (.A(n_0_87), .B1(n_0_70), .B2(n_0_169), .ZN(n_0_69));
   NAND2_X1 i_0_104 (.A1(n_0_198), .A2(n_0_151), .ZN(n_0_70));
   OAI21_X1 i_0_105 (.A(n_0_138), .B1(n_0_149), .B2(n_0_72), .ZN(n_0_71));
   NAND2_X1 i_0_106 (.A1(n_19), .A2(n_0_170), .ZN(n_0_72));
   NAND4_X1 i_0_107 (.A1(n_0_80), .A2(n_0_79), .A3(n_0_74), .A4(n_0_73), 
      .ZN(n_65));
   NAND3_X1 i_0_108 (.A1(n_0_143), .A2(n_0_170), .A3(n_18), .ZN(n_0_73));
   OAI21_X1 i_0_109 (.A(n_0_78), .B1(n_0_76), .B2(n_0_75), .ZN(n_0_74));
   NOR2_X1 i_0_110 (.A1(n_0_94), .A2(n_19), .ZN(n_0_75));
   NOR2_X1 i_0_111 (.A1(n_0_198), .A2(n_0_90), .ZN(n_0_76));
   INV_X1 i_0_112 (.A(n_0_78), .ZN(n_0_77));
   NOR2_X1 i_0_113 (.A1(n_0_171), .A2(n_20), .ZN(n_0_78));
   NAND2_X1 i_0_114 (.A1(n_2), .A2(n_0_85), .ZN(n_0_79));
   NAND2_X1 i_0_115 (.A1(n_0_81), .A2(new_adr[13]), .ZN(n_0_80));
   NAND3_X1 i_0_116 (.A1(n_0_171), .A2(n_0_142), .A3(n_0_82), .ZN(n_0_81));
   NAND2_X1 i_0_117 (.A1(n_0_120), .A2(n_19), .ZN(n_0_82));
   INV_X1 i_0_118 (.A(n_0_83), .ZN(n_66));
   AOI22_X1 i_0_119 (.A1(n_0_86), .A2(new_adr[14]), .B1(n_1), .B2(n_0_85), 
      .ZN(n_0_83));
   INV_X1 i_0_120 (.A(n_0_84), .ZN(n_67));
   AOI22_X1 i_0_121 (.A1(n_0_86), .A2(new_adr[15]), .B1(n_0), .B2(n_0_85), 
      .ZN(n_0_84));
   OAI21_X1 i_0_122 (.A(enbl), .B1(n_0_176), .B2(n_0_200), .ZN(n_0_85));
   OAI211_X1 i_0_123 (.A(n_0_119), .B(n_0_87), .C1(n_0_169), .C2(n_0_143), 
      .ZN(n_0_86));
   OR2_X1 i_0_124 (.A1(n_0_88), .A2(n_20), .ZN(n_0_87));
   OR2_X1 i_0_125 (.A1(n_0_173), .A2(n_0_89), .ZN(n_0_88));
   AOI22_X1 i_0_126 (.A1(n_0_94), .A2(n_0_93), .B1(n_0_90), .B2(n_19), .ZN(
      n_0_89));
   NAND4_X1 i_0_127 (.A1(n_0_115), .A2(n_0_92), .A3(n_0_91), .A4(n_0_117), 
      .ZN(n_0_90));
   NOR4_X1 i_0_128 (.A1(n_0_165), .A2(n_0_118), .A3(n_0_116), .A4(n_0_112), 
      .ZN(n_0_91));
   NOR2_X1 i_0_129 (.A1(n_0_114), .A2(n_0_113), .ZN(n_0_92));
   NOR2_X1 i_0_130 (.A1(n_0_199), .A2(n_19), .ZN(n_0_93));
   NAND3_X1 i_0_131 (.A1(n_0_97), .A2(n_0_96), .A3(n_0_95), .ZN(n_0_94));
   NOR4_X1 i_0_132 (.A1(n_0_110), .A2(n_0_108), .A3(n_0_106), .A4(n_0_101), 
      .ZN(n_0_95));
   NOR4_X1 i_0_133 (.A1(n_0_111), .A2(n_0_107), .A3(n_0_103), .A4(n_0_99), 
      .ZN(n_0_96));
   NOR3_X1 i_0_134 (.A1(n_0_195), .A2(n_0_105), .A3(n_0_98), .ZN(n_0_97));
   NAND4_X1 i_0_135 (.A1(n_0_109), .A2(n_0_104), .A3(n_0_102), .A4(n_0_100), 
      .ZN(n_0_98));
   XOR2_X1 i_0_136 (.A(new_adr[4]), .B(max_b_adr[4]), .Z(n_0_99));
   XNOR2_X1 i_0_137 (.A(new_adr[13]), .B(max_b_adr[13]), .ZN(n_0_100));
   XOR2_X1 i_0_138 (.A(new_adr[1]), .B(hdr_n_m[0]), .Z(n_0_101));
   XNOR2_X1 i_0_139 (.A(new_adr[10]), .B(max_b_adr[10]), .ZN(n_0_102));
   XOR2_X1 i_0_140 (.A(new_adr[5]), .B(max_b_adr[5]), .Z(n_0_103));
   XNOR2_X1 i_0_141 (.A(new_adr[8]), .B(max_b_adr[8]), .ZN(n_0_104));
   XOR2_X1 i_0_142 (.A(new_adr[2]), .B(max_b_adr[2]), .Z(n_0_105));
   XOR2_X1 i_0_143 (.A(new_adr[7]), .B(max_b_adr[7]), .Z(n_0_106));
   XOR2_X1 i_0_144 (.A(new_adr[11]), .B(max_b_adr[11]), .Z(n_0_107));
   XOR2_X1 i_0_145 (.A(new_adr[6]), .B(max_b_adr[6]), .Z(n_0_108));
   XNOR2_X1 i_0_146 (.A(new_adr[3]), .B(max_b_adr[3]), .ZN(n_0_109));
   XOR2_X1 i_0_147 (.A(new_adr[9]), .B(max_b_adr[9]), .Z(n_0_110));
   XOR2_X1 i_0_148 (.A(new_adr[12]), .B(max_b_adr[12]), .Z(n_0_111));
   XOR2_X1 i_0_149 (.A(new_adr[2]), .B(max_u0_adr[2]), .Z(n_0_112));
   XOR2_X1 i_0_150 (.A(new_adr[7]), .B(max_u0_adr[7]), .Z(n_0_113));
   XOR2_X1 i_0_151 (.A(new_adr[3]), .B(max_u0_adr[3]), .Z(n_0_114));
   XNOR2_X1 i_0_152 (.A(new_adr[4]), .B(max_u0_adr[4]), .ZN(n_0_115));
   XOR2_X1 i_0_153 (.A(new_adr[6]), .B(max_u0_adr[6]), .Z(n_0_116));
   XNOR2_X1 i_0_154 (.A(new_adr[1]), .B(i[20]), .ZN(n_0_117));
   XOR2_X1 i_0_155 (.A(new_adr[5]), .B(max_u0_adr[5]), .Z(n_0_118));
   AOI21_X1 i_0_156 (.A(n_0_204), .B1(n_0_120), .B2(n_0_141), .ZN(n_0_119));
   AOI21_X1 i_0_157 (.A(n_0_173), .B1(n_0_121), .B2(n_20), .ZN(n_0_120));
   INV_X1 i_0_158 (.A(n_0_122), .ZN(n_0_121));
   NAND3_X1 i_0_159 (.A1(n_0_133), .A2(n_0_129), .A3(n_0_123), .ZN(n_0_122));
   NOR3_X1 i_0_160 (.A1(n_0_157), .A2(n_0_127), .A3(n_0_124), .ZN(n_0_123));
   NAND4_X1 i_0_161 (.A1(n_0_135), .A2(n_0_132), .A3(n_0_126), .A4(n_0_125), 
      .ZN(n_0_124));
   NOR4_X1 i_0_162 (.A1(n_0_136), .A2(n_0_134), .A3(n_0_130), .A4(n_0_128), 
      .ZN(n_0_125));
   XNOR2_X1 i_0_163 (.A(new_adr[9]), .B(hdr_n_square[8]), .ZN(n_0_126));
   NAND4_X1 i_0_164 (.A1(new_adr[2]), .A2(n_0_196), .A3(n_0_137), .A4(n_0_201), 
      .ZN(n_0_127));
   XOR2_X1 i_0_165 (.A(new_adr[11]), .B(hdr_n_square[10]), .Z(n_0_128));
   XNOR2_X1 i_0_166 (.A(new_adr[10]), .B(hdr_n_square[9]), .ZN(n_0_129));
   XOR2_X1 i_0_167 (.A(new_adr[12]), .B(hdr_n_square[11]), .Z(n_0_130));
   NOR2_X1 i_0_168 (.A1(n_0_173), .A2(n_20), .ZN(n_0_131));
   XNOR2_X1 i_0_169 (.A(new_adr[8]), .B(hdr_n_square[7]), .ZN(n_0_132));
   XNOR2_X1 i_0_170 (.A(new_adr[5]), .B(hdr_n_square[4]), .ZN(n_0_133));
   XOR2_X1 i_0_171 (.A(new_adr[6]), .B(hdr_n_square[5]), .Z(n_0_134));
   XNOR2_X1 i_0_172 (.A(new_adr[4]), .B(hdr_n_square[3]), .ZN(n_0_135));
   XOR2_X1 i_0_173 (.A(new_adr[3]), .B(hdr_n_square[2]), .Z(n_0_136));
   XNOR2_X1 i_0_174 (.A(new_adr[7]), .B(hdr_n_square[6]), .ZN(n_0_137));
   INV_X1 i_0_175 (.A(n_0_139), .ZN(n_0_138));
   OAI21_X1 i_0_176 (.A(n_0_142), .B1(n_0_140), .B2(n_18), .ZN(n_0_139));
   NAND2_X1 i_0_177 (.A1(n_19), .A2(n_0_202), .ZN(n_0_140));
   NOR2_X1 i_0_178 (.A1(n_0_198), .A2(n_18), .ZN(n_0_141));
   OR3_X1 i_0_179 (.A1(n_0_175), .A2(n_0_174), .A3(n_20), .ZN(n_0_142));
   NAND2_X1 i_0_180 (.A1(n_0_147), .A2(n_0_144), .ZN(n_0_143));
   OR4_X1 i_0_181 (.A1(n_0_157), .A2(n_0_153), .A3(n_0_145), .A4(n_19), .ZN(
      n_0_144));
   NAND2_X1 i_0_182 (.A1(new_adr[8]), .A2(n_0_146), .ZN(n_0_145));
   NOR2_X1 i_0_183 (.A1(n_0_168), .A2(n_0_152), .ZN(n_0_146));
   NAND2_X1 i_0_184 (.A1(n_19), .A2(n_0_149), .ZN(n_0_147));
   INV_X1 i_0_185 (.A(n_0_149), .ZN(n_0_148));
   NOR4_X1 i_0_186 (.A1(n_0_165), .A2(n_0_163), .A3(n_0_154), .A4(n_0_150), 
      .ZN(n_0_149));
   NAND4_X1 i_0_187 (.A1(new_adr[7]), .A2(new_adr[6]), .A3(new_adr[4]), .A4(
      n_0_164), .ZN(n_0_150));
   OR4_X1 i_0_188 (.A1(n_0_167), .A2(n_0_157), .A3(n_0_153), .A4(n_0_152), 
      .ZN(n_0_151));
   NAND4_X1 i_0_189 (.A1(n_0_159), .A2(n_0_155), .A3(new_adr[10]), .A4(
      new_adr[9]), .ZN(n_0_152));
   NAND4_X1 i_0_190 (.A1(n_0_162), .A2(n_0_161), .A3(n_0_160), .A4(n_0_156), 
      .ZN(n_0_153));
   XOR2_X1 i_0_191 (.A(new_adr[1]), .B(n_29), .Z(n_0_154));
   NOR2_X1 i_0_192 (.A1(new_adr[11]), .A2(new_adr[7]), .ZN(n_0_155));
   XNOR2_X1 i_0_193 (.A(new_adr[4]), .B(max_x_adr[4]), .ZN(n_0_156));
   NAND2_X1 i_0_194 (.A1(n_0_158), .A2(new_adr[0]), .ZN(n_0_157));
   XNOR2_X1 i_0_195 (.A(new_adr[1]), .B(n_26), .ZN(n_0_158));
   XNOR2_X1 i_0_196 (.A(new_adr[6]), .B(max_x_adr[6]), .ZN(n_0_159));
   XNOR2_X1 i_0_197 (.A(new_adr[2]), .B(max_x_adr[2]), .ZN(n_0_160));
   XNOR2_X1 i_0_198 (.A(new_adr[3]), .B(max_x_adr[3]), .ZN(n_0_161));
   XNOR2_X1 i_0_199 (.A(new_adr[5]), .B(max_x_adr[5]), .ZN(n_0_162));
   XOR2_X1 i_0_200 (.A(new_adr[2]), .B(n_28), .Z(n_0_163));
   NOR2_X1 i_0_201 (.A1(new_adr[5]), .A2(new_adr[3]), .ZN(n_0_164));
   OR4_X1 i_0_202 (.A1(n_0_167), .A2(n_0_166), .A3(new_adr[10]), .A4(new_adr[9]), 
      .ZN(n_0_165));
   NAND2_X1 i_0_203 (.A1(new_adr[11]), .A2(new_adr[0]), .ZN(n_0_166));
   NAND3_X1 i_0_204 (.A1(new_adr[8]), .A2(n_0_196), .A3(n_0_190), .ZN(n_0_167));
   NAND2_X1 i_0_205 (.A1(n_0_196), .A2(n_0_190), .ZN(n_0_168));
   NAND2_X1 i_0_206 (.A1(n_18), .A2(n_0_170), .ZN(n_0_169));
   AND2_X1 i_0_207 (.A1(n_20), .A2(n_0_202), .ZN(n_0_170));
   NAND2_X1 i_0_208 (.A1(n_18), .A2(n_0_202), .ZN(n_0_171));
   OR2_X1 i_0_209 (.A1(done), .A2(n_0_172), .ZN(n_68));
   NOR3_X1 i_0_210 (.A1(n_0_177), .A2(n_0_175), .A3(n_0_174), .ZN(n_0_172));
   NAND2_X1 i_0_211 (.A1(n_0_200), .A2(enbl), .ZN(n_0_173));
   NAND2_X1 i_0_212 (.A1(n_17), .A2(enbl), .ZN(n_0_174));
   NAND2_X1 i_0_213 (.A1(n_0_199), .A2(n_0_198), .ZN(n_0_175));
   NOR2_X1 i_0_214 (.A1(n_18), .A2(n_19), .ZN(n_0_176));
   NOR2_X1 i_0_215 (.A1(n_20), .A2(n_0_178), .ZN(n_0_177));
   INV_X1 i_0_216 (.A(n_0_179), .ZN(n_0_178));
   NAND3_X1 i_0_217 (.A1(n_0_186), .A2(n_0_182), .A3(n_0_180), .ZN(n_0_179));
   NOR3_X1 i_0_218 (.A1(n_0_181), .A2(n_0_193), .A3(n_0_191), .ZN(n_0_180));
   NAND3_X1 i_0_219 (.A1(new_adr[11]), .A2(n_0_190), .A3(n_0_189), .ZN(n_0_181));
   NOR4_X1 i_0_220 (.A1(n_0_195), .A2(n_0_185), .A3(n_0_184), .A4(n_0_183), 
      .ZN(n_0_182));
   XOR2_X1 i_0_221 (.A(max_us_adr[6]), .B(new_adr[6]), .Z(n_0_183));
   XOR2_X1 i_0_222 (.A(max_us_adr[2]), .B(new_adr[2]), .Z(n_0_184));
   XOR2_X1 i_0_223 (.A(max_us_adr[10]), .B(new_adr[10]), .Z(n_0_185));
   NOR4_X1 i_0_224 (.A1(n_0_194), .A2(n_0_192), .A3(n_0_188), .A4(n_0_187), 
      .ZN(n_0_186));
   XOR2_X1 i_0_225 (.A(max_us_adr[5]), .B(new_adr[5]), .Z(n_0_187));
   XOR2_X1 i_0_226 (.A(max_us_adr[8]), .B(new_adr[8]), .Z(n_0_188));
   XNOR2_X1 i_0_227 (.A(max_us_adr[1]), .B(new_adr[1]), .ZN(n_0_189));
   NOR2_X1 i_0_228 (.A1(n_0_201), .A2(new_adr[12]), .ZN(n_0_190));
   XOR2_X1 i_0_229 (.A(max_us_adr[4]), .B(new_adr[4]), .Z(n_0_191));
   XOR2_X1 i_0_230 (.A(max_us_adr[7]), .B(new_adr[7]), .Z(n_0_192));
   XOR2_X1 i_0_231 (.A(max_us_adr[9]), .B(new_adr[9]), .Z(n_0_193));
   XOR2_X1 i_0_232 (.A(max_us_adr[3]), .B(new_adr[3]), .Z(n_0_194));
   NAND2_X1 i_0_233 (.A1(new_adr[0]), .A2(n_0_196), .ZN(n_0_195));
   NOR2_X1 i_0_234 (.A1(new_adr[15]), .A2(new_adr[14]), .ZN(n_0_196));
   INV_X1 i_0_235 (.A(fpu_mode[17]), .ZN(n_69));
   INV_X1 i_0_236 (.A(n_16), .ZN(n_0_197));
   INV_X1 i_0_237 (.A(clk), .ZN(n_70));
   INV_X1 i_0_238 (.A(rst), .ZN(n_71));
   INV_X1 i_0_239 (.A(n_19), .ZN(n_0_198));
   INV_X1 i_0_240 (.A(n_18), .ZN(n_0_199));
   INV_X1 i_0_241 (.A(n_17), .ZN(n_0_200));
   INV_X1 i_0_242 (.A(new_adr[13]), .ZN(n_0_201));
   INV_X1 i_0_243 (.A(n_0_173), .ZN(n_0_202));
   INV_X1 i_0_244 (.A(n_0_170), .ZN(n_0_203));
   INV_X1 i_0_245 (.A(n_0_142), .ZN(n_0_204));
endmodule

module io(in_state, clk, rst, cpu_data, in_data, adr, interrupt, error_success);
   input [1:0]in_state;
   input clk;
   input rst;
   inout [31:0]cpu_data;
   inout [31:0]in_data;
   output [15:0]adr;
   output interrupt;
   output error_success;

   wire dcm_error_success;
   wire [31:0]dcm_out_data;
   wire dcm_out_ready;
   wire nau_done;
   wire [15:0]nau_out_adr;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_0_7;
   wire n_0_0_8;
   wire n_0_0;
   wire n_0_0_11;
   wire to_std_logic;
   wire n_0_0_16;
   wire n_0_0_12;
   wire n_0_0_9;
   wire n_0_0_10;
   wire n_0_0_13;
   wire n_0_21;
   wire n_0_1;
   wire n_0_0_15;
   wire n_0_0_17;
   wire n_0_88;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_0_18;
   wire n_0_0_19;
   wire n_0_20;
   wire n_0_0_14;
   wire n_0_0_20;
   wire n_0_0_21;
   wire n_0_0_22;
   wire n_0_0_23;

   decompressor decompressor (.in_data(cpu_data), .rst(rst), .enbl_in(
      to_std_logic), .clk(clk), .state_wait(n_0), .out_ready(dcm_out_ready), 
      .out_data(dcm_out_data), .error_success(dcm_error_success), .buf_test());
   next_adr nau (.in_data({dcm_out_data[31], dcm_out_data[30], dcm_out_data[29], 
      dcm_out_data[28], dcm_out_data[27], dcm_out_data[26], dcm_out_data[25], 
      dcm_out_data[24], dcm_out_data[23], dcm_out_data[22], dcm_out_data[21], 
      dcm_out_data[20], uc_0, uc_1, dcm_out_data[17], dcm_out_data[16], 
      dcm_out_data[15], dcm_out_data[14], uc_2, uc_3, uc_4, uc_5, uc_6, uc_7, 
      uc_8, uc_9, uc_10, uc_11, uc_12, uc_13, uc_14, uc_15}), .enbl(
      dcm_out_ready), .clk(clk), .rst(rst), .out_adr(nau_out_adr), .done(
      nau_done), .state_test());
   DLH_X1 \adr_reg[15]  (.D(nau_out_adr[15]), .G(n_0_20), .Q(n_0_2));
   DLH_X1 \adr_reg[14]  (.D(nau_out_adr[14]), .G(n_0_20), .Q(n_0_3));
   DLH_X1 \adr_reg[13]  (.D(nau_out_adr[13]), .G(n_0_20), .Q(n_0_4));
   DLH_X1 \adr_reg[12]  (.D(nau_out_adr[12]), .G(n_0_20), .Q(n_0_5));
   DLH_X1 \adr_reg[11]  (.D(nau_out_adr[11]), .G(n_0_20), .Q(n_0_6));
   DLH_X1 \adr_reg[10]  (.D(nau_out_adr[10]), .G(n_0_20), .Q(n_0_7));
   DLH_X1 \adr_reg[9]  (.D(nau_out_adr[9]), .G(n_0_20), .Q(n_0_8));
   DLH_X1 \adr_reg[8]  (.D(nau_out_adr[8]), .G(n_0_20), .Q(n_0_9));
   DLH_X1 \adr_reg[7]  (.D(nau_out_adr[7]), .G(n_0_20), .Q(n_0_10));
   DLH_X1 \adr_reg[6]  (.D(nau_out_adr[6]), .G(n_0_20), .Q(n_0_11));
   DLH_X1 \adr_reg[5]  (.D(nau_out_adr[5]), .G(n_0_20), .Q(n_0_12));
   DLH_X1 \adr_reg[4]  (.D(nau_out_adr[4]), .G(n_0_20), .Q(n_0_13));
   DLH_X1 \adr_reg[3]  (.D(nau_out_adr[3]), .G(n_0_20), .Q(n_0_14));
   DLH_X1 \adr_reg[2]  (.D(nau_out_adr[2]), .G(n_0_20), .Q(n_0_15));
   DLH_X1 \adr_reg[1]  (.D(nau_out_adr[1]), .G(n_0_20), .Q(n_0_16));
   DLH_X1 \adr_reg[0]  (.D(nau_out_adr[0]), .G(n_0_20), .Q(n_0_17));
   TBUF_X1 i_0_5 (.A(n_0_17), .EN(n_0_18), .Z(adr[0]));
   TBUF_X1 i_0_7 (.A(n_0_16), .EN(n_0_18), .Z(adr[1]));
   TBUF_X1 i_0_9 (.A(n_0_15), .EN(n_0_18), .Z(adr[2]));
   TBUF_X1 i_0_11 (.A(n_0_14), .EN(n_0_18), .Z(adr[3]));
   TBUF_X1 i_0_13 (.A(n_0_13), .EN(n_0_18), .Z(adr[4]));
   TBUF_X1 i_0_15 (.A(n_0_12), .EN(n_0_18), .Z(adr[5]));
   TBUF_X1 i_0_17 (.A(n_0_11), .EN(n_0_18), .Z(adr[6]));
   TBUF_X1 i_0_19 (.A(n_0_10), .EN(n_0_18), .Z(adr[7]));
   TBUF_X1 i_0_21 (.A(n_0_9), .EN(n_0_18), .Z(adr[8]));
   TBUF_X1 i_0_23 (.A(n_0_8), .EN(n_0_18), .Z(adr[9]));
   TBUF_X1 i_0_25 (.A(n_0_7), .EN(n_0_18), .Z(adr[10]));
   TBUF_X1 i_0_27 (.A(n_0_6), .EN(n_0_18), .Z(adr[11]));
   TBUF_X1 i_0_29 (.A(n_0_5), .EN(n_0_18), .Z(adr[12]));
   TBUF_X1 i_0_31 (.A(n_0_4), .EN(n_0_18), .Z(adr[13]));
   TBUF_X1 i_0_33 (.A(n_0_3), .EN(n_0_18), .Z(adr[14]));
   TBUF_X1 i_0_35 (.A(n_0_2), .EN(n_0_18), .Z(adr[15]));
   INV_X1 i_0_36 (.A(n_0_19), .ZN(n_0_18));
   DLH_X1 i_0_37 (.D(n_0_21), .G(n_0_20), .Q(n_0_19));
   DLH_X1 \cpu_data_reg[31]  (.D(n_0_87), .G(n_0_88), .Q(n_0_22));
   DLH_X1 \cpu_data_reg[30]  (.D(n_0_86), .G(n_0_88), .Q(n_0_23));
   DLH_X1 \cpu_data_reg[29]  (.D(n_0_85), .G(n_0_88), .Q(n_0_24));
   DLH_X1 \cpu_data_reg[28]  (.D(n_0_84), .G(n_0_88), .Q(n_0_25));
   DLH_X1 \cpu_data_reg[27]  (.D(n_0_83), .G(n_0_88), .Q(n_0_26));
   DLH_X1 \cpu_data_reg[26]  (.D(n_0_82), .G(n_0_88), .Q(n_0_27));
   DLH_X1 \cpu_data_reg[25]  (.D(n_0_81), .G(n_0_88), .Q(n_0_28));
   DLH_X1 \cpu_data_reg[24]  (.D(n_0_80), .G(n_0_88), .Q(n_0_29));
   DLH_X1 \cpu_data_reg[23]  (.D(n_0_79), .G(n_0_88), .Q(n_0_30));
   DLH_X1 \cpu_data_reg[22]  (.D(n_0_78), .G(n_0_88), .Q(n_0_31));
   DLH_X1 \cpu_data_reg[21]  (.D(n_0_77), .G(n_0_88), .Q(n_0_32));
   DLH_X1 \cpu_data_reg[20]  (.D(n_0_76), .G(n_0_88), .Q(n_0_33));
   DLH_X1 \cpu_data_reg[19]  (.D(n_0_75), .G(n_0_88), .Q(n_0_34));
   DLH_X1 \cpu_data_reg[18]  (.D(n_0_74), .G(n_0_88), .Q(n_0_35));
   DLH_X1 \cpu_data_reg[17]  (.D(n_0_73), .G(n_0_88), .Q(n_0_36));
   DLH_X1 \cpu_data_reg[16]  (.D(n_0_72), .G(n_0_88), .Q(n_0_37));
   DLH_X1 \cpu_data_reg[15]  (.D(n_0_71), .G(n_0_88), .Q(n_0_38));
   DLH_X1 \cpu_data_reg[14]  (.D(n_0_70), .G(n_0_88), .Q(n_0_39));
   DLH_X1 \cpu_data_reg[13]  (.D(n_0_69), .G(n_0_88), .Q(n_0_40));
   DLH_X1 \cpu_data_reg[12]  (.D(n_0_68), .G(n_0_88), .Q(n_0_41));
   DLH_X1 \cpu_data_reg[11]  (.D(n_0_67), .G(n_0_88), .Q(n_0_42));
   DLH_X1 \cpu_data_reg[10]  (.D(n_0_66), .G(n_0_88), .Q(n_0_43));
   DLH_X1 \cpu_data_reg[9]  (.D(n_0_65), .G(n_0_88), .Q(n_0_44));
   DLH_X1 \cpu_data_reg[8]  (.D(n_0_64), .G(n_0_88), .Q(n_0_45));
   DLH_X1 \cpu_data_reg[7]  (.D(n_0_63), .G(n_0_88), .Q(n_0_46));
   DLH_X1 \cpu_data_reg[6]  (.D(n_0_62), .G(n_0_88), .Q(n_0_47));
   DLH_X1 \cpu_data_reg[5]  (.D(n_0_61), .G(n_0_88), .Q(n_0_48));
   DLH_X1 \cpu_data_reg[4]  (.D(n_0_60), .G(n_0_88), .Q(n_0_49));
   DLH_X1 \cpu_data_reg[3]  (.D(n_0_59), .G(n_0_88), .Q(n_0_50));
   DLH_X1 \cpu_data_reg[2]  (.D(n_0_58), .G(n_0_88), .Q(n_0_51));
   DLH_X1 \cpu_data_reg[1]  (.D(n_0_57), .G(n_0_88), .Q(n_0_52));
   DLH_X1 \cpu_data_reg[0]  (.D(n_0_56), .G(n_0_88), .Q(n_0_53));
   TBUF_X1 i_0_55 (.A(n_0_53), .EN(n_0_54), .Z(cpu_data[0]));
   TBUF_X1 i_0_57 (.A(n_0_52), .EN(n_0_54), .Z(cpu_data[1]));
   TBUF_X1 i_0_59 (.A(n_0_51), .EN(n_0_54), .Z(cpu_data[2]));
   TBUF_X1 i_0_61 (.A(n_0_50), .EN(n_0_54), .Z(cpu_data[3]));
   TBUF_X1 i_0_63 (.A(n_0_49), .EN(n_0_54), .Z(cpu_data[4]));
   TBUF_X1 i_0_65 (.A(n_0_48), .EN(n_0_54), .Z(cpu_data[5]));
   TBUF_X1 i_0_67 (.A(n_0_47), .EN(n_0_54), .Z(cpu_data[6]));
   TBUF_X1 i_0_69 (.A(n_0_46), .EN(n_0_54), .Z(cpu_data[7]));
   TBUF_X1 i_0_71 (.A(n_0_45), .EN(n_0_54), .Z(cpu_data[8]));
   TBUF_X1 i_0_73 (.A(n_0_44), .EN(n_0_54), .Z(cpu_data[9]));
   TBUF_X1 i_0_75 (.A(n_0_43), .EN(n_0_54), .Z(cpu_data[10]));
   TBUF_X1 i_0_77 (.A(n_0_42), .EN(n_0_54), .Z(cpu_data[11]));
   TBUF_X1 i_0_79 (.A(n_0_41), .EN(n_0_54), .Z(cpu_data[12]));
   TBUF_X1 i_0_81 (.A(n_0_40), .EN(n_0_54), .Z(cpu_data[13]));
   TBUF_X1 i_0_83 (.A(n_0_39), .EN(n_0_54), .Z(cpu_data[14]));
   TBUF_X1 i_0_85 (.A(n_0_38), .EN(n_0_54), .Z(cpu_data[15]));
   TBUF_X1 i_0_87 (.A(n_0_37), .EN(n_0_54), .Z(cpu_data[16]));
   TBUF_X1 i_0_89 (.A(n_0_36), .EN(n_0_54), .Z(cpu_data[17]));
   TBUF_X1 i_0_91 (.A(n_0_35), .EN(n_0_54), .Z(cpu_data[18]));
   TBUF_X1 i_0_93 (.A(n_0_34), .EN(n_0_54), .Z(cpu_data[19]));
   TBUF_X1 i_0_95 (.A(n_0_33), .EN(n_0_54), .Z(cpu_data[20]));
   TBUF_X1 i_0_97 (.A(n_0_32), .EN(n_0_54), .Z(cpu_data[21]));
   TBUF_X1 i_0_99 (.A(n_0_31), .EN(n_0_54), .Z(cpu_data[22]));
   TBUF_X1 i_0_101 (.A(n_0_30), .EN(n_0_54), .Z(cpu_data[23]));
   TBUF_X1 i_0_103 (.A(n_0_29), .EN(n_0_54), .Z(cpu_data[24]));
   TBUF_X1 i_0_105 (.A(n_0_28), .EN(n_0_54), .Z(cpu_data[25]));
   TBUF_X1 i_0_107 (.A(n_0_27), .EN(n_0_54), .Z(cpu_data[26]));
   TBUF_X1 i_0_109 (.A(n_0_26), .EN(n_0_54), .Z(cpu_data[27]));
   TBUF_X1 i_0_111 (.A(n_0_25), .EN(n_0_54), .Z(cpu_data[28]));
   TBUF_X1 i_0_113 (.A(n_0_24), .EN(n_0_54), .Z(cpu_data[29]));
   TBUF_X1 i_0_115 (.A(n_0_23), .EN(n_0_54), .Z(cpu_data[30]));
   TBUF_X1 i_0_117 (.A(n_0_22), .EN(n_0_54), .Z(cpu_data[31]));
   INV_X1 i_0_118 (.A(n_0_55), .ZN(n_0_54));
   DLH_X1 i_0_119 (.D(n_0_1), .G(n_0_88), .Q(n_0_55));
   DFF_X1 \in_data_reg[31]  (.D(dcm_out_data[31]), .CK(n_0_0), .Q(in_data[31]), 
      .QN());
   DFF_X1 \in_data_reg[30]  (.D(dcm_out_data[30]), .CK(n_0_0), .Q(in_data[30]), 
      .QN());
   DFF_X1 \in_data_reg[29]  (.D(dcm_out_data[29]), .CK(n_0_0), .Q(in_data[29]), 
      .QN());
   DFF_X1 \in_data_reg[28]  (.D(dcm_out_data[28]), .CK(n_0_0), .Q(in_data[28]), 
      .QN());
   DFF_X1 \in_data_reg[27]  (.D(dcm_out_data[27]), .CK(n_0_0), .Q(in_data[27]), 
      .QN());
   DFF_X1 \in_data_reg[26]  (.D(dcm_out_data[26]), .CK(n_0_0), .Q(in_data[26]), 
      .QN());
   DFF_X1 \in_data_reg[25]  (.D(dcm_out_data[25]), .CK(n_0_0), .Q(in_data[25]), 
      .QN());
   DFF_X1 \in_data_reg[24]  (.D(dcm_out_data[24]), .CK(n_0_0), .Q(in_data[24]), 
      .QN());
   DFF_X1 \in_data_reg[23]  (.D(dcm_out_data[23]), .CK(n_0_0), .Q(in_data[23]), 
      .QN());
   DFF_X1 \in_data_reg[22]  (.D(dcm_out_data[22]), .CK(n_0_0), .Q(in_data[22]), 
      .QN());
   DFF_X1 \in_data_reg[21]  (.D(dcm_out_data[21]), .CK(n_0_0), .Q(in_data[21]), 
      .QN());
   DFF_X1 \in_data_reg[20]  (.D(dcm_out_data[20]), .CK(n_0_0), .Q(in_data[20]), 
      .QN());
   DFF_X1 \in_data_reg[19]  (.D(dcm_out_data[19]), .CK(n_0_0), .Q(in_data[19]), 
      .QN());
   DFF_X1 \in_data_reg[18]  (.D(dcm_out_data[18]), .CK(n_0_0), .Q(in_data[18]), 
      .QN());
   DFF_X1 \in_data_reg[17]  (.D(dcm_out_data[17]), .CK(n_0_0), .Q(in_data[17]), 
      .QN());
   DFF_X1 \in_data_reg[16]  (.D(dcm_out_data[16]), .CK(n_0_0), .Q(in_data[16]), 
      .QN());
   DFF_X1 \in_data_reg[15]  (.D(dcm_out_data[15]), .CK(n_0_0), .Q(in_data[15]), 
      .QN());
   DFF_X1 \in_data_reg[14]  (.D(dcm_out_data[14]), .CK(n_0_0), .Q(in_data[14]), 
      .QN());
   DFF_X1 \in_data_reg[13]  (.D(dcm_out_data[13]), .CK(n_0_0), .Q(in_data[13]), 
      .QN());
   DFF_X1 \in_data_reg[12]  (.D(dcm_out_data[12]), .CK(n_0_0), .Q(in_data[12]), 
      .QN());
   DFF_X1 \in_data_reg[11]  (.D(dcm_out_data[11]), .CK(n_0_0), .Q(in_data[11]), 
      .QN());
   DFF_X1 \in_data_reg[10]  (.D(dcm_out_data[10]), .CK(n_0_0), .Q(in_data[10]), 
      .QN());
   DFF_X1 \in_data_reg[9]  (.D(dcm_out_data[9]), .CK(n_0_0), .Q(in_data[9]), 
      .QN());
   DFF_X1 \in_data_reg[8]  (.D(dcm_out_data[8]), .CK(n_0_0), .Q(in_data[8]), 
      .QN());
   DFF_X1 \in_data_reg[7]  (.D(dcm_out_data[7]), .CK(n_0_0), .Q(in_data[7]), 
      .QN());
   DFF_X1 \in_data_reg[6]  (.D(dcm_out_data[6]), .CK(n_0_0), .Q(in_data[6]), 
      .QN());
   DFF_X1 \in_data_reg[5]  (.D(dcm_out_data[5]), .CK(n_0_0), .Q(in_data[5]), 
      .QN());
   DFF_X1 \in_data_reg[4]  (.D(dcm_out_data[4]), .CK(n_0_0), .Q(in_data[4]), 
      .QN());
   DFF_X1 \in_data_reg[3]  (.D(dcm_out_data[3]), .CK(n_0_0), .Q(in_data[3]), 
      .QN());
   DFF_X1 \in_data_reg[2]  (.D(dcm_out_data[2]), .CK(n_0_0), .Q(in_data[2]), 
      .QN());
   DFF_X1 \in_data_reg[1]  (.D(dcm_out_data[1]), .CK(n_0_0), .Q(in_data[1]), 
      .QN());
   DFF_X1 \in_data_reg[0]  (.D(dcm_out_data[0]), .CK(n_0_0), .Q(in_data[0]), 
      .QN());
   MUX2_X1 i_0_0_0 (.A(to_std_logic), .B(n_0), .S(n_0_0_0), .Z(n_0_0_0));
   MUX2_X1 i_0_0_1 (.A(to_std_logic), .B(n_0), .S(n_0_0_1), .Z(n_0_0_1));
   MUX2_X1 i_0_0_2 (.A(to_std_logic), .B(n_0), .S(n_0_0_2), .Z(n_0_0_2));
   MUX2_X1 i_0_0_3 (.A(to_std_logic), .B(n_0), .S(n_0_0_3), .Z(n_0_0_3));
   MUX2_X1 i_0_0_4 (.A(to_std_logic), .B(n_0), .S(n_0_0_4), .Z(n_0_0_4));
   MUX2_X1 i_0_0_5 (.A(to_std_logic), .B(n_0), .S(n_0_0_5), .Z(n_0_0_5));
   MUX2_X1 i_0_0_58 (.A(n_0_0_10), .B(n_0_0_9), .S(n_0_0_6), .Z(n_0_0_6));
   MUX2_X1 i_0_0_59 (.A(n_0_0_10), .B(n_0_0_9), .S(n_0_0_7), .Z(n_0_0_7));
   NOR3_X1 i_0_0_10 (.A1(in_state[1]), .A2(n_0_0_8), .A3(n_0_0_14), .ZN(
      interrupt));
   NOR2_X1 i_0_0_11 (.A1(n_0_0_16), .A2(nau_done), .ZN(n_0_0_8));
   INV_X1 i_0_0_54 (.A(clk), .ZN(n_0_0));
   BUF_X1 rt_shieldBuf__4 (.A(in_state[1]), .Z(n_0_0_11));
   BUF_X1 rt_shieldBuf__4__4__0 (.A(n_0_0_10), .Z(to_std_logic));
   BUF_X1 rt_shieldBuf__4__4__1 (.A(n_0_0_9), .Z(n_0));
   INV_X1 i_0_0_8 (.A(dcm_error_success), .ZN(n_0_0_16));
   INV_X1 i_0_0_6 (.A(in_state[0]), .ZN(n_0_0_12));
   NOR2_X1 i_0_0_61 (.A1(n_0_0_12), .A2(in_state[1]), .ZN(n_0_0_9));
   NOR2_X1 i_0_0_13 (.A1(in_state[0]), .A2(in_state[1]), .ZN(n_0_0_10));
   INV_X1 i_0_0_14 (.A(rst), .ZN(n_0_0_13));
   NOR2_X1 i_0_0_15 (.A1(n_0_0_11), .A2(n_0_0_13), .ZN(n_0_21));
   AND2_X1 i_0_0_16 (.A1(n_0_0_0), .A2(rst), .ZN(n_0_1));
   NAND2_X1 i_0_0_17 (.A1(n_0_0_1), .A2(rst), .ZN(n_0_0_15));
   NOR2_X1 i_0_0_18 (.A1(n_0_0_2), .A2(n_0_0_13), .ZN(n_0_0_17));
   OAI211_X1 i_0_0_19 (.A(n_0_0_11), .B(n_0_0_15), .C1(n_0_0_17), .C2(
      in_state[0]), .ZN(n_0_88));
   AND2_X1 i_0_0_20 (.A1(n_0_0_3), .A2(in_data[0]), .ZN(n_0_56));
   AND2_X1 i_0_0_21 (.A1(n_0_0_3), .A2(in_data[1]), .ZN(n_0_57));
   AND2_X1 i_0_0_22 (.A1(n_0_0_3), .A2(in_data[2]), .ZN(n_0_58));
   AND2_X1 i_0_0_23 (.A1(n_0_0_3), .A2(in_data[3]), .ZN(n_0_59));
   AND2_X1 i_0_0_24 (.A1(n_0_0_3), .A2(in_data[4]), .ZN(n_0_60));
   AND2_X1 i_0_0_25 (.A1(n_0_0_3), .A2(in_data[5]), .ZN(n_0_61));
   AND2_X1 i_0_0_26 (.A1(n_0_0_3), .A2(in_data[6]), .ZN(n_0_62));
   AND2_X1 i_0_0_27 (.A1(n_0_0_3), .A2(in_data[7]), .ZN(n_0_63));
   AND2_X1 i_0_0_28 (.A1(n_0_0_3), .A2(in_data[8]), .ZN(n_0_64));
   AND2_X1 i_0_0_29 (.A1(n_0_0_3), .A2(in_data[9]), .ZN(n_0_65));
   AND2_X1 i_0_0_30 (.A1(n_0_0_3), .A2(in_data[10]), .ZN(n_0_66));
   AND2_X1 i_0_0_31 (.A1(n_0_0_3), .A2(in_data[11]), .ZN(n_0_67));
   AND2_X1 i_0_0_32 (.A1(n_0_0_3), .A2(in_data[12]), .ZN(n_0_68));
   AND2_X1 i_0_0_33 (.A1(n_0_0_3), .A2(in_data[13]), .ZN(n_0_69));
   AND2_X1 i_0_0_34 (.A1(n_0_0_3), .A2(in_data[14]), .ZN(n_0_70));
   AND2_X1 i_0_0_35 (.A1(n_0_0_3), .A2(in_data[15]), .ZN(n_0_71));
   AND2_X1 i_0_0_36 (.A1(n_0_0_3), .A2(in_data[16]), .ZN(n_0_72));
   AND2_X1 i_0_0_37 (.A1(n_0_0_3), .A2(in_data[17]), .ZN(n_0_73));
   AND2_X1 i_0_0_38 (.A1(n_0_0_3), .A2(in_data[18]), .ZN(n_0_74));
   AND2_X1 i_0_0_39 (.A1(n_0_0_3), .A2(in_data[19]), .ZN(n_0_75));
   AND2_X1 i_0_0_40 (.A1(n_0_0_3), .A2(in_data[20]), .ZN(n_0_76));
   AND2_X1 i_0_0_41 (.A1(n_0_0_3), .A2(in_data[21]), .ZN(n_0_77));
   AND2_X1 i_0_0_42 (.A1(n_0_0_3), .A2(in_data[22]), .ZN(n_0_78));
   AND2_X1 i_0_0_43 (.A1(n_0_0_3), .A2(in_data[23]), .ZN(n_0_79));
   AND2_X1 i_0_0_44 (.A1(n_0_0_3), .A2(in_data[24]), .ZN(n_0_80));
   AND2_X1 i_0_0_45 (.A1(n_0_0_3), .A2(in_data[25]), .ZN(n_0_81));
   AND2_X1 i_0_0_46 (.A1(n_0_0_3), .A2(in_data[26]), .ZN(n_0_82));
   AND2_X1 i_0_0_47 (.A1(n_0_0_3), .A2(in_data[27]), .ZN(n_0_83));
   AND2_X1 i_0_0_48 (.A1(n_0_0_3), .A2(in_data[28]), .ZN(n_0_84));
   AND2_X1 i_0_0_49 (.A1(n_0_0_3), .A2(in_data[29]), .ZN(n_0_85));
   AND2_X1 i_0_0_50 (.A1(n_0_0_3), .A2(in_data[30]), .ZN(n_0_86));
   AND2_X1 i_0_0_51 (.A1(n_0_0_3), .A2(in_data[31]), .ZN(n_0_87));
   INV_X1 i_0_0_7 (.A(n_0_0_11), .ZN(n_0_0_18));
   NOR4_X1 i_0_0_53 (.A1(n_0_0_4), .A2(n_0_0_5), .A3(n_0_0_13), .A4(n_0_0_18), 
      .ZN(n_0_0_19));
   AOI21_X1 i_0_0_55 (.A(n_0_0_19), .B1(n_0_0_18), .B2(n_0_0_13), .ZN(n_0_20));
   BUF_X1 i_0_0_60 (.A(n_0_0_13), .Z(n_0_0_14));
   INV_X1 i_0_0_9 (.A(n_0_0_6), .ZN(n_0_0_20));
   NAND2_X1 i_0_0_12 (.A1(n_0_0_18), .A2(dcm_error_success), .ZN(n_0_0_21));
   INV_X1 i_0_0_52 (.A(rst), .ZN(n_0_0_22));
   AOI21_X1 i_0_0_56 (.A(n_0_0_22), .B1(n_0_0_7), .B2(in_state[1]), .ZN(n_0_0_23));
   NAND3_X1 i_0_0_57 (.A1(n_0_0_20), .A2(n_0_0_21), .A3(n_0_0_23), .ZN(
      error_success));
endmodule
