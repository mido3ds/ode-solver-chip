/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sat Apr 25 22:05:33 2020
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 1371104287 */

module datapath(in_b, p_0);
   input [22:0]in_b;
   output [22:0]p_0;

   XOR2_X1 i_0 (.A(in_b[1]), .B(in_b[0]), .Z(p_0[1]));
   AND2_X1 i_1 (.A1(n_20), .A2(n_0), .ZN(p_0[2]));
   OAI21_X1 i_2 (.A(in_b[2]), .B1(in_b[1]), .B2(in_b[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(in_b[3]), .B(n_20), .Z(p_0[3]));
   XOR2_X1 i_4 (.A(in_b[4]), .B(n_19), .Z(p_0[4]));
   XOR2_X1 i_5 (.A(in_b[5]), .B(n_18), .Z(p_0[5]));
   AND2_X1 i_6 (.A1(n_17), .A2(n_1), .ZN(p_0[6]));
   OAI21_X1 i_7 (.A(in_b[6]), .B1(n_18), .B2(in_b[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(in_b[7]), .B(n_17), .Z(p_0[7]));
   XOR2_X1 i_9 (.A(in_b[8]), .B(n_16), .Z(p_0[8]));
   AND2_X1 i_10 (.A1(n_15), .A2(n_2), .ZN(p_0[9]));
   OAI21_X1 i_11 (.A(in_b[9]), .B1(n_16), .B2(in_b[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(in_b[10]), .B(n_15), .Z(p_0[10]));
   XNOR2_X1 i_13 (.A(in_b[11]), .B(n_14), .ZN(p_0[11]));
   XOR2_X1 i_14 (.A(in_b[12]), .B(n_13), .Z(p_0[12]));
   XOR2_X1 i_15 (.A(in_b[13]), .B(n_12), .Z(p_0[13]));
   XNOR2_X1 i_16 (.A(in_b[14]), .B(n_11), .ZN(p_0[14]));
   XNOR2_X1 i_17 (.A(in_b[15]), .B(n_10), .ZN(p_0[15]));
   XOR2_X1 i_18 (.A(in_b[16]), .B(n_9), .Z(p_0[16]));
   XOR2_X1 i_19 (.A(in_b[17]), .B(n_8), .Z(p_0[17]));
   XNOR2_X1 i_20 (.A(in_b[18]), .B(n_7), .ZN(p_0[18]));
   XNOR2_X1 i_21 (.A(in_b[19]), .B(n_6), .ZN(p_0[19]));
   XOR2_X1 i_22 (.A(in_b[20]), .B(n_5), .Z(p_0[20]));
   XNOR2_X1 i_23 (.A(in_b[21]), .B(n_4), .ZN(p_0[21]));
   XNOR2_X1 i_24 (.A(in_b[22]), .B(n_3), .ZN(p_0[22]));
   NOR3_X1 i_25 (.A1(n_5), .A2(in_b[20]), .A3(in_b[21]), .ZN(n_3));
   NOR2_X1 i_26 (.A1(n_5), .A2(in_b[20]), .ZN(n_4));
   NAND2_X1 i_27 (.A1(n_6), .A2(n_23), .ZN(n_5));
   NOR3_X1 i_28 (.A1(n_8), .A2(in_b[17]), .A3(in_b[18]), .ZN(n_6));
   NOR2_X1 i_29 (.A1(n_8), .A2(in_b[17]), .ZN(n_7));
   OR2_X1 i_30 (.A1(n_9), .A2(in_b[16]), .ZN(n_8));
   NAND2_X1 i_31 (.A1(n_10), .A2(n_22), .ZN(n_9));
   NOR3_X1 i_32 (.A1(n_12), .A2(in_b[13]), .A3(in_b[14]), .ZN(n_10));
   NOR2_X1 i_33 (.A1(n_12), .A2(in_b[13]), .ZN(n_11));
   OR2_X1 i_34 (.A1(n_13), .A2(in_b[12]), .ZN(n_12));
   NAND2_X1 i_35 (.A1(n_14), .A2(n_21), .ZN(n_13));
   NOR2_X1 i_36 (.A1(n_15), .A2(in_b[10]), .ZN(n_14));
   OR3_X1 i_37 (.A1(n_16), .A2(in_b[8]), .A3(in_b[9]), .ZN(n_15));
   OR2_X1 i_38 (.A1(n_17), .A2(in_b[7]), .ZN(n_16));
   OR3_X1 i_39 (.A1(n_18), .A2(in_b[5]), .A3(in_b[6]), .ZN(n_17));
   OR2_X1 i_40 (.A1(n_19), .A2(in_b[4]), .ZN(n_18));
   OR2_X1 i_41 (.A1(n_20), .A2(in_b[3]), .ZN(n_19));
   OR3_X1 i_42 (.A1(in_b[2]), .A2(in_b[1]), .A3(in_b[0]), .ZN(n_20));
   INV_X1 i_43 (.A(in_b[11]), .ZN(n_21));
   INV_X1 i_44 (.A(in_b[15]), .ZN(n_22));
   INV_X1 i_45 (.A(in_b[19]), .ZN(n_23));
endmodule

module datapath__0_7(p_0, p_1);
   input [22:0]p_0;
   output [22:0]p_1;

   XOR2_X1 i_0 (.A(p_0[1]), .B(p_0[0]), .Z(p_1[1]));
   AND2_X1 i_1 (.A1(n_19), .A2(n_0), .ZN(p_1[2]));
   OAI21_X1 i_2 (.A(p_0[2]), .B1(p_0[1]), .B2(p_0[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(p_0[3]), .B(n_19), .Z(p_1[3]));
   XOR2_X1 i_4 (.A(p_0[4]), .B(n_18), .Z(p_1[4]));
   XOR2_X1 i_5 (.A(p_0[5]), .B(n_17), .Z(p_1[5]));
   AND2_X1 i_6 (.A1(n_16), .A2(n_1), .ZN(p_1[6]));
   OAI21_X1 i_7 (.A(p_0[6]), .B1(n_17), .B2(p_0[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(p_0[7]), .B(n_16), .Z(p_1[7]));
   XOR2_X1 i_9 (.A(p_0[8]), .B(n_15), .Z(p_1[8]));
   AND2_X1 i_10 (.A1(n_14), .A2(n_2), .ZN(p_1[9]));
   OAI21_X1 i_11 (.A(p_0[9]), .B1(n_15), .B2(p_0[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(p_0[10]), .B(n_14), .Z(p_1[10]));
   XNOR2_X1 i_13 (.A(p_0[11]), .B(n_13), .ZN(p_1[11]));
   XOR2_X1 i_14 (.A(p_0[12]), .B(n_12), .Z(p_1[12]));
   XOR2_X1 i_15 (.A(p_0[13]), .B(n_11), .Z(p_1[13]));
   XNOR2_X1 i_16 (.A(p_0[14]), .B(n_10), .ZN(p_1[14]));
   XNOR2_X1 i_17 (.A(p_0[15]), .B(n_9), .ZN(p_1[15]));
   XOR2_X1 i_18 (.A(p_0[16]), .B(n_8), .Z(p_1[16]));
   XOR2_X1 i_19 (.A(p_0[17]), .B(n_7), .Z(p_1[17]));
   XNOR2_X1 i_20 (.A(p_0[18]), .B(n_6), .ZN(p_1[18]));
   XNOR2_X1 i_21 (.A(p_0[19]), .B(n_5), .ZN(p_1[19]));
   XOR2_X1 i_22 (.A(p_0[20]), .B(n_4), .Z(p_1[20]));
   XNOR2_X1 i_23 (.A(p_0[21]), .B(n_3), .ZN(p_1[21]));
   NOR2_X1 i_24 (.A1(n_4), .A2(p_0[20]), .ZN(n_3));
   NAND2_X1 i_25 (.A1(n_5), .A2(n_22), .ZN(n_4));
   NOR3_X1 i_26 (.A1(n_7), .A2(p_0[17]), .A3(p_0[18]), .ZN(n_5));
   NOR2_X1 i_27 (.A1(n_7), .A2(p_0[17]), .ZN(n_6));
   OR2_X1 i_28 (.A1(n_8), .A2(p_0[16]), .ZN(n_7));
   NAND2_X1 i_29 (.A1(n_9), .A2(n_21), .ZN(n_8));
   NOR3_X1 i_30 (.A1(n_11), .A2(p_0[13]), .A3(p_0[14]), .ZN(n_9));
   NOR2_X1 i_31 (.A1(n_11), .A2(p_0[13]), .ZN(n_10));
   OR2_X1 i_32 (.A1(n_12), .A2(p_0[12]), .ZN(n_11));
   NAND2_X1 i_33 (.A1(n_13), .A2(n_20), .ZN(n_12));
   NOR2_X1 i_34 (.A1(n_14), .A2(p_0[10]), .ZN(n_13));
   OR3_X1 i_35 (.A1(n_15), .A2(p_0[8]), .A3(p_0[9]), .ZN(n_14));
   OR2_X1 i_36 (.A1(n_16), .A2(p_0[7]), .ZN(n_15));
   OR3_X1 i_37 (.A1(n_17), .A2(p_0[5]), .A3(p_0[6]), .ZN(n_16));
   OR2_X1 i_38 (.A1(n_18), .A2(p_0[4]), .ZN(n_17));
   OR2_X1 i_39 (.A1(n_19), .A2(p_0[3]), .ZN(n_18));
   OR3_X1 i_40 (.A1(p_0[2]), .A2(p_0[1]), .A3(p_0[0]), .ZN(n_19));
   INV_X1 i_41 (.A(p_0[11]), .ZN(n_20));
   INV_X1 i_42 (.A(p_0[15]), .ZN(n_21));
   INV_X1 i_43 (.A(p_0[19]), .ZN(n_22));
endmodule

module datapath__0_9(p_0, p_1, divider);
   input [22:0]p_0;
   input [22:0]p_1;
   output [22:0]divider;

   HA_X1 i_0 (.A(p_0[0]), .B(p_1[0]), .CO(n_0), .S(divider[0]));
   HA_X1 i_1 (.A(p_0[1]), .B(n_0), .CO(n_1), .S(divider[1]));
   HA_X1 i_2 (.A(p_0[2]), .B(n_1), .CO(n_2), .S(divider[2]));
   HA_X1 i_3 (.A(p_0[3]), .B(n_2), .CO(n_3), .S(divider[3]));
   HA_X1 i_4 (.A(p_0[4]), .B(n_3), .CO(n_4), .S(divider[4]));
   HA_X1 i_5 (.A(p_0[5]), .B(n_4), .CO(n_5), .S(divider[5]));
   HA_X1 i_6 (.A(p_0[6]), .B(n_5), .CO(n_6), .S(divider[6]));
   HA_X1 i_7 (.A(p_0[7]), .B(n_6), .CO(n_7), .S(divider[7]));
   HA_X1 i_8 (.A(p_0[8]), .B(n_7), .CO(n_8), .S(divider[8]));
   HA_X1 i_9 (.A(p_0[9]), .B(n_8), .CO(n_9), .S(divider[9]));
   HA_X1 i_10 (.A(p_0[10]), .B(n_9), .CO(n_10), .S(divider[10]));
   HA_X1 i_11 (.A(p_0[11]), .B(n_10), .CO(n_11), .S(divider[11]));
   HA_X1 i_12 (.A(p_0[12]), .B(n_11), .CO(n_12), .S(divider[12]));
   HA_X1 i_13 (.A(p_0[13]), .B(n_12), .CO(n_13), .S(divider[13]));
   HA_X1 i_14 (.A(p_0[14]), .B(n_13), .CO(n_14), .S(divider[14]));
   HA_X1 i_15 (.A(p_0[15]), .B(n_14), .CO(n_15), .S(divider[15]));
   HA_X1 i_16 (.A(p_0[16]), .B(n_15), .CO(n_16), .S(divider[16]));
   HA_X1 i_17 (.A(p_0[17]), .B(n_16), .CO(n_17), .S(divider[17]));
   HA_X1 i_18 (.A(p_0[18]), .B(n_17), .CO(n_18), .S(divider[18]));
   HA_X1 i_19 (.A(p_0[19]), .B(n_18), .CO(n_19), .S(divider[19]));
   HA_X1 i_20 (.A(p_0[20]), .B(n_19), .CO(n_20), .S(divider[20]));
   HA_X1 i_21 (.A(p_0[21]), .B(n_20), .CO(n_21), .S(divider[21]));
endmodule

module datapath__0_13(p_0, p_1, divider);
   input [22:0]p_0;
   input [22:0]p_1;
   output [22:0]divider;

   HA_X1 i_0 (.A(p_0[0]), .B(p_1[0]), .CO(n_0), .S(divider[0]));
   FA_X1 i_1 (.A(p_0[1]), .B(p_1[1]), .CI(n_0), .CO(n_1), .S(divider[1]));
   FA_X1 i_2 (.A(p_0[2]), .B(p_1[2]), .CI(n_1), .CO(n_2), .S(divider[2]));
   FA_X1 i_3 (.A(p_0[3]), .B(p_1[3]), .CI(n_2), .CO(n_3), .S(divider[3]));
   FA_X1 i_4 (.A(p_0[4]), .B(p_1[4]), .CI(n_3), .CO(n_4), .S(divider[4]));
   FA_X1 i_5 (.A(p_0[5]), .B(p_1[5]), .CI(n_4), .CO(n_5), .S(divider[5]));
   FA_X1 i_6 (.A(p_0[6]), .B(p_1[6]), .CI(n_5), .CO(n_6), .S(divider[6]));
   FA_X1 i_7 (.A(p_0[7]), .B(p_1[7]), .CI(n_6), .CO(n_7), .S(divider[7]));
   FA_X1 i_8 (.A(p_0[8]), .B(p_1[8]), .CI(n_7), .CO(n_8), .S(divider[8]));
   FA_X1 i_9 (.A(p_0[9]), .B(p_1[9]), .CI(n_8), .CO(n_9), .S(divider[9]));
   FA_X1 i_10 (.A(p_0[10]), .B(p_1[10]), .CI(n_9), .CO(n_10), .S(divider[10]));
   FA_X1 i_11 (.A(p_0[11]), .B(p_1[11]), .CI(n_10), .CO(n_11), .S(divider[11]));
   FA_X1 i_12 (.A(p_0[12]), .B(p_1[12]), .CI(n_11), .CO(n_12), .S(divider[12]));
   FA_X1 i_13 (.A(p_0[13]), .B(p_1[13]), .CI(n_12), .CO(n_13), .S(divider[13]));
   FA_X1 i_14 (.A(p_0[14]), .B(p_1[14]), .CI(n_13), .CO(n_14), .S(divider[14]));
   FA_X1 i_15 (.A(p_0[15]), .B(p_1[15]), .CI(n_14), .CO(n_15), .S(divider[15]));
   FA_X1 i_16 (.A(p_0[16]), .B(p_1[16]), .CI(n_15), .CO(n_16), .S(divider[16]));
   FA_X1 i_17 (.A(p_0[17]), .B(p_1[17]), .CI(n_16), .CO(n_17), .S(divider[17]));
   FA_X1 i_18 (.A(p_0[18]), .B(p_1[18]), .CI(n_17), .CO(n_18), .S(divider[18]));
   FA_X1 i_19 (.A(p_0[19]), .B(p_1[19]), .CI(n_18), .CO(n_19), .S(divider[19]));
   FA_X1 i_20 (.A(p_0[20]), .B(p_1[20]), .CI(n_19), .CO(n_20), .S(divider[20]));
   FA_X1 i_21 (.A(p_0[21]), .B(p_1[21]), .CI(n_20), .CO(n_21), .S(divider[21]));
endmodule

module datapath__0_17(p_0, p_1, divider);
   input [22:0]p_0;
   input [22:0]p_1;
   output [22:0]divider;

   HA_X1 i_0 (.A(p_0[0]), .B(p_1[0]), .CO(n_0), .S(divider[0]));
   FA_X1 i_1 (.A(p_0[1]), .B(p_1[1]), .CI(n_0), .CO(n_1), .S(divider[1]));
   FA_X1 i_2 (.A(p_0[2]), .B(p_1[2]), .CI(n_1), .CO(n_2), .S(divider[2]));
   FA_X1 i_3 (.A(p_0[3]), .B(p_1[3]), .CI(n_2), .CO(n_3), .S(divider[3]));
   FA_X1 i_4 (.A(p_0[4]), .B(p_1[4]), .CI(n_3), .CO(n_4), .S(divider[4]));
   FA_X1 i_5 (.A(p_0[5]), .B(p_1[5]), .CI(n_4), .CO(n_5), .S(divider[5]));
   FA_X1 i_6 (.A(p_0[6]), .B(p_1[6]), .CI(n_5), .CO(n_6), .S(divider[6]));
   FA_X1 i_7 (.A(p_0[7]), .B(p_1[7]), .CI(n_6), .CO(n_7), .S(divider[7]));
   FA_X1 i_8 (.A(p_0[8]), .B(p_1[8]), .CI(n_7), .CO(n_8), .S(divider[8]));
   FA_X1 i_9 (.A(p_0[9]), .B(p_1[9]), .CI(n_8), .CO(n_9), .S(divider[9]));
   FA_X1 i_10 (.A(p_0[10]), .B(p_1[10]), .CI(n_9), .CO(n_10), .S(divider[10]));
   FA_X1 i_11 (.A(p_0[11]), .B(p_1[11]), .CI(n_10), .CO(n_11), .S(divider[11]));
   FA_X1 i_12 (.A(p_0[12]), .B(p_1[12]), .CI(n_11), .CO(n_12), .S(divider[12]));
   FA_X1 i_13 (.A(p_0[13]), .B(p_1[13]), .CI(n_12), .CO(n_13), .S(divider[13]));
   FA_X1 i_14 (.A(p_0[14]), .B(p_1[14]), .CI(n_13), .CO(n_14), .S(divider[14]));
   FA_X1 i_15 (.A(p_0[15]), .B(p_1[15]), .CI(n_14), .CO(n_15), .S(divider[15]));
   FA_X1 i_16 (.A(p_0[16]), .B(p_1[16]), .CI(n_15), .CO(n_16), .S(divider[16]));
   FA_X1 i_17 (.A(p_0[17]), .B(p_1[17]), .CI(n_16), .CO(n_17), .S(divider[17]));
   FA_X1 i_18 (.A(p_0[18]), .B(p_1[18]), .CI(n_17), .CO(n_18), .S(divider[18]));
   FA_X1 i_19 (.A(p_0[19]), .B(p_1[19]), .CI(n_18), .CO(n_19), .S(divider[19]));
   FA_X1 i_20 (.A(p_0[20]), .B(p_1[20]), .CI(n_19), .CO(n_20), .S(divider[20]));
   FA_X1 i_21 (.A(p_0[21]), .B(p_1[21]), .CI(n_20), .CO(n_21), .S(divider[21]));
endmodule

module datapath__0_21(p_0, p_1, divider);
   input [22:0]p_0;
   input [22:0]p_1;
   output [22:0]divider;

   HA_X1 i_0 (.A(p_0[0]), .B(p_1[0]), .CO(n_0), .S(divider[0]));
   FA_X1 i_1 (.A(p_0[1]), .B(p_1[1]), .CI(n_0), .CO(n_1), .S(divider[1]));
   FA_X1 i_2 (.A(p_0[2]), .B(p_1[2]), .CI(n_1), .CO(n_2), .S(divider[2]));
   FA_X1 i_3 (.A(p_0[3]), .B(p_1[3]), .CI(n_2), .CO(n_3), .S(divider[3]));
   FA_X1 i_4 (.A(p_0[4]), .B(p_1[4]), .CI(n_3), .CO(n_4), .S(divider[4]));
   FA_X1 i_5 (.A(p_0[5]), .B(p_1[5]), .CI(n_4), .CO(n_5), .S(divider[5]));
   FA_X1 i_6 (.A(p_0[6]), .B(p_1[6]), .CI(n_5), .CO(n_6), .S(divider[6]));
   FA_X1 i_7 (.A(p_0[7]), .B(p_1[7]), .CI(n_6), .CO(n_7), .S(divider[7]));
   FA_X1 i_8 (.A(p_0[8]), .B(p_1[8]), .CI(n_7), .CO(n_8), .S(divider[8]));
   FA_X1 i_9 (.A(p_0[9]), .B(p_1[9]), .CI(n_8), .CO(n_9), .S(divider[9]));
   FA_X1 i_10 (.A(p_0[10]), .B(p_1[10]), .CI(n_9), .CO(n_10), .S(divider[10]));
   FA_X1 i_11 (.A(p_0[11]), .B(p_1[11]), .CI(n_10), .CO(n_11), .S(divider[11]));
   FA_X1 i_12 (.A(p_0[12]), .B(p_1[12]), .CI(n_11), .CO(n_12), .S(divider[12]));
   FA_X1 i_13 (.A(p_0[13]), .B(p_1[13]), .CI(n_12), .CO(n_13), .S(divider[13]));
   FA_X1 i_14 (.A(p_0[14]), .B(p_1[14]), .CI(n_13), .CO(n_14), .S(divider[14]));
   FA_X1 i_15 (.A(p_0[15]), .B(p_1[15]), .CI(n_14), .CO(n_15), .S(divider[15]));
   FA_X1 i_16 (.A(p_0[16]), .B(p_1[16]), .CI(n_15), .CO(n_16), .S(divider[16]));
   FA_X1 i_17 (.A(p_0[17]), .B(p_1[17]), .CI(n_16), .CO(n_17), .S(divider[17]));
   FA_X1 i_18 (.A(p_0[18]), .B(p_1[18]), .CI(n_17), .CO(n_18), .S(divider[18]));
   FA_X1 i_19 (.A(p_0[19]), .B(p_1[19]), .CI(n_18), .CO(n_19), .S(divider[19]));
   FA_X1 i_20 (.A(p_0[20]), .B(p_1[20]), .CI(n_19), .CO(n_20), .S(divider[20]));
   FA_X1 i_21 (.A(p_0[21]), .B(p_1[21]), .CI(n_20), .CO(n_21), .S(divider[21]));
endmodule

module datapath__0_25(p_0, p_1, divider);
   input [22:0]p_0;
   input [22:0]p_1;
   output [22:0]divider;

   HA_X1 i_0 (.A(p_0[0]), .B(p_1[0]), .CO(n_0), .S(divider[0]));
   FA_X1 i_1 (.A(p_0[1]), .B(p_1[1]), .CI(n_0), .CO(n_1), .S(divider[1]));
   FA_X1 i_2 (.A(p_0[2]), .B(p_1[2]), .CI(n_1), .CO(n_2), .S(divider[2]));
   FA_X1 i_3 (.A(p_0[3]), .B(p_1[3]), .CI(n_2), .CO(n_3), .S(divider[3]));
   FA_X1 i_4 (.A(p_0[4]), .B(p_1[4]), .CI(n_3), .CO(n_4), .S(divider[4]));
   FA_X1 i_5 (.A(p_0[5]), .B(p_1[5]), .CI(n_4), .CO(n_5), .S(divider[5]));
   FA_X1 i_6 (.A(p_0[6]), .B(p_1[6]), .CI(n_5), .CO(n_6), .S(divider[6]));
   FA_X1 i_7 (.A(p_0[7]), .B(p_1[7]), .CI(n_6), .CO(n_7), .S(divider[7]));
   FA_X1 i_8 (.A(p_0[8]), .B(p_1[8]), .CI(n_7), .CO(n_8), .S(divider[8]));
   FA_X1 i_9 (.A(p_0[9]), .B(p_1[9]), .CI(n_8), .CO(n_9), .S(divider[9]));
   FA_X1 i_10 (.A(p_0[10]), .B(p_1[10]), .CI(n_9), .CO(n_10), .S(divider[10]));
   FA_X1 i_11 (.A(p_0[11]), .B(p_1[11]), .CI(n_10), .CO(n_11), .S(divider[11]));
   FA_X1 i_12 (.A(p_0[12]), .B(p_1[12]), .CI(n_11), .CO(n_12), .S(divider[12]));
   FA_X1 i_13 (.A(p_0[13]), .B(p_1[13]), .CI(n_12), .CO(n_13), .S(divider[13]));
   FA_X1 i_14 (.A(p_0[14]), .B(p_1[14]), .CI(n_13), .CO(n_14), .S(divider[14]));
   FA_X1 i_15 (.A(p_0[15]), .B(p_1[15]), .CI(n_14), .CO(n_15), .S(divider[15]));
   FA_X1 i_16 (.A(p_0[16]), .B(p_1[16]), .CI(n_15), .CO(n_16), .S(divider[16]));
   FA_X1 i_17 (.A(p_0[17]), .B(p_1[17]), .CI(n_16), .CO(n_17), .S(divider[17]));
   FA_X1 i_18 (.A(p_0[18]), .B(p_1[18]), .CI(n_17), .CO(n_18), .S(divider[18]));
   FA_X1 i_19 (.A(p_0[19]), .B(p_1[19]), .CI(n_18), .CO(n_19), .S(divider[19]));
   FA_X1 i_20 (.A(p_0[20]), .B(p_1[20]), .CI(n_19), .CO(n_20), .S(divider[20]));
   FA_X1 i_21 (.A(p_0[21]), .B(p_1[21]), .CI(n_20), .CO(n_21), .S(divider[21]));
endmodule

module datapath__0_29(p_0, p_1, divider);
   input [22:0]p_0;
   input [22:0]p_1;
   output [22:0]divider;

   HA_X1 i_0 (.A(p_0[0]), .B(p_1[0]), .CO(n_0), .S(divider[0]));
   FA_X1 i_1 (.A(p_0[1]), .B(p_1[1]), .CI(n_0), .CO(n_1), .S(divider[1]));
   FA_X1 i_2 (.A(p_0[2]), .B(p_1[2]), .CI(n_1), .CO(n_2), .S(divider[2]));
   FA_X1 i_3 (.A(p_0[3]), .B(p_1[3]), .CI(n_2), .CO(n_3), .S(divider[3]));
   FA_X1 i_4 (.A(p_0[4]), .B(p_1[4]), .CI(n_3), .CO(n_4), .S(divider[4]));
   FA_X1 i_5 (.A(p_0[5]), .B(p_1[5]), .CI(n_4), .CO(n_5), .S(divider[5]));
   FA_X1 i_6 (.A(p_0[6]), .B(p_1[6]), .CI(n_5), .CO(n_6), .S(divider[6]));
   FA_X1 i_7 (.A(p_0[7]), .B(p_1[7]), .CI(n_6), .CO(n_7), .S(divider[7]));
   FA_X1 i_8 (.A(p_0[8]), .B(p_1[8]), .CI(n_7), .CO(n_8), .S(divider[8]));
   FA_X1 i_9 (.A(p_0[9]), .B(p_1[9]), .CI(n_8), .CO(n_9), .S(divider[9]));
   FA_X1 i_10 (.A(p_0[10]), .B(p_1[10]), .CI(n_9), .CO(n_10), .S(divider[10]));
   FA_X1 i_11 (.A(p_0[11]), .B(p_1[11]), .CI(n_10), .CO(n_11), .S(divider[11]));
   FA_X1 i_12 (.A(p_0[12]), .B(p_1[12]), .CI(n_11), .CO(n_12), .S(divider[12]));
   FA_X1 i_13 (.A(p_0[13]), .B(p_1[13]), .CI(n_12), .CO(n_13), .S(divider[13]));
   FA_X1 i_14 (.A(p_0[14]), .B(p_1[14]), .CI(n_13), .CO(n_14), .S(divider[14]));
   FA_X1 i_15 (.A(p_0[15]), .B(p_1[15]), .CI(n_14), .CO(n_15), .S(divider[15]));
   FA_X1 i_16 (.A(p_0[16]), .B(p_1[16]), .CI(n_15), .CO(n_16), .S(divider[16]));
   FA_X1 i_17 (.A(p_0[17]), .B(p_1[17]), .CI(n_16), .CO(n_17), .S(divider[17]));
   FA_X1 i_18 (.A(p_0[18]), .B(p_1[18]), .CI(n_17), .CO(n_18), .S(divider[18]));
   FA_X1 i_19 (.A(p_0[19]), .B(p_1[19]), .CI(n_18), .CO(n_19), .S(divider[19]));
   FA_X1 i_20 (.A(p_0[20]), .B(p_1[20]), .CI(n_19), .CO(n_20), .S(divider[20]));
   FA_X1 i_21 (.A(p_0[21]), .B(p_1[21]), .CI(n_20), .CO(n_21), .S(divider[21]));
endmodule

module datapath__0_33(p_0, p_1, divider);
   input [22:0]p_0;
   input [22:0]p_1;
   output [22:0]divider;

   HA_X1 i_0 (.A(p_0[0]), .B(p_1[0]), .CO(n_0), .S(divider[0]));
   FA_X1 i_1 (.A(p_0[1]), .B(p_1[1]), .CI(n_0), .CO(n_1), .S(divider[1]));
   FA_X1 i_2 (.A(p_0[2]), .B(p_1[2]), .CI(n_1), .CO(n_2), .S(divider[2]));
   FA_X1 i_3 (.A(p_0[3]), .B(p_1[3]), .CI(n_2), .CO(n_3), .S(divider[3]));
   FA_X1 i_4 (.A(p_0[4]), .B(p_1[4]), .CI(n_3), .CO(n_4), .S(divider[4]));
   FA_X1 i_5 (.A(p_0[5]), .B(p_1[5]), .CI(n_4), .CO(n_5), .S(divider[5]));
   FA_X1 i_6 (.A(p_0[6]), .B(p_1[6]), .CI(n_5), .CO(n_6), .S(divider[6]));
   FA_X1 i_7 (.A(p_0[7]), .B(p_1[7]), .CI(n_6), .CO(n_7), .S(divider[7]));
   FA_X1 i_8 (.A(p_0[8]), .B(p_1[8]), .CI(n_7), .CO(n_8), .S(divider[8]));
   FA_X1 i_9 (.A(p_0[9]), .B(p_1[9]), .CI(n_8), .CO(n_9), .S(divider[9]));
   FA_X1 i_10 (.A(p_0[10]), .B(p_1[10]), .CI(n_9), .CO(n_10), .S(divider[10]));
   FA_X1 i_11 (.A(p_0[11]), .B(p_1[11]), .CI(n_10), .CO(n_11), .S(divider[11]));
   FA_X1 i_12 (.A(p_0[12]), .B(p_1[12]), .CI(n_11), .CO(n_12), .S(divider[12]));
   FA_X1 i_13 (.A(p_0[13]), .B(p_1[13]), .CI(n_12), .CO(n_13), .S(divider[13]));
   FA_X1 i_14 (.A(p_0[14]), .B(p_1[14]), .CI(n_13), .CO(n_14), .S(divider[14]));
   FA_X1 i_15 (.A(p_0[15]), .B(p_1[15]), .CI(n_14), .CO(n_15), .S(divider[15]));
   FA_X1 i_16 (.A(p_0[16]), .B(p_1[16]), .CI(n_15), .CO(n_16), .S(divider[16]));
   FA_X1 i_17 (.A(p_0[17]), .B(p_1[17]), .CI(n_16), .CO(n_17), .S(divider[17]));
   FA_X1 i_18 (.A(p_0[18]), .B(p_1[18]), .CI(n_17), .CO(n_18), .S(divider[18]));
   FA_X1 i_19 (.A(p_0[19]), .B(p_1[19]), .CI(n_18), .CO(n_19), .S(divider[19]));
   FA_X1 i_20 (.A(p_0[20]), .B(p_1[20]), .CI(n_19), .CO(n_20), .S(divider[20]));
   FA_X1 i_21 (.A(p_0[21]), .B(p_1[21]), .CI(n_20), .CO(n_21), .S(divider[21]));
endmodule

module datapath__0_37(p_0, p_1, divider);
   input [22:0]p_0;
   input [22:0]p_1;
   output [22:0]divider;

   HA_X1 i_0 (.A(p_0[0]), .B(p_1[0]), .CO(n_0), .S(divider[0]));
   FA_X1 i_1 (.A(p_0[1]), .B(p_1[1]), .CI(n_0), .CO(n_1), .S(divider[1]));
   FA_X1 i_2 (.A(p_0[2]), .B(p_1[2]), .CI(n_1), .CO(n_2), .S(divider[2]));
   FA_X1 i_3 (.A(p_0[3]), .B(p_1[3]), .CI(n_2), .CO(n_3), .S(divider[3]));
   FA_X1 i_4 (.A(p_0[4]), .B(p_1[4]), .CI(n_3), .CO(n_4), .S(divider[4]));
   FA_X1 i_5 (.A(p_0[5]), .B(p_1[5]), .CI(n_4), .CO(n_5), .S(divider[5]));
   FA_X1 i_6 (.A(p_0[6]), .B(p_1[6]), .CI(n_5), .CO(n_6), .S(divider[6]));
   FA_X1 i_7 (.A(p_0[7]), .B(p_1[7]), .CI(n_6), .CO(n_7), .S(divider[7]));
   FA_X1 i_8 (.A(p_0[8]), .B(p_1[8]), .CI(n_7), .CO(n_8), .S(divider[8]));
   FA_X1 i_9 (.A(p_0[9]), .B(p_1[9]), .CI(n_8), .CO(n_9), .S(divider[9]));
   FA_X1 i_10 (.A(p_0[10]), .B(p_1[10]), .CI(n_9), .CO(n_10), .S(divider[10]));
   FA_X1 i_11 (.A(p_0[11]), .B(p_1[11]), .CI(n_10), .CO(n_11), .S(divider[11]));
   FA_X1 i_12 (.A(p_0[12]), .B(p_1[12]), .CI(n_11), .CO(n_12), .S(divider[12]));
   FA_X1 i_13 (.A(p_0[13]), .B(p_1[13]), .CI(n_12), .CO(n_13), .S(divider[13]));
   FA_X1 i_14 (.A(p_0[14]), .B(p_1[14]), .CI(n_13), .CO(n_14), .S(divider[14]));
   FA_X1 i_15 (.A(p_0[15]), .B(p_1[15]), .CI(n_14), .CO(n_15), .S(divider[15]));
   FA_X1 i_16 (.A(p_0[16]), .B(p_1[16]), .CI(n_15), .CO(n_16), .S(divider[16]));
   FA_X1 i_17 (.A(p_0[17]), .B(p_1[17]), .CI(n_16), .CO(n_17), .S(divider[17]));
   FA_X1 i_18 (.A(p_0[18]), .B(p_1[18]), .CI(n_17), .CO(n_18), .S(divider[18]));
   FA_X1 i_19 (.A(p_0[19]), .B(p_1[19]), .CI(n_18), .CO(n_19), .S(divider[19]));
   FA_X1 i_20 (.A(p_0[20]), .B(p_1[20]), .CI(n_19), .CO(n_20), .S(divider[20]));
   FA_X1 i_21 (.A(p_0[21]), .B(p_1[21]), .CI(n_20), .CO(n_21), .S(divider[21]));
endmodule

module datapath__0_41(p_0, p_1, divider);
   input [22:0]p_0;
   input [22:0]p_1;
   output [22:0]divider;

   HA_X1 i_0 (.A(p_0[0]), .B(p_1[0]), .CO(n_0), .S(divider[0]));
   FA_X1 i_1 (.A(p_0[1]), .B(p_1[1]), .CI(n_0), .CO(n_1), .S(divider[1]));
   FA_X1 i_2 (.A(p_0[2]), .B(p_1[2]), .CI(n_1), .CO(n_2), .S(divider[2]));
   FA_X1 i_3 (.A(p_0[3]), .B(p_1[3]), .CI(n_2), .CO(n_3), .S(divider[3]));
   FA_X1 i_4 (.A(p_0[4]), .B(p_1[4]), .CI(n_3), .CO(n_4), .S(divider[4]));
   FA_X1 i_5 (.A(p_0[5]), .B(p_1[5]), .CI(n_4), .CO(n_5), .S(divider[5]));
   FA_X1 i_6 (.A(p_0[6]), .B(p_1[6]), .CI(n_5), .CO(n_6), .S(divider[6]));
   FA_X1 i_7 (.A(p_0[7]), .B(p_1[7]), .CI(n_6), .CO(n_7), .S(divider[7]));
   FA_X1 i_8 (.A(p_0[8]), .B(p_1[8]), .CI(n_7), .CO(n_8), .S(divider[8]));
   FA_X1 i_9 (.A(p_0[9]), .B(p_1[9]), .CI(n_8), .CO(n_9), .S(divider[9]));
   FA_X1 i_10 (.A(p_0[10]), .B(p_1[10]), .CI(n_9), .CO(n_10), .S(divider[10]));
   FA_X1 i_11 (.A(p_0[11]), .B(p_1[11]), .CI(n_10), .CO(n_11), .S(divider[11]));
   FA_X1 i_12 (.A(p_0[12]), .B(p_1[12]), .CI(n_11), .CO(n_12), .S(divider[12]));
   FA_X1 i_13 (.A(p_0[13]), .B(p_1[13]), .CI(n_12), .CO(n_13), .S(divider[13]));
   FA_X1 i_14 (.A(p_0[14]), .B(p_1[14]), .CI(n_13), .CO(n_14), .S(divider[14]));
   FA_X1 i_15 (.A(p_0[15]), .B(p_1[15]), .CI(n_14), .CO(n_15), .S(divider[15]));
   FA_X1 i_16 (.A(p_0[16]), .B(p_1[16]), .CI(n_15), .CO(n_16), .S(divider[16]));
   FA_X1 i_17 (.A(p_0[17]), .B(p_1[17]), .CI(n_16), .CO(n_17), .S(divider[17]));
   FA_X1 i_18 (.A(p_0[18]), .B(p_1[18]), .CI(n_17), .CO(n_18), .S(divider[18]));
   FA_X1 i_19 (.A(p_0[19]), .B(p_1[19]), .CI(n_18), .CO(n_19), .S(divider[19]));
   FA_X1 i_20 (.A(p_0[20]), .B(p_1[20]), .CI(n_19), .CO(n_20), .S(divider[20]));
   FA_X1 i_21 (.A(p_0[21]), .B(p_1[21]), .CI(n_20), .CO(n_21), .S(divider[21]));
endmodule

module datapath__0_45(p_0, p_1, divider);
   input [22:0]p_0;
   input [22:0]p_1;
   output [22:0]divider;

   HA_X1 i_0 (.A(p_0[0]), .B(p_1[0]), .CO(n_0), .S(divider[0]));
   FA_X1 i_1 (.A(p_0[1]), .B(p_1[1]), .CI(n_0), .CO(n_1), .S(divider[1]));
   FA_X1 i_2 (.A(p_0[2]), .B(p_1[2]), .CI(n_1), .CO(n_2), .S(divider[2]));
   FA_X1 i_3 (.A(p_0[3]), .B(p_1[3]), .CI(n_2), .CO(n_3), .S(divider[3]));
   FA_X1 i_4 (.A(p_0[4]), .B(p_1[4]), .CI(n_3), .CO(n_4), .S(divider[4]));
   FA_X1 i_5 (.A(p_0[5]), .B(p_1[5]), .CI(n_4), .CO(n_5), .S(divider[5]));
   FA_X1 i_6 (.A(p_0[6]), .B(p_1[6]), .CI(n_5), .CO(n_6), .S(divider[6]));
   FA_X1 i_7 (.A(p_0[7]), .B(p_1[7]), .CI(n_6), .CO(n_7), .S(divider[7]));
   FA_X1 i_8 (.A(p_0[8]), .B(p_1[8]), .CI(n_7), .CO(n_8), .S(divider[8]));
   FA_X1 i_9 (.A(p_0[9]), .B(p_1[9]), .CI(n_8), .CO(n_9), .S(divider[9]));
   FA_X1 i_10 (.A(p_0[10]), .B(p_1[10]), .CI(n_9), .CO(n_10), .S(divider[10]));
   FA_X1 i_11 (.A(p_0[11]), .B(p_1[11]), .CI(n_10), .CO(n_11), .S(divider[11]));
   FA_X1 i_12 (.A(p_0[12]), .B(p_1[12]), .CI(n_11), .CO(n_12), .S(divider[12]));
   FA_X1 i_13 (.A(p_0[13]), .B(p_1[13]), .CI(n_12), .CO(n_13), .S(divider[13]));
   FA_X1 i_14 (.A(p_0[14]), .B(p_1[14]), .CI(n_13), .CO(n_14), .S(divider[14]));
   FA_X1 i_15 (.A(p_0[15]), .B(p_1[15]), .CI(n_14), .CO(n_15), .S(divider[15]));
   FA_X1 i_16 (.A(p_0[16]), .B(p_1[16]), .CI(n_15), .CO(n_16), .S(divider[16]));
   FA_X1 i_17 (.A(p_0[17]), .B(p_1[17]), .CI(n_16), .CO(n_17), .S(divider[17]));
   FA_X1 i_18 (.A(p_0[18]), .B(p_1[18]), .CI(n_17), .CO(n_18), .S(divider[18]));
   FA_X1 i_19 (.A(p_0[19]), .B(p_1[19]), .CI(n_18), .CO(n_19), .S(divider[19]));
   FA_X1 i_20 (.A(p_0[20]), .B(p_1[20]), .CI(n_19), .CO(n_20), .S(divider[20]));
   FA_X1 i_21 (.A(p_0[21]), .B(p_1[21]), .CI(n_20), .CO(n_21), .S(divider[21]));
endmodule

module datapath__0_49(p_0, p_1, divider);
   input [22:0]p_0;
   input [22:0]p_1;
   output [22:0]divider;

   HA_X1 i_0 (.A(p_0[0]), .B(p_1[0]), .CO(n_0), .S(divider[0]));
   FA_X1 i_1 (.A(p_0[1]), .B(p_1[1]), .CI(n_0), .CO(n_1), .S(divider[1]));
   FA_X1 i_2 (.A(p_0[2]), .B(p_1[2]), .CI(n_1), .CO(n_2), .S(divider[2]));
   FA_X1 i_3 (.A(p_0[3]), .B(p_1[3]), .CI(n_2), .CO(n_3), .S(divider[3]));
   FA_X1 i_4 (.A(p_0[4]), .B(p_1[4]), .CI(n_3), .CO(n_4), .S(divider[4]));
   FA_X1 i_5 (.A(p_0[5]), .B(p_1[5]), .CI(n_4), .CO(n_5), .S(divider[5]));
   FA_X1 i_6 (.A(p_0[6]), .B(p_1[6]), .CI(n_5), .CO(n_6), .S(divider[6]));
   FA_X1 i_7 (.A(p_0[7]), .B(p_1[7]), .CI(n_6), .CO(n_7), .S(divider[7]));
   FA_X1 i_8 (.A(p_0[8]), .B(p_1[8]), .CI(n_7), .CO(n_8), .S(divider[8]));
   FA_X1 i_9 (.A(p_0[9]), .B(p_1[9]), .CI(n_8), .CO(n_9), .S(divider[9]));
   FA_X1 i_10 (.A(p_0[10]), .B(p_1[10]), .CI(n_9), .CO(n_10), .S(divider[10]));
   FA_X1 i_11 (.A(p_0[11]), .B(p_1[11]), .CI(n_10), .CO(n_11), .S(divider[11]));
   FA_X1 i_12 (.A(p_0[12]), .B(p_1[12]), .CI(n_11), .CO(n_12), .S(divider[12]));
   FA_X1 i_13 (.A(p_0[13]), .B(p_1[13]), .CI(n_12), .CO(n_13), .S(divider[13]));
   FA_X1 i_14 (.A(p_0[14]), .B(p_1[14]), .CI(n_13), .CO(n_14), .S(divider[14]));
   FA_X1 i_15 (.A(p_0[15]), .B(p_1[15]), .CI(n_14), .CO(n_15), .S(divider[15]));
   FA_X1 i_16 (.A(p_0[16]), .B(p_1[16]), .CI(n_15), .CO(n_16), .S(divider[16]));
   FA_X1 i_17 (.A(p_0[17]), .B(p_1[17]), .CI(n_16), .CO(n_17), .S(divider[17]));
   FA_X1 i_18 (.A(p_0[18]), .B(p_1[18]), .CI(n_17), .CO(n_18), .S(divider[18]));
   FA_X1 i_19 (.A(p_0[19]), .B(p_1[19]), .CI(n_18), .CO(n_19), .S(divider[19]));
   FA_X1 i_20 (.A(p_0[20]), .B(p_1[20]), .CI(n_19), .CO(n_20), .S(divider[20]));
   FA_X1 i_21 (.A(p_0[21]), .B(p_1[21]), .CI(n_20), .CO(n_21), .S(divider[21]));
endmodule

module datapath__0_53(p_0, p_1, divider);
   input [22:0]p_0;
   input [22:0]p_1;
   output [22:0]divider;

   HA_X1 i_0 (.A(p_0[0]), .B(p_1[0]), .CO(n_0), .S(divider[0]));
   FA_X1 i_1 (.A(p_0[1]), .B(p_1[1]), .CI(n_0), .CO(n_1), .S(divider[1]));
   FA_X1 i_2 (.A(p_0[2]), .B(p_1[2]), .CI(n_1), .CO(n_2), .S(divider[2]));
   FA_X1 i_3 (.A(p_0[3]), .B(p_1[3]), .CI(n_2), .CO(n_3), .S(divider[3]));
   FA_X1 i_4 (.A(p_0[4]), .B(p_1[4]), .CI(n_3), .CO(n_4), .S(divider[4]));
   FA_X1 i_5 (.A(p_0[5]), .B(p_1[5]), .CI(n_4), .CO(n_5), .S(divider[5]));
   FA_X1 i_6 (.A(p_0[6]), .B(p_1[6]), .CI(n_5), .CO(n_6), .S(divider[6]));
   FA_X1 i_7 (.A(p_0[7]), .B(p_1[7]), .CI(n_6), .CO(n_7), .S(divider[7]));
   FA_X1 i_8 (.A(p_0[8]), .B(p_1[8]), .CI(n_7), .CO(n_8), .S(divider[8]));
   FA_X1 i_9 (.A(p_0[9]), .B(p_1[9]), .CI(n_8), .CO(n_9), .S(divider[9]));
   FA_X1 i_10 (.A(p_0[10]), .B(p_1[10]), .CI(n_9), .CO(n_10), .S(divider[10]));
   FA_X1 i_11 (.A(p_0[11]), .B(p_1[11]), .CI(n_10), .CO(n_11), .S(divider[11]));
   FA_X1 i_12 (.A(p_0[12]), .B(p_1[12]), .CI(n_11), .CO(n_12), .S(divider[12]));
   FA_X1 i_13 (.A(p_0[13]), .B(p_1[13]), .CI(n_12), .CO(n_13), .S(divider[13]));
   FA_X1 i_14 (.A(p_0[14]), .B(p_1[14]), .CI(n_13), .CO(n_14), .S(divider[14]));
   FA_X1 i_15 (.A(p_0[15]), .B(p_1[15]), .CI(n_14), .CO(n_15), .S(divider[15]));
   FA_X1 i_16 (.A(p_0[16]), .B(p_1[16]), .CI(n_15), .CO(n_16), .S(divider[16]));
   FA_X1 i_17 (.A(p_0[17]), .B(p_1[17]), .CI(n_16), .CO(n_17), .S(divider[17]));
   FA_X1 i_18 (.A(p_0[18]), .B(p_1[18]), .CI(n_17), .CO(n_18), .S(divider[18]));
   FA_X1 i_19 (.A(p_0[19]), .B(p_1[19]), .CI(n_18), .CO(n_19), .S(divider[19]));
   FA_X1 i_20 (.A(p_0[20]), .B(p_1[20]), .CI(n_19), .CO(n_20), .S(divider[20]));
   FA_X1 i_21 (.A(p_0[21]), .B(p_1[21]), .CI(n_20), .CO(n_21), .S(divider[21]));
endmodule

module datapath__0_57(p_0, p_1, divider);
   input [22:0]p_0;
   input [22:0]p_1;
   output [22:0]divider;

   HA_X1 i_0 (.A(p_0[0]), .B(p_1[0]), .CO(n_0), .S(divider[0]));
   FA_X1 i_1 (.A(p_0[1]), .B(p_1[1]), .CI(n_0), .CO(n_1), .S(divider[1]));
   FA_X1 i_2 (.A(p_0[2]), .B(p_1[2]), .CI(n_1), .CO(n_2), .S(divider[2]));
   FA_X1 i_3 (.A(p_0[3]), .B(p_1[3]), .CI(n_2), .CO(n_3), .S(divider[3]));
   FA_X1 i_4 (.A(p_0[4]), .B(p_1[4]), .CI(n_3), .CO(n_4), .S(divider[4]));
   FA_X1 i_5 (.A(p_0[5]), .B(p_1[5]), .CI(n_4), .CO(n_5), .S(divider[5]));
   FA_X1 i_6 (.A(p_0[6]), .B(p_1[6]), .CI(n_5), .CO(n_6), .S(divider[6]));
   FA_X1 i_7 (.A(p_0[7]), .B(p_1[7]), .CI(n_6), .CO(n_7), .S(divider[7]));
   FA_X1 i_8 (.A(p_0[8]), .B(p_1[8]), .CI(n_7), .CO(n_8), .S(divider[8]));
   FA_X1 i_9 (.A(p_0[9]), .B(p_1[9]), .CI(n_8), .CO(n_9), .S(divider[9]));
   FA_X1 i_10 (.A(p_0[10]), .B(p_1[10]), .CI(n_9), .CO(n_10), .S(divider[10]));
   FA_X1 i_11 (.A(p_0[11]), .B(p_1[11]), .CI(n_10), .CO(n_11), .S(divider[11]));
   FA_X1 i_12 (.A(p_0[12]), .B(p_1[12]), .CI(n_11), .CO(n_12), .S(divider[12]));
   FA_X1 i_13 (.A(p_0[13]), .B(p_1[13]), .CI(n_12), .CO(n_13), .S(divider[13]));
   FA_X1 i_14 (.A(p_0[14]), .B(p_1[14]), .CI(n_13), .CO(n_14), .S(divider[14]));
   FA_X1 i_15 (.A(p_0[15]), .B(p_1[15]), .CI(n_14), .CO(n_15), .S(divider[15]));
   FA_X1 i_16 (.A(p_0[16]), .B(p_1[16]), .CI(n_15), .CO(n_16), .S(divider[16]));
   FA_X1 i_17 (.A(p_0[17]), .B(p_1[17]), .CI(n_16), .CO(n_17), .S(divider[17]));
   FA_X1 i_18 (.A(p_0[18]), .B(p_1[18]), .CI(n_17), .CO(n_18), .S(divider[18]));
   FA_X1 i_19 (.A(p_0[19]), .B(p_1[19]), .CI(n_18), .CO(n_19), .S(divider[19]));
   FA_X1 i_20 (.A(p_0[20]), .B(p_1[20]), .CI(n_19), .CO(n_20), .S(divider[20]));
   FA_X1 i_21 (.A(p_0[21]), .B(p_1[21]), .CI(n_20), .CO(n_21), .S(divider[21]));
endmodule

module datapath__0_61(p_0, p_1, divider);
   input [22:0]p_0;
   input [22:0]p_1;
   output [22:0]divider;

   HA_X1 i_0 (.A(p_0[0]), .B(p_1[0]), .CO(n_0), .S(divider[0]));
   FA_X1 i_1 (.A(p_0[1]), .B(p_1[1]), .CI(n_0), .CO(n_1), .S(divider[1]));
   FA_X1 i_2 (.A(p_0[2]), .B(p_1[2]), .CI(n_1), .CO(n_2), .S(divider[2]));
   FA_X1 i_3 (.A(p_0[3]), .B(p_1[3]), .CI(n_2), .CO(n_3), .S(divider[3]));
   FA_X1 i_4 (.A(p_0[4]), .B(p_1[4]), .CI(n_3), .CO(n_4), .S(divider[4]));
   FA_X1 i_5 (.A(p_0[5]), .B(p_1[5]), .CI(n_4), .CO(n_5), .S(divider[5]));
   FA_X1 i_6 (.A(p_0[6]), .B(p_1[6]), .CI(n_5), .CO(n_6), .S(divider[6]));
   FA_X1 i_7 (.A(p_0[7]), .B(p_1[7]), .CI(n_6), .CO(n_7), .S(divider[7]));
   FA_X1 i_8 (.A(p_0[8]), .B(p_1[8]), .CI(n_7), .CO(n_8), .S(divider[8]));
   FA_X1 i_9 (.A(p_0[9]), .B(p_1[9]), .CI(n_8), .CO(n_9), .S(divider[9]));
   FA_X1 i_10 (.A(p_0[10]), .B(p_1[10]), .CI(n_9), .CO(n_10), .S(divider[10]));
   FA_X1 i_11 (.A(p_0[11]), .B(p_1[11]), .CI(n_10), .CO(n_11), .S(divider[11]));
   FA_X1 i_12 (.A(p_0[12]), .B(p_1[12]), .CI(n_11), .CO(n_12), .S(divider[12]));
   FA_X1 i_13 (.A(p_0[13]), .B(p_1[13]), .CI(n_12), .CO(n_13), .S(divider[13]));
   FA_X1 i_14 (.A(p_0[14]), .B(p_1[14]), .CI(n_13), .CO(n_14), .S(divider[14]));
   FA_X1 i_15 (.A(p_0[15]), .B(p_1[15]), .CI(n_14), .CO(n_15), .S(divider[15]));
   FA_X1 i_16 (.A(p_0[16]), .B(p_1[16]), .CI(n_15), .CO(n_16), .S(divider[16]));
   FA_X1 i_17 (.A(p_0[17]), .B(p_1[17]), .CI(n_16), .CO(n_17), .S(divider[17]));
   FA_X1 i_18 (.A(p_0[18]), .B(p_1[18]), .CI(n_17), .CO(n_18), .S(divider[18]));
   FA_X1 i_19 (.A(p_0[19]), .B(p_1[19]), .CI(n_18), .CO(n_19), .S(divider[19]));
   FA_X1 i_20 (.A(p_0[20]), .B(p_1[20]), .CI(n_19), .CO(n_20), .S(divider[20]));
   FA_X1 i_21 (.A(p_0[21]), .B(p_1[21]), .CI(n_20), .CO(n_21), .S(divider[21]));
endmodule

module datapath__0_65(p_0, p_1, divider);
   input [22:0]p_0;
   input [22:0]p_1;
   output [22:0]divider;

   HA_X1 i_0 (.A(p_0[0]), .B(p_1[0]), .CO(n_0), .S(divider[0]));
   FA_X1 i_1 (.A(p_0[1]), .B(p_1[1]), .CI(n_0), .CO(n_1), .S(divider[1]));
   FA_X1 i_2 (.A(p_0[2]), .B(p_1[2]), .CI(n_1), .CO(n_2), .S(divider[2]));
   FA_X1 i_3 (.A(p_0[3]), .B(p_1[3]), .CI(n_2), .CO(n_3), .S(divider[3]));
   FA_X1 i_4 (.A(p_0[4]), .B(p_1[4]), .CI(n_3), .CO(n_4), .S(divider[4]));
   FA_X1 i_5 (.A(p_0[5]), .B(p_1[5]), .CI(n_4), .CO(n_5), .S(divider[5]));
   FA_X1 i_6 (.A(p_0[6]), .B(p_1[6]), .CI(n_5), .CO(n_6), .S(divider[6]));
   FA_X1 i_7 (.A(p_0[7]), .B(p_1[7]), .CI(n_6), .CO(n_7), .S(divider[7]));
   FA_X1 i_8 (.A(p_0[8]), .B(p_1[8]), .CI(n_7), .CO(n_8), .S(divider[8]));
   FA_X1 i_9 (.A(p_0[9]), .B(p_1[9]), .CI(n_8), .CO(n_9), .S(divider[9]));
   FA_X1 i_10 (.A(p_0[10]), .B(p_1[10]), .CI(n_9), .CO(n_10), .S(divider[10]));
   FA_X1 i_11 (.A(p_0[11]), .B(p_1[11]), .CI(n_10), .CO(n_11), .S(divider[11]));
   FA_X1 i_12 (.A(p_0[12]), .B(p_1[12]), .CI(n_11), .CO(n_12), .S(divider[12]));
   FA_X1 i_13 (.A(p_0[13]), .B(p_1[13]), .CI(n_12), .CO(n_13), .S(divider[13]));
   FA_X1 i_14 (.A(p_0[14]), .B(p_1[14]), .CI(n_13), .CO(n_14), .S(divider[14]));
   FA_X1 i_15 (.A(p_0[15]), .B(p_1[15]), .CI(n_14), .CO(n_15), .S(divider[15]));
   FA_X1 i_16 (.A(p_0[16]), .B(p_1[16]), .CI(n_15), .CO(n_16), .S(divider[16]));
   FA_X1 i_17 (.A(p_0[17]), .B(p_1[17]), .CI(n_16), .CO(n_17), .S(divider[17]));
   FA_X1 i_18 (.A(p_0[18]), .B(p_1[18]), .CI(n_17), .CO(n_18), .S(divider[18]));
   FA_X1 i_19 (.A(p_0[19]), .B(p_1[19]), .CI(n_18), .CO(n_19), .S(divider[19]));
   FA_X1 i_20 (.A(p_0[20]), .B(p_1[20]), .CI(n_19), .CO(n_20), .S(divider[20]));
   FA_X1 i_21 (.A(p_0[21]), .B(p_1[21]), .CI(n_20), .CO(n_21), .S(divider[21]));
endmodule

module datapath__0_69(p_0, p_1, divider);
   input [22:0]p_0;
   input [22:0]p_1;
   output [22:0]divider;

   HA_X1 i_0 (.A(p_0[0]), .B(p_1[0]), .CO(n_0), .S(divider[0]));
   FA_X1 i_1 (.A(p_0[1]), .B(p_1[1]), .CI(n_0), .CO(n_1), .S(divider[1]));
   FA_X1 i_2 (.A(p_0[2]), .B(p_1[2]), .CI(n_1), .CO(n_2), .S(divider[2]));
   FA_X1 i_3 (.A(p_0[3]), .B(p_1[3]), .CI(n_2), .CO(n_3), .S(divider[3]));
   FA_X1 i_4 (.A(p_0[4]), .B(p_1[4]), .CI(n_3), .CO(n_4), .S(divider[4]));
   FA_X1 i_5 (.A(p_0[5]), .B(p_1[5]), .CI(n_4), .CO(n_5), .S(divider[5]));
   FA_X1 i_6 (.A(p_0[6]), .B(p_1[6]), .CI(n_5), .CO(n_6), .S(divider[6]));
   FA_X1 i_7 (.A(p_0[7]), .B(p_1[7]), .CI(n_6), .CO(n_7), .S(divider[7]));
   FA_X1 i_8 (.A(p_0[8]), .B(p_1[8]), .CI(n_7), .CO(n_8), .S(divider[8]));
   FA_X1 i_9 (.A(p_0[9]), .B(p_1[9]), .CI(n_8), .CO(n_9), .S(divider[9]));
   FA_X1 i_10 (.A(p_0[10]), .B(p_1[10]), .CI(n_9), .CO(n_10), .S(divider[10]));
   FA_X1 i_11 (.A(p_0[11]), .B(p_1[11]), .CI(n_10), .CO(n_11), .S(divider[11]));
   FA_X1 i_12 (.A(p_0[12]), .B(p_1[12]), .CI(n_11), .CO(n_12), .S(divider[12]));
   FA_X1 i_13 (.A(p_0[13]), .B(p_1[13]), .CI(n_12), .CO(n_13), .S(divider[13]));
   FA_X1 i_14 (.A(p_0[14]), .B(p_1[14]), .CI(n_13), .CO(n_14), .S(divider[14]));
   FA_X1 i_15 (.A(p_0[15]), .B(p_1[15]), .CI(n_14), .CO(n_15), .S(divider[15]));
   FA_X1 i_16 (.A(p_0[16]), .B(p_1[16]), .CI(n_15), .CO(n_16), .S(divider[16]));
   FA_X1 i_17 (.A(p_0[17]), .B(p_1[17]), .CI(n_16), .CO(n_17), .S(divider[17]));
   FA_X1 i_18 (.A(p_0[18]), .B(p_1[18]), .CI(n_17), .CO(n_18), .S(divider[18]));
   FA_X1 i_19 (.A(p_0[19]), .B(p_1[19]), .CI(n_18), .CO(n_19), .S(divider[19]));
   FA_X1 i_20 (.A(p_0[20]), .B(p_1[20]), .CI(n_19), .CO(n_20), .S(divider[20]));
   FA_X1 i_21 (.A(p_0[21]), .B(p_1[21]), .CI(n_20), .CO(n_21), .S(divider[21]));
endmodule

module datapath__0_73(p_0, p_1, divider);
   input [22:0]p_0;
   input [22:0]p_1;
   output [22:0]divider;

   HA_X1 i_0 (.A(p_0[1]), .B(p_1[1]), .CO(n_0), .S(divider[1]));
   FA_X1 i_1 (.A(p_0[2]), .B(p_1[2]), .CI(n_0), .CO(n_1), .S(divider[2]));
   FA_X1 i_2 (.A(p_0[3]), .B(p_1[3]), .CI(n_1), .CO(n_2), .S(divider[3]));
   FA_X1 i_3 (.A(p_0[4]), .B(p_1[4]), .CI(n_2), .CO(n_3), .S(divider[4]));
   FA_X1 i_4 (.A(p_0[5]), .B(p_1[5]), .CI(n_3), .CO(n_4), .S(divider[5]));
   FA_X1 i_5 (.A(p_0[6]), .B(p_1[6]), .CI(n_4), .CO(n_5), .S(divider[6]));
   FA_X1 i_6 (.A(p_0[7]), .B(p_1[7]), .CI(n_5), .CO(n_6), .S(divider[7]));
   FA_X1 i_7 (.A(p_0[8]), .B(p_1[8]), .CI(n_6), .CO(n_7), .S(divider[8]));
   FA_X1 i_8 (.A(p_0[9]), .B(p_1[9]), .CI(n_7), .CO(n_8), .S(divider[9]));
   FA_X1 i_9 (.A(p_0[10]), .B(p_1[10]), .CI(n_8), .CO(n_9), .S(divider[10]));
   FA_X1 i_10 (.A(p_0[11]), .B(p_1[11]), .CI(n_9), .CO(n_10), .S(divider[11]));
   FA_X1 i_11 (.A(p_0[12]), .B(p_1[12]), .CI(n_10), .CO(n_11), .S(divider[12]));
   FA_X1 i_12 (.A(p_0[13]), .B(p_1[13]), .CI(n_11), .CO(n_12), .S(divider[13]));
   FA_X1 i_13 (.A(p_0[14]), .B(p_1[14]), .CI(n_12), .CO(n_13), .S(divider[14]));
   FA_X1 i_14 (.A(p_0[15]), .B(p_1[15]), .CI(n_13), .CO(n_14), .S(divider[15]));
   FA_X1 i_15 (.A(p_0[16]), .B(p_1[16]), .CI(n_14), .CO(n_15), .S(divider[16]));
   FA_X1 i_16 (.A(p_0[17]), .B(p_1[17]), .CI(n_15), .CO(n_16), .S(divider[17]));
   FA_X1 i_17 (.A(p_0[18]), .B(p_1[18]), .CI(n_16), .CO(n_17), .S(divider[18]));
   FA_X1 i_18 (.A(p_0[19]), .B(p_1[19]), .CI(n_17), .CO(n_18), .S(divider[19]));
   FA_X1 i_19 (.A(p_0[20]), .B(p_1[20]), .CI(n_18), .CO(n_19), .S(divider[20]));
   FA_X1 i_20 (.A(p_0[21]), .B(p_1[21]), .CI(n_19), .CO(n_20), .S(divider[21]));
endmodule

module datapath__0_77(p_0, p_1, divider);
   input [22:0]p_0;
   input [22:0]p_1;
   output [22:0]divider;

   HA_X1 i_0 (.A(p_0[1]), .B(p_1[1]), .CO(n_0), .S(divider[1]));
   FA_X1 i_1 (.A(p_0[2]), .B(p_1[2]), .CI(n_0), .CO(n_1), .S(divider[2]));
   FA_X1 i_2 (.A(p_0[3]), .B(p_1[3]), .CI(n_1), .CO(n_2), .S(divider[3]));
   FA_X1 i_3 (.A(p_0[4]), .B(p_1[4]), .CI(n_2), .CO(n_3), .S(divider[4]));
   FA_X1 i_4 (.A(p_0[5]), .B(p_1[5]), .CI(n_3), .CO(n_4), .S(divider[5]));
   FA_X1 i_5 (.A(p_0[6]), .B(p_1[6]), .CI(n_4), .CO(n_5), .S(divider[6]));
   FA_X1 i_6 (.A(p_0[7]), .B(p_1[7]), .CI(n_5), .CO(n_6), .S(divider[7]));
   FA_X1 i_7 (.A(p_0[8]), .B(p_1[8]), .CI(n_6), .CO(n_7), .S(divider[8]));
   FA_X1 i_8 (.A(p_0[9]), .B(p_1[9]), .CI(n_7), .CO(n_8), .S(divider[9]));
   FA_X1 i_9 (.A(p_0[10]), .B(p_1[10]), .CI(n_8), .CO(n_9), .S(divider[10]));
   FA_X1 i_10 (.A(p_0[11]), .B(p_1[11]), .CI(n_9), .CO(n_10), .S(divider[11]));
   FA_X1 i_11 (.A(p_0[12]), .B(p_1[12]), .CI(n_10), .CO(n_11), .S(divider[12]));
   FA_X1 i_12 (.A(p_0[13]), .B(p_1[13]), .CI(n_11), .CO(n_12), .S(divider[13]));
   FA_X1 i_13 (.A(p_0[14]), .B(p_1[14]), .CI(n_12), .CO(n_13), .S(divider[14]));
   FA_X1 i_14 (.A(p_0[15]), .B(p_1[15]), .CI(n_13), .CO(n_14), .S(divider[15]));
   FA_X1 i_15 (.A(p_0[16]), .B(p_1[16]), .CI(n_14), .CO(n_15), .S(divider[16]));
   FA_X1 i_16 (.A(p_0[17]), .B(p_1[17]), .CI(n_15), .CO(n_16), .S(divider[17]));
   FA_X1 i_17 (.A(p_0[18]), .B(p_1[18]), .CI(n_16), .CO(n_17), .S(divider[18]));
   FA_X1 i_18 (.A(p_0[19]), .B(p_1[19]), .CI(n_17), .CO(n_18), .S(divider[19]));
   FA_X1 i_19 (.A(p_0[20]), .B(p_1[20]), .CI(n_18), .CO(n_19), .S(divider[20]));
   FA_X1 i_20 (.A(p_0[21]), .B(p_1[21]), .CI(n_19), .CO(n_20), .S(divider[21]));
endmodule

module datapath__0_81(p_0, p_1, divider);
   input [22:0]p_0;
   input [22:0]p_1;
   output [22:0]divider;

   HA_X1 i_0 (.A(p_0[1]), .B(p_1[1]), .CO(n_0), .S(divider[1]));
   FA_X1 i_1 (.A(p_0[2]), .B(p_1[2]), .CI(n_0), .CO(n_1), .S(divider[2]));
   FA_X1 i_2 (.A(p_0[3]), .B(p_1[3]), .CI(n_1), .CO(n_2), .S(divider[3]));
   FA_X1 i_3 (.A(p_0[4]), .B(p_1[4]), .CI(n_2), .CO(n_3), .S(divider[4]));
   FA_X1 i_4 (.A(p_0[5]), .B(p_1[5]), .CI(n_3), .CO(n_4), .S(divider[5]));
   FA_X1 i_5 (.A(p_0[6]), .B(p_1[6]), .CI(n_4), .CO(n_5), .S(divider[6]));
   FA_X1 i_6 (.A(p_0[7]), .B(p_1[7]), .CI(n_5), .CO(n_6), .S(divider[7]));
   FA_X1 i_7 (.A(p_0[8]), .B(p_1[8]), .CI(n_6), .CO(n_7), .S(divider[8]));
   FA_X1 i_8 (.A(p_0[9]), .B(p_1[9]), .CI(n_7), .CO(n_8), .S(divider[9]));
   FA_X1 i_9 (.A(p_0[10]), .B(p_1[10]), .CI(n_8), .CO(n_9), .S(divider[10]));
   FA_X1 i_10 (.A(p_0[11]), .B(p_1[11]), .CI(n_9), .CO(n_10), .S(divider[11]));
   FA_X1 i_11 (.A(p_0[12]), .B(p_1[12]), .CI(n_10), .CO(n_11), .S(divider[12]));
   FA_X1 i_12 (.A(p_0[13]), .B(p_1[13]), .CI(n_11), .CO(n_12), .S(divider[13]));
   FA_X1 i_13 (.A(p_0[14]), .B(p_1[14]), .CI(n_12), .CO(n_13), .S(divider[14]));
   FA_X1 i_14 (.A(p_0[15]), .B(p_1[15]), .CI(n_13), .CO(n_14), .S(divider[15]));
   FA_X1 i_15 (.A(p_0[16]), .B(p_1[16]), .CI(n_14), .CO(n_15), .S(divider[16]));
   FA_X1 i_16 (.A(p_0[17]), .B(p_1[17]), .CI(n_15), .CO(n_16), .S(divider[17]));
   FA_X1 i_17 (.A(p_0[18]), .B(p_1[18]), .CI(n_16), .CO(n_17), .S(divider[18]));
   FA_X1 i_18 (.A(p_0[19]), .B(p_1[19]), .CI(n_17), .CO(n_18), .S(divider[19]));
   FA_X1 i_19 (.A(p_0[20]), .B(p_1[20]), .CI(n_18), .CO(n_19), .S(divider[20]));
   FA_X1 i_20 (.A(p_0[21]), .B(p_1[21]), .CI(n_19), .CO(n_20), .S(divider[21]));
endmodule

module datapath__0_85(p_0, p_1, divider);
   input [22:0]p_0;
   input [22:0]p_1;
   output [22:0]divider;

   HA_X1 i_0 (.A(p_0[1]), .B(p_1[1]), .CO(n_0), .S(divider[1]));
   FA_X1 i_1 (.A(p_0[2]), .B(p_1[2]), .CI(n_0), .CO(n_1), .S(divider[2]));
   FA_X1 i_2 (.A(p_0[3]), .B(p_1[3]), .CI(n_1), .CO(n_2), .S(divider[3]));
   FA_X1 i_3 (.A(p_0[4]), .B(p_1[4]), .CI(n_2), .CO(n_3), .S(divider[4]));
   FA_X1 i_4 (.A(p_0[5]), .B(p_1[5]), .CI(n_3), .CO(n_4), .S(divider[5]));
   FA_X1 i_5 (.A(p_0[6]), .B(p_1[6]), .CI(n_4), .CO(n_5), .S(divider[6]));
   FA_X1 i_6 (.A(p_0[7]), .B(p_1[7]), .CI(n_5), .CO(n_6), .S(divider[7]));
   FA_X1 i_7 (.A(p_0[8]), .B(p_1[8]), .CI(n_6), .CO(n_7), .S(divider[8]));
   FA_X1 i_8 (.A(p_0[9]), .B(p_1[9]), .CI(n_7), .CO(n_8), .S(divider[9]));
   FA_X1 i_9 (.A(p_0[10]), .B(p_1[10]), .CI(n_8), .CO(n_9), .S(divider[10]));
   FA_X1 i_10 (.A(p_0[11]), .B(p_1[11]), .CI(n_9), .CO(n_10), .S(divider[11]));
   FA_X1 i_11 (.A(p_0[12]), .B(p_1[12]), .CI(n_10), .CO(n_11), .S(divider[12]));
   FA_X1 i_12 (.A(p_0[13]), .B(p_1[13]), .CI(n_11), .CO(n_12), .S(divider[13]));
   FA_X1 i_13 (.A(p_0[14]), .B(p_1[14]), .CI(n_12), .CO(n_13), .S(divider[14]));
   FA_X1 i_14 (.A(p_0[15]), .B(p_1[15]), .CI(n_13), .CO(n_14), .S(divider[15]));
   FA_X1 i_15 (.A(p_0[16]), .B(p_1[16]), .CI(n_14), .CO(n_15), .S(divider[16]));
   FA_X1 i_16 (.A(p_0[17]), .B(p_1[17]), .CI(n_15), .CO(n_16), .S(divider[17]));
   FA_X1 i_17 (.A(p_0[18]), .B(p_1[18]), .CI(n_16), .CO(n_17), .S(divider[18]));
   FA_X1 i_18 (.A(p_0[19]), .B(p_1[19]), .CI(n_17), .CO(n_18), .S(divider[19]));
   FA_X1 i_19 (.A(p_0[20]), .B(p_1[20]), .CI(n_18), .CO(n_19), .S(divider[20]));
   FA_X1 i_20 (.A(p_0[21]), .B(p_1[21]), .CI(n_19), .CO(n_20), .S(divider[21]));
endmodule

module datapath__0_89(p_0, p_1, divider);
   input [22:0]p_0;
   input [22:0]p_1;
   output [22:0]divider;

   HA_X1 i_0 (.A(p_0[1]), .B(p_1[1]), .CO(n_0), .S(divider[1]));
   FA_X1 i_1 (.A(p_0[2]), .B(p_1[2]), .CI(n_0), .CO(n_1), .S(divider[2]));
   FA_X1 i_2 (.A(p_0[3]), .B(p_1[3]), .CI(n_1), .CO(n_2), .S(divider[3]));
   FA_X1 i_3 (.A(p_0[4]), .B(p_1[4]), .CI(n_2), .CO(n_3), .S(divider[4]));
   FA_X1 i_4 (.A(p_0[5]), .B(p_1[5]), .CI(n_3), .CO(n_4), .S(divider[5]));
   FA_X1 i_5 (.A(p_0[6]), .B(p_1[6]), .CI(n_4), .CO(n_5), .S(divider[6]));
   FA_X1 i_6 (.A(p_0[7]), .B(p_1[7]), .CI(n_5), .CO(n_6), .S(divider[7]));
   FA_X1 i_7 (.A(p_0[8]), .B(p_1[8]), .CI(n_6), .CO(n_7), .S(divider[8]));
   FA_X1 i_8 (.A(p_0[9]), .B(p_1[9]), .CI(n_7), .CO(n_8), .S(divider[9]));
   FA_X1 i_9 (.A(p_0[10]), .B(p_1[10]), .CI(n_8), .CO(n_9), .S(divider[10]));
   FA_X1 i_10 (.A(p_0[11]), .B(p_1[11]), .CI(n_9), .CO(n_10), .S(divider[11]));
   FA_X1 i_11 (.A(p_0[12]), .B(p_1[12]), .CI(n_10), .CO(n_11), .S(divider[12]));
   FA_X1 i_12 (.A(p_0[13]), .B(p_1[13]), .CI(n_11), .CO(n_12), .S(divider[13]));
   FA_X1 i_13 (.A(p_0[14]), .B(p_1[14]), .CI(n_12), .CO(n_13), .S(divider[14]));
   FA_X1 i_14 (.A(p_0[15]), .B(p_1[15]), .CI(n_13), .CO(n_14), .S(divider[15]));
   FA_X1 i_15 (.A(p_0[16]), .B(p_1[16]), .CI(n_14), .CO(n_15), .S(divider[16]));
   FA_X1 i_16 (.A(p_0[17]), .B(p_1[17]), .CI(n_15), .CO(n_16), .S(divider[17]));
   FA_X1 i_17 (.A(p_0[18]), .B(p_1[18]), .CI(n_16), .CO(n_17), .S(divider[18]));
   FA_X1 i_18 (.A(p_0[19]), .B(p_1[19]), .CI(n_17), .CO(n_18), .S(divider[19]));
   FA_X1 i_19 (.A(p_0[20]), .B(p_1[20]), .CI(n_18), .CO(n_19), .S(divider[20]));
   FA_X1 i_20 (.A(p_0[21]), .B(p_1[21]), .CI(n_19), .CO(n_20), .S(divider[21]));
endmodule

module datapath__0_93(p_0, p_1, divider);
   input [22:0]p_0;
   input [22:0]p_1;
   output [22:0]divider;

   HA_X1 i_0 (.A(p_0[1]), .B(p_1[1]), .CO(n_0), .S(divider[1]));
   FA_X1 i_1 (.A(p_0[2]), .B(p_1[2]), .CI(n_0), .CO(n_1), .S(divider[2]));
   FA_X1 i_2 (.A(p_0[3]), .B(p_1[3]), .CI(n_1), .CO(n_2), .S(divider[3]));
   FA_X1 i_3 (.A(p_0[4]), .B(p_1[4]), .CI(n_2), .CO(n_3), .S(divider[4]));
   FA_X1 i_4 (.A(p_0[5]), .B(p_1[5]), .CI(n_3), .CO(n_4), .S(divider[5]));
   FA_X1 i_5 (.A(p_0[6]), .B(p_1[6]), .CI(n_4), .CO(n_5), .S(divider[6]));
   FA_X1 i_6 (.A(p_0[7]), .B(p_1[7]), .CI(n_5), .CO(n_6), .S(divider[7]));
   FA_X1 i_7 (.A(p_0[8]), .B(p_1[8]), .CI(n_6), .CO(n_7), .S(divider[8]));
   FA_X1 i_8 (.A(p_0[9]), .B(p_1[9]), .CI(n_7), .CO(n_8), .S(divider[9]));
   FA_X1 i_9 (.A(p_0[10]), .B(p_1[10]), .CI(n_8), .CO(n_9), .S(divider[10]));
   FA_X1 i_10 (.A(p_0[11]), .B(p_1[11]), .CI(n_9), .CO(n_10), .S(divider[11]));
   FA_X1 i_11 (.A(p_0[12]), .B(p_1[12]), .CI(n_10), .CO(n_11), .S(divider[12]));
   FA_X1 i_12 (.A(p_0[13]), .B(p_1[13]), .CI(n_11), .CO(n_12), .S(divider[13]));
   FA_X1 i_13 (.A(p_0[14]), .B(p_1[14]), .CI(n_12), .CO(n_13), .S(divider[14]));
   FA_X1 i_14 (.A(p_0[15]), .B(p_1[15]), .CI(n_13), .CO(n_14), .S(divider[15]));
   FA_X1 i_15 (.A(p_0[16]), .B(p_1[16]), .CI(n_14), .CO(n_15), .S(divider[16]));
   FA_X1 i_16 (.A(p_0[17]), .B(p_1[17]), .CI(n_15), .CO(n_16), .S(divider[17]));
   FA_X1 i_17 (.A(p_0[18]), .B(p_1[18]), .CI(n_16), .CO(n_17), .S(divider[18]));
   FA_X1 i_18 (.A(p_0[19]), .B(p_1[19]), .CI(n_17), .CO(n_18), .S(divider[19]));
   FA_X1 i_19 (.A(p_0[20]), .B(p_1[20]), .CI(n_18), .CO(n_19), .S(divider[20]));
   FA_X1 i_20 (.A(p_0[21]), .B(p_1[21]), .CI(n_19), .CO(n_20), .S(divider[21]));
endmodule

module datapath__0_103(plus, p_0);
   output [63:0]plus;
   input [63:0]p_0;

   XOR2_X1 i_0 (.A(p_0[1]), .B(p_0[0]), .Z(plus[1]));
   AND2_X1 i_1 (.A1(n_13), .A2(n_0), .ZN(plus[2]));
   OAI21_X1 i_2 (.A(p_0[2]), .B1(p_0[1]), .B2(p_0[0]), .ZN(n_0));
   XOR2_X1 i_3 (.A(p_0[3]), .B(n_13), .Z(plus[3]));
   XOR2_X1 i_4 (.A(p_0[4]), .B(n_12), .Z(plus[4]));
   XOR2_X1 i_5 (.A(p_0[5]), .B(n_11), .Z(plus[5]));
   AND2_X1 i_6 (.A1(n_10), .A2(n_1), .ZN(plus[6]));
   OAI21_X1 i_7 (.A(p_0[6]), .B1(n_11), .B2(p_0[5]), .ZN(n_1));
   XOR2_X1 i_8 (.A(p_0[7]), .B(n_10), .Z(plus[7]));
   XOR2_X1 i_9 (.A(p_0[8]), .B(n_9), .Z(plus[8]));
   AND2_X1 i_10 (.A1(n_8), .A2(n_2), .ZN(plus[9]));
   OAI21_X1 i_11 (.A(p_0[9]), .B1(n_9), .B2(p_0[8]), .ZN(n_2));
   XOR2_X1 i_12 (.A(p_0[10]), .B(n_8), .Z(plus[10]));
   XOR2_X1 i_13 (.A(p_0[11]), .B(n_7), .Z(plus[11]));
   XOR2_X1 i_14 (.A(p_0[12]), .B(n_6), .Z(plus[12]));
   XNOR2_X1 i_15 (.A(p_0[13]), .B(n_5), .ZN(plus[13]));
   XOR2_X1 i_16 (.A(p_0[14]), .B(n_4), .Z(plus[14]));
   AND2_X1 i_17 (.A1(plus[63]), .A2(n_3), .ZN(plus[15]));
   OAI21_X1 i_18 (.A(p_0[15]), .B1(n_4), .B2(p_0[14]), .ZN(n_3));
   OR3_X1 i_19 (.A1(n_4), .A2(p_0[14]), .A3(p_0[15]), .ZN(plus[63]));
   NAND2_X1 i_20 (.A1(n_5), .A2(n_14), .ZN(n_4));
   NOR2_X1 i_21 (.A1(n_6), .A2(p_0[12]), .ZN(n_5));
   OR2_X1 i_22 (.A1(n_7), .A2(p_0[11]), .ZN(n_6));
   OR2_X1 i_23 (.A1(n_8), .A2(p_0[10]), .ZN(n_7));
   OR3_X1 i_24 (.A1(n_9), .A2(p_0[8]), .A3(p_0[9]), .ZN(n_8));
   OR2_X1 i_25 (.A1(n_10), .A2(p_0[7]), .ZN(n_9));
   OR3_X1 i_26 (.A1(n_11), .A2(p_0[5]), .A3(p_0[6]), .ZN(n_10));
   OR2_X1 i_27 (.A1(n_12), .A2(p_0[4]), .ZN(n_11));
   OR2_X1 i_28 (.A1(n_13), .A2(p_0[3]), .ZN(n_12));
   OR3_X1 i_29 (.A1(p_0[2]), .A2(p_0[1]), .A3(p_0[0]), .ZN(n_13));
   INV_X1 i_30 (.A(p_0[13]), .ZN(n_14));
endmodule

module fpu_divider(mode, clk, rst, enbl, in_a, in_b, out_c, done, err, zero, 
      posv);
   input [1:0]mode;
   input clk;
   input rst;
   input enbl;
   input [63:0]in_a;
   input [63:0]in_b;
   output [63:0]out_c;
   output done;
   output err;
   output zero;
   output posv;

   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_4;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire [22:0]divider;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_189;
   wire n_0_190;
   wire n_0_191;
   wire n_0_192;
   wire n_0_193;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_200;
   wire n_0_201;
   wire n_0_202;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_207;
   wire n_0_208;
   wire n_0_209;
   wire n_0_210;
   wire n_0_234;
   wire n_0_235;
   wire n_0_236;
   wire n_0_237;
   wire n_0_238;
   wire n_0_239;
   wire n_0_240;
   wire n_0_241;
   wire n_0_242;
   wire n_0_243;
   wire n_0_244;
   wire n_0_245;
   wire n_0_246;
   wire n_0_247;
   wire n_0_248;
   wire n_0_249;
   wire n_0_250;
   wire n_0_251;
   wire n_0_252;
   wire n_0_253;
   wire n_0_254;
   wire n_0_255;
   wire n_0_279;
   wire n_0_280;
   wire n_0_281;
   wire n_0_282;
   wire n_0_283;
   wire n_0_284;
   wire n_0_285;
   wire n_0_286;
   wire n_0_287;
   wire n_0_288;
   wire n_0_289;
   wire n_0_290;
   wire n_0_291;
   wire n_0_292;
   wire n_0_293;
   wire n_0_294;
   wire n_0_295;
   wire n_0_296;
   wire n_0_297;
   wire n_0_298;
   wire n_0_299;
   wire n_0_300;
   wire n_0_324;
   wire n_0_325;
   wire n_0_326;
   wire n_0_327;
   wire n_0_328;
   wire n_0_329;
   wire n_0_330;
   wire n_0_331;
   wire n_0_332;
   wire n_0_333;
   wire n_0_334;
   wire n_0_335;
   wire n_0_336;
   wire n_0_337;
   wire n_0_338;
   wire n_0_339;
   wire n_0_340;
   wire n_0_341;
   wire n_0_342;
   wire n_0_343;
   wire n_0_344;
   wire n_0_345;
   wire n_0_369;
   wire n_0_370;
   wire n_0_371;
   wire n_0_372;
   wire n_0_373;
   wire n_0_374;
   wire n_0_375;
   wire n_0_376;
   wire n_0_377;
   wire n_0_378;
   wire n_0_379;
   wire n_0_380;
   wire n_0_381;
   wire n_0_382;
   wire n_0_383;
   wire n_0_384;
   wire n_0_385;
   wire n_0_386;
   wire n_0_387;
   wire n_0_388;
   wire n_0_389;
   wire n_0_390;
   wire n_0_414;
   wire n_0_415;
   wire n_0_416;
   wire n_0_417;
   wire n_0_418;
   wire n_0_419;
   wire n_0_420;
   wire n_0_421;
   wire n_0_422;
   wire n_0_423;
   wire n_0_424;
   wire n_0_425;
   wire n_0_426;
   wire n_0_427;
   wire n_0_428;
   wire n_0_429;
   wire n_0_430;
   wire n_0_431;
   wire n_0_432;
   wire n_0_433;
   wire n_0_434;
   wire n_0_435;
   wire n_0_459;
   wire n_0_460;
   wire n_0_461;
   wire n_0_462;
   wire n_0_463;
   wire n_0_464;
   wire n_0_465;
   wire n_0_466;
   wire n_0_467;
   wire n_0_468;
   wire n_0_469;
   wire n_0_470;
   wire n_0_471;
   wire n_0_472;
   wire n_0_473;
   wire n_0_474;
   wire n_0_475;
   wire n_0_476;
   wire n_0_477;
   wire n_0_478;
   wire n_0_479;
   wire n_0_480;
   wire n_0_504;
   wire n_0_505;
   wire n_0_506;
   wire n_0_507;
   wire n_0_508;
   wire n_0_509;
   wire n_0_510;
   wire n_0_511;
   wire n_0_512;
   wire n_0_513;
   wire n_0_514;
   wire n_0_515;
   wire n_0_516;
   wire n_0_517;
   wire n_0_518;
   wire n_0_519;
   wire n_0_520;
   wire n_0_521;
   wire n_0_522;
   wire n_0_523;
   wire n_0_524;
   wire n_0_525;
   wire n_0_549;
   wire n_0_550;
   wire n_0_551;
   wire n_0_552;
   wire n_0_553;
   wire n_0_554;
   wire n_0_555;
   wire n_0_556;
   wire n_0_557;
   wire n_0_558;
   wire n_0_559;
   wire n_0_560;
   wire n_0_561;
   wire n_0_562;
   wire n_0_563;
   wire n_0_564;
   wire n_0_565;
   wire n_0_566;
   wire n_0_567;
   wire n_0_568;
   wire n_0_569;
   wire n_0_570;
   wire n_0_594;
   wire n_0_595;
   wire n_0_596;
   wire n_0_597;
   wire n_0_598;
   wire n_0_599;
   wire n_0_600;
   wire n_0_601;
   wire n_0_602;
   wire n_0_603;
   wire n_0_604;
   wire n_0_605;
   wire n_0_606;
   wire n_0_607;
   wire n_0_608;
   wire n_0_609;
   wire n_0_610;
   wire n_0_611;
   wire n_0_612;
   wire n_0_613;
   wire n_0_614;
   wire n_0_615;
   wire n_0_639;
   wire n_0_640;
   wire n_0_641;
   wire n_0_642;
   wire n_0_643;
   wire n_0_644;
   wire n_0_645;
   wire n_0_646;
   wire n_0_647;
   wire n_0_648;
   wire n_0_649;
   wire n_0_650;
   wire n_0_651;
   wire n_0_652;
   wire n_0_653;
   wire n_0_654;
   wire n_0_655;
   wire n_0_656;
   wire n_0_657;
   wire n_0_658;
   wire n_0_659;
   wire n_0_660;
   wire n_0_684;
   wire n_0_685;
   wire n_0_686;
   wire n_0_687;
   wire n_0_688;
   wire n_0_689;
   wire n_0_690;
   wire n_0_691;
   wire n_0_692;
   wire n_0_693;
   wire n_0_694;
   wire n_0_695;
   wire n_0_696;
   wire n_0_697;
   wire n_0_698;
   wire n_0_699;
   wire n_0_700;
   wire n_0_701;
   wire n_0_702;
   wire n_0_703;
   wire n_0_704;
   wire n_0_705;
   wire n_0_729;
   wire n_0_730;
   wire n_0_731;
   wire n_0_732;
   wire n_0_733;
   wire n_0_734;
   wire n_0_735;
   wire n_0_736;
   wire n_0_737;
   wire n_0_738;
   wire n_0_739;
   wire n_0_740;
   wire n_0_741;
   wire n_0_742;
   wire n_0_743;
   wire n_0_744;
   wire n_0_745;
   wire n_0_746;
   wire n_0_747;
   wire n_0_748;
   wire n_0_749;
   wire n_0_750;
   wire n_0_774;
   wire n_0_775;
   wire n_0_776;
   wire n_0_777;
   wire n_0_778;
   wire n_0_779;
   wire n_0_780;
   wire n_0_781;
   wire n_0_782;
   wire n_0_783;
   wire n_0_784;
   wire n_0_785;
   wire n_0_786;
   wire n_0_787;
   wire n_0_788;
   wire n_0_789;
   wire n_0_790;
   wire n_0_791;
   wire n_0_792;
   wire n_0_793;
   wire n_0_794;
   wire n_0_795;
   wire n_0_819;
   wire n_0_820;
   wire n_0_821;
   wire n_0_822;
   wire n_0_823;
   wire n_0_824;
   wire n_0_825;
   wire n_0_826;
   wire n_0_827;
   wire n_0_828;
   wire n_0_829;
   wire n_0_830;
   wire n_0_831;
   wire n_0_832;
   wire n_0_833;
   wire n_0_834;
   wire n_0_835;
   wire n_0_836;
   wire n_0_837;
   wire n_0_838;
   wire n_0_839;
   wire n_0_863;
   wire n_0_864;
   wire n_0_865;
   wire n_0_866;
   wire n_0_867;
   wire n_0_868;
   wire n_0_869;
   wire n_0_870;
   wire n_0_871;
   wire n_0_872;
   wire n_0_873;
   wire n_0_874;
   wire n_0_875;
   wire n_0_876;
   wire n_0_877;
   wire n_0_878;
   wire n_0_879;
   wire n_0_880;
   wire n_0_881;
   wire n_0_882;
   wire n_0_883;
   wire n_0_907;
   wire n_0_908;
   wire n_0_909;
   wire n_0_910;
   wire n_0_911;
   wire n_0_912;
   wire n_0_913;
   wire n_0_914;
   wire n_0_915;
   wire n_0_916;
   wire n_0_917;
   wire n_0_918;
   wire n_0_919;
   wire n_0_920;
   wire n_0_921;
   wire n_0_922;
   wire n_0_923;
   wire n_0_924;
   wire n_0_925;
   wire n_0_926;
   wire n_0_927;
   wire n_0_951;
   wire n_0_952;
   wire n_0_953;
   wire n_0_954;
   wire n_0_955;
   wire n_0_956;
   wire n_0_957;
   wire n_0_958;
   wire n_0_959;
   wire n_0_960;
   wire n_0_961;
   wire n_0_962;
   wire n_0_963;
   wire n_0_964;
   wire n_0_965;
   wire n_0_966;
   wire n_0_967;
   wire n_0_968;
   wire n_0_969;
   wire n_0_970;
   wire n_0_971;
   wire n_0_995;
   wire n_0_996;
   wire n_0_997;
   wire n_0_998;
   wire n_0_999;
   wire n_0_1000;
   wire n_0_1001;
   wire n_0_1002;
   wire n_0_1003;
   wire n_0_1004;
   wire n_0_1005;
   wire n_0_1006;
   wire n_0_1007;
   wire n_0_1008;
   wire n_0_1009;
   wire n_0_1010;
   wire n_0_1011;
   wire n_0_1012;
   wire n_0_1013;
   wire n_0_1014;
   wire n_0_1015;
   wire n_0_1039;
   wire n_0_1040;
   wire n_0_1041;
   wire n_0_1042;
   wire n_0_1043;
   wire n_0_1044;
   wire n_0_1045;
   wire n_0_1046;
   wire n_0_1047;
   wire n_0_1048;
   wire n_0_1049;
   wire n_0_1050;
   wire n_0_1051;
   wire n_0_1052;
   wire n_0_1053;
   wire n_0_1054;
   wire n_0_1055;
   wire n_0_1056;
   wire n_0_1057;
   wire n_0_1058;
   wire n_0_1059;
   wire n_0_0;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire ovfl_flag;
   wire divide_by_zero_error;
   wire n_0_1065;
   wire n_0_38;
   wire n_0_40;
   wire n_0_0_0;
   wire n_0_0_1;
   wire n_0_0_2;
   wire n_0_0_3;
   wire n_0_0_4;
   wire n_0_0_5;
   wire n_0_0_6;
   wire n_0_0_7;
   wire n_0_0_8;
   wire n_0_0_9;
   wire n_0_0_10;
   wire n_0_0_11;
   wire n_0_0_12;
   wire n_0_0_13;
   wire n_0_0_14;
   wire n_0_0_15;
   wire n_0_0_16;
   wire n_0_0_17;
   wire n_0_0_18;
   wire n_0_0_19;
   wire n_0_0_20;
   wire n_0_41;
   wire n_0_0_21;
   wire n_0_42;
   wire n_0_43;
   wire n_0_0_22;
   wire n_0_0_23;
   wire n_0_0_24;
   wire n_0_0_25;
   wire n_0_0_26;
   wire n_0_0_27;
   wire n_0_0_28;
   wire n_0_0_29;
   wire n_0_0_30;
   wire n_0_0_31;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_0_32;
   wire n_0_48;
   wire n_0_0_33;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_0_34;
   wire n_0_52;
   wire n_0_53;
   wire n_0_0_35;
   wire n_0_54;
   wire n_0_0_36;
   wire n_0_55;
   wire n_0_0_37;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_0_38;
   wire n_0_0_39;
   wire n_0_0_40;
   wire n_0_59;
   wire n_0_0_41;
   wire n_0_1066;
   wire n_0_0_42;
   wire n_0_0_43;
   wire n_0_0_44;
   wire n_0_0_45;
   wire n_0_0_46;
   wire n_0_0_47;
   wire n_0_0_48;
   wire n_0_0_49;
   wire n_0_0_50;
   wire n_0_0_51;
   wire n_0_0_52;
   wire n_0_0_53;
   wire n_0_0_54;
   wire n_0_0_55;
   wire n_0_0_56;
   wire n_0_0_57;
   wire n_0_0_58;
   wire n_0_0_59;
   wire n_0_0_60;
   wire n_0_0_61;
   wire n_0_0_62;
   wire n_0_0_63;
   wire n_0_0_64;
   wire n_0_0_65;
   wire n_0_0_66;
   wire n_0_0_67;
   wire n_0_0_68;
   wire n_0_0_69;
   wire n_0_0_70;
   wire n_0_0_71;
   wire n_0_0_72;
   wire n_0_1018;
   wire n_0_1019;
   wire n_0_1020;
   wire n_0_1021;
   wire n_0_1022;
   wire n_0_1023;
   wire n_0_1024;
   wire n_0_1025;
   wire n_0_1026;
   wire n_0_1027;
   wire n_0_1028;
   wire n_0_1029;
   wire n_0_1030;
   wire n_0_1031;
   wire n_0_1032;
   wire n_0_1033;
   wire n_0_1034;
   wire n_0_1035;
   wire n_0_1036;
   wire n_0_1037;
   wire n_0_1038;
   wire n_0_1067;
   wire n_0_0_73;
   wire n_0_0_74;
   wire n_0_0_75;
   wire n_0_0_76;
   wire n_0_0_77;
   wire n_0_0_78;
   wire n_0_0_79;
   wire n_0_0_80;
   wire n_0_0_81;
   wire n_0_0_82;
   wire n_0_0_83;
   wire n_0_0_84;
   wire n_0_0_85;
   wire n_0_0_86;
   wire n_0_0_87;
   wire n_0_0_88;
   wire n_0_0_89;
   wire n_0_0_90;
   wire n_0_0_91;
   wire n_0_0_92;
   wire n_0_0_93;
   wire n_0_0_94;
   wire n_0_0_95;
   wire n_0_0_96;
   wire n_0_0_97;
   wire n_0_0_98;
   wire n_0_0_99;
   wire n_0_0_100;
   wire n_0_0_101;
   wire n_0_0_102;
   wire n_0_0_103;
   wire n_0_0_104;
   wire n_0_0_105;
   wire n_0_0_106;
   wire n_0_752;
   wire n_0_753;
   wire n_0_754;
   wire n_0_755;
   wire n_0_756;
   wire n_0_757;
   wire n_0_758;
   wire n_0_759;
   wire n_0_760;
   wire n_0_761;
   wire n_0_762;
   wire n_0_763;
   wire n_0_764;
   wire n_0_765;
   wire n_0_766;
   wire n_0_767;
   wire n_0_768;
   wire n_0_769;
   wire n_0_770;
   wire n_0_771;
   wire n_0_772;
   wire n_0_773;
   wire n_0_60;
   wire n_0_0_107;
   wire n_0_0_108;
   wire n_0_0_109;
   wire n_0_0_110;
   wire n_0_0_111;
   wire n_0_0_112;
   wire n_0_0_113;
   wire n_0_0_114;
   wire n_0_0_115;
   wire n_0_0_116;
   wire n_0_0_117;
   wire n_0_0_118;
   wire n_0_0_119;
   wire n_0_0_120;
   wire n_0_0_121;
   wire n_0_0_122;
   wire n_0_0_123;
   wire n_0_0_124;
   wire n_0_0_125;
   wire n_0_0_126;
   wire n_0_0_127;
   wire n_0_0_128;
   wire n_0_0_129;
   wire n_0_0_130;
   wire n_0_0_131;
   wire n_0_0_132;
   wire n_0_0_133;
   wire n_0_0_134;
   wire n_0_0_135;
   wire n_0_0_136;
   wire n_0_0_137;
   wire n_0_0_138;
   wire n_0_707;
   wire n_0_708;
   wire n_0_709;
   wire n_0_710;
   wire n_0_711;
   wire n_0_712;
   wire n_0_713;
   wire n_0_714;
   wire n_0_715;
   wire n_0_716;
   wire n_0_717;
   wire n_0_718;
   wire n_0_719;
   wire n_0_720;
   wire n_0_721;
   wire n_0_722;
   wire n_0_723;
   wire n_0_724;
   wire n_0_725;
   wire n_0_726;
   wire n_0_727;
   wire n_0_728;
   wire n_0_61;
   wire n_0_0_139;
   wire n_0_0_140;
   wire n_0_0_141;
   wire n_0_0_142;
   wire n_0_0_143;
   wire n_0_0_144;
   wire n_0_0_145;
   wire n_0_0_146;
   wire n_0_0_147;
   wire n_0_0_148;
   wire n_0_0_149;
   wire n_0_0_150;
   wire n_0_0_151;
   wire n_0_0_152;
   wire n_0_0_153;
   wire n_0_0_154;
   wire n_0_0_155;
   wire n_0_0_156;
   wire n_0_0_157;
   wire n_0_0_158;
   wire n_0_0_159;
   wire n_0_0_160;
   wire n_0_0_161;
   wire n_0_0_162;
   wire n_0_0_163;
   wire n_0_0_164;
   wire n_0_0_165;
   wire n_0_0_166;
   wire n_0_0_167;
   wire n_0_0_168;
   wire n_0_0_169;
   wire n_0_0_170;
   wire n_0_0_171;
   wire n_0_0_172;
   wire n_0_662;
   wire n_0_663;
   wire n_0_664;
   wire n_0_665;
   wire n_0_666;
   wire n_0_667;
   wire n_0_668;
   wire n_0_669;
   wire n_0_670;
   wire n_0_671;
   wire n_0_672;
   wire n_0_673;
   wire n_0_674;
   wire n_0_675;
   wire n_0_676;
   wire n_0_677;
   wire n_0_678;
   wire n_0_679;
   wire n_0_680;
   wire n_0_681;
   wire n_0_682;
   wire n_0_683;
   wire n_0_62;
   wire n_0_0_173;
   wire n_0_0_174;
   wire n_0_0_175;
   wire n_0_0_176;
   wire n_0_0_177;
   wire n_0_0_178;
   wire n_0_0_179;
   wire n_0_0_180;
   wire n_0_0_181;
   wire n_0_0_182;
   wire n_0_0_183;
   wire n_0_0_184;
   wire n_0_0_185;
   wire n_0_0_186;
   wire n_0_0_187;
   wire n_0_0_188;
   wire n_0_0_189;
   wire n_0_0_190;
   wire n_0_0_191;
   wire n_0_0_192;
   wire n_0_0_193;
   wire n_0_0_194;
   wire n_0_0_195;
   wire n_0_0_196;
   wire n_0_0_197;
   wire n_0_0_198;
   wire n_0_0_199;
   wire n_0_0_200;
   wire n_0_0_201;
   wire n_0_0_202;
   wire n_0_0_203;
   wire n_0_0_204;
   wire n_0_0_205;
   wire n_0_617;
   wire n_0_618;
   wire n_0_619;
   wire n_0_620;
   wire n_0_621;
   wire n_0_622;
   wire n_0_623;
   wire n_0_624;
   wire n_0_625;
   wire n_0_626;
   wire n_0_627;
   wire n_0_628;
   wire n_0_629;
   wire n_0_630;
   wire n_0_631;
   wire n_0_632;
   wire n_0_633;
   wire n_0_634;
   wire n_0_635;
   wire n_0_636;
   wire n_0_637;
   wire n_0_638;
   wire n_0_63;
   wire n_0_0_206;
   wire n_0_0_207;
   wire n_0_0_208;
   wire n_0_0_209;
   wire n_0_0_210;
   wire n_0_0_211;
   wire n_0_0_212;
   wire n_0_0_213;
   wire n_0_0_214;
   wire n_0_0_215;
   wire n_0_0_216;
   wire n_0_0_217;
   wire n_0_0_218;
   wire n_0_0_219;
   wire n_0_0_220;
   wire n_0_0_221;
   wire n_0_0_222;
   wire n_0_0_223;
   wire n_0_0_224;
   wire n_0_0_225;
   wire n_0_0_226;
   wire n_0_0_227;
   wire n_0_0_228;
   wire n_0_0_229;
   wire n_0_0_230;
   wire n_0_0_231;
   wire n_0_0_232;
   wire n_0_0_233;
   wire n_0_0_234;
   wire n_0_0_235;
   wire n_0_0_236;
   wire n_0_0_237;
   wire n_0_572;
   wire n_0_573;
   wire n_0_574;
   wire n_0_575;
   wire n_0_576;
   wire n_0_577;
   wire n_0_578;
   wire n_0_579;
   wire n_0_580;
   wire n_0_581;
   wire n_0_582;
   wire n_0_583;
   wire n_0_584;
   wire n_0_585;
   wire n_0_586;
   wire n_0_587;
   wire n_0_588;
   wire n_0_589;
   wire n_0_590;
   wire n_0_591;
   wire n_0_592;
   wire n_0_593;
   wire n_0_0_238;
   wire n_0_64;
   wire n_0_0_239;
   wire n_0_0_240;
   wire n_0_0_241;
   wire n_0_0_242;
   wire n_0_0_243;
   wire n_0_0_244;
   wire n_0_0_245;
   wire n_0_0_246;
   wire n_0_0_247;
   wire n_0_0_248;
   wire n_0_0_249;
   wire n_0_0_250;
   wire n_0_0_251;
   wire n_0_0_252;
   wire n_0_0_253;
   wire n_0_0_254;
   wire n_0_0_255;
   wire n_0_0_256;
   wire n_0_0_257;
   wire n_0_0_258;
   wire n_0_0_259;
   wire n_0_0_260;
   wire n_0_0_261;
   wire n_0_0_262;
   wire n_0_0_263;
   wire n_0_0_264;
   wire n_0_0_265;
   wire n_0_0_266;
   wire n_0_0_267;
   wire n_0_0_268;
   wire n_0_0_269;
   wire n_0_527;
   wire n_0_528;
   wire n_0_529;
   wire n_0_530;
   wire n_0_531;
   wire n_0_532;
   wire n_0_533;
   wire n_0_534;
   wire n_0_535;
   wire n_0_536;
   wire n_0_537;
   wire n_0_538;
   wire n_0_539;
   wire n_0_540;
   wire n_0_541;
   wire n_0_542;
   wire n_0_543;
   wire n_0_544;
   wire n_0_545;
   wire n_0_546;
   wire n_0_547;
   wire n_0_548;
   wire n_0_65;
   wire n_0_0_270;
   wire n_0_0_271;
   wire n_0_0_272;
   wire n_0_0_273;
   wire n_0_0_274;
   wire n_0_0_275;
   wire n_0_0_276;
   wire n_0_0_277;
   wire n_0_0_278;
   wire n_0_0_279;
   wire n_0_0_280;
   wire n_0_0_281;
   wire n_0_0_282;
   wire n_0_0_283;
   wire n_0_0_284;
   wire n_0_0_285;
   wire n_0_0_286;
   wire n_0_0_287;
   wire n_0_0_288;
   wire n_0_0_289;
   wire n_0_0_290;
   wire n_0_0_291;
   wire n_0_0_292;
   wire n_0_0_293;
   wire n_0_0_294;
   wire n_0_0_295;
   wire n_0_0_296;
   wire n_0_0_297;
   wire n_0_0_298;
   wire n_0_0_299;
   wire n_0_0_300;
   wire n_0_0_301;
   wire n_0_0_302;
   wire n_0_482;
   wire n_0_483;
   wire n_0_484;
   wire n_0_485;
   wire n_0_486;
   wire n_0_487;
   wire n_0_488;
   wire n_0_489;
   wire n_0_490;
   wire n_0_491;
   wire n_0_492;
   wire n_0_493;
   wire n_0_494;
   wire n_0_495;
   wire n_0_496;
   wire n_0_497;
   wire n_0_498;
   wire n_0_499;
   wire n_0_500;
   wire n_0_501;
   wire n_0_502;
   wire n_0_503;
   wire n_0_66;
   wire n_0_0_303;
   wire n_0_0_304;
   wire n_0_0_305;
   wire n_0_0_306;
   wire n_0_0_307;
   wire n_0_0_308;
   wire n_0_0_309;
   wire n_0_0_310;
   wire n_0_0_311;
   wire n_0_0_312;
   wire n_0_0_313;
   wire n_0_0_314;
   wire n_0_0_315;
   wire n_0_0_316;
   wire n_0_0_317;
   wire n_0_0_318;
   wire n_0_0_319;
   wire n_0_0_320;
   wire n_0_0_321;
   wire n_0_0_322;
   wire n_0_0_323;
   wire n_0_0_324;
   wire n_0_0_325;
   wire n_0_0_326;
   wire n_0_0_327;
   wire n_0_0_328;
   wire n_0_0_329;
   wire n_0_0_330;
   wire n_0_0_331;
   wire n_0_0_332;
   wire n_0_0_333;
   wire n_0_0_334;
   wire n_0_0_335;
   wire n_0_437;
   wire n_0_438;
   wire n_0_439;
   wire n_0_440;
   wire n_0_441;
   wire n_0_442;
   wire n_0_443;
   wire n_0_444;
   wire n_0_445;
   wire n_0_446;
   wire n_0_447;
   wire n_0_448;
   wire n_0_449;
   wire n_0_450;
   wire n_0_451;
   wire n_0_452;
   wire n_0_453;
   wire n_0_454;
   wire n_0_455;
   wire n_0_456;
   wire n_0_457;
   wire n_0_458;
   wire n_0_67;
   wire n_0_0_336;
   wire n_0_0_337;
   wire n_0_0_338;
   wire n_0_0_339;
   wire n_0_0_340;
   wire n_0_0_341;
   wire n_0_0_342;
   wire n_0_0_343;
   wire n_0_0_344;
   wire n_0_0_345;
   wire n_0_0_346;
   wire n_0_0_347;
   wire n_0_0_348;
   wire n_0_0_349;
   wire n_0_0_350;
   wire n_0_0_351;
   wire n_0_0_352;
   wire n_0_0_353;
   wire n_0_0_354;
   wire n_0_0_355;
   wire n_0_0_356;
   wire n_0_0_357;
   wire n_0_0_358;
   wire n_0_0_359;
   wire n_0_0_360;
   wire n_0_0_361;
   wire n_0_0_362;
   wire n_0_0_363;
   wire n_0_0_364;
   wire n_0_0_365;
   wire n_0_0_366;
   wire n_0_0_367;
   wire n_0_392;
   wire n_0_393;
   wire n_0_394;
   wire n_0_395;
   wire n_0_396;
   wire n_0_397;
   wire n_0_398;
   wire n_0_399;
   wire n_0_400;
   wire n_0_401;
   wire n_0_402;
   wire n_0_403;
   wire n_0_404;
   wire n_0_405;
   wire n_0_406;
   wire n_0_407;
   wire n_0_408;
   wire n_0_409;
   wire n_0_410;
   wire n_0_411;
   wire n_0_412;
   wire n_0_413;
   wire n_0_68;
   wire n_0_0_368;
   wire n_0_0_369;
   wire n_0_0_370;
   wire n_0_0_371;
   wire n_0_0_372;
   wire n_0_0_373;
   wire n_0_0_374;
   wire n_0_0_375;
   wire n_0_0_376;
   wire n_0_0_377;
   wire n_0_0_378;
   wire n_0_0_379;
   wire n_0_0_380;
   wire n_0_0_381;
   wire n_0_0_382;
   wire n_0_0_383;
   wire n_0_0_384;
   wire n_0_0_385;
   wire n_0_0_386;
   wire n_0_0_387;
   wire n_0_0_388;
   wire n_0_0_389;
   wire n_0_0_390;
   wire n_0_0_391;
   wire n_0_0_392;
   wire n_0_0_393;
   wire n_0_0_394;
   wire n_0_0_395;
   wire n_0_0_396;
   wire n_0_0_397;
   wire n_0_0_398;
   wire n_0_0_399;
   wire n_0_347;
   wire n_0_348;
   wire n_0_349;
   wire n_0_350;
   wire n_0_351;
   wire n_0_352;
   wire n_0_353;
   wire n_0_354;
   wire n_0_355;
   wire n_0_356;
   wire n_0_357;
   wire n_0_358;
   wire n_0_359;
   wire n_0_360;
   wire n_0_361;
   wire n_0_362;
   wire n_0_363;
   wire n_0_364;
   wire n_0_365;
   wire n_0_366;
   wire n_0_367;
   wire n_0_368;
   wire n_0_0_400;
   wire n_0_0_401;
   wire n_0_0_402;
   wire n_0_0_403;
   wire n_0_0_404;
   wire n_0_0_405;
   wire n_0_0_406;
   wire n_0_0_407;
   wire n_0_0_408;
   wire n_0_0_409;
   wire n_0_0_410;
   wire n_0_0_411;
   wire n_0_0_412;
   wire n_0_0_413;
   wire n_0_0_414;
   wire n_0_0_415;
   wire n_0_0_416;
   wire n_0_0_417;
   wire n_0_0_418;
   wire n_0_0_419;
   wire n_0_0_420;
   wire n_0_0_421;
   wire n_0_0_422;
   wire n_0_0_423;
   wire n_0_0_424;
   wire n_0_0_425;
   wire n_0_0_426;
   wire n_0_0_427;
   wire n_0_0_428;
   wire n_0_0_429;
   wire n_0_0_430;
   wire n_0_0_431;
   wire n_0_302;
   wire n_0_303;
   wire n_0_304;
   wire n_0_305;
   wire n_0_306;
   wire n_0_307;
   wire n_0_308;
   wire n_0_309;
   wire n_0_310;
   wire n_0_311;
   wire n_0_312;
   wire n_0_313;
   wire n_0_314;
   wire n_0_315;
   wire n_0_316;
   wire n_0_317;
   wire n_0_318;
   wire n_0_319;
   wire n_0_320;
   wire n_0_321;
   wire n_0_322;
   wire n_0_323;
   wire n_0_0_432;
   wire n_0_0_433;
   wire n_0_0_434;
   wire n_0_0_435;
   wire n_0_0_436;
   wire n_0_0_437;
   wire n_0_0_438;
   wire n_0_0_439;
   wire n_0_0_440;
   wire n_0_0_441;
   wire n_0_0_442;
   wire n_0_0_443;
   wire n_0_0_444;
   wire n_0_0_445;
   wire n_0_0_446;
   wire n_0_0_447;
   wire n_0_0_448;
   wire n_0_0_449;
   wire n_0_0_450;
   wire n_0_0_451;
   wire n_0_0_452;
   wire n_0_0_453;
   wire n_0_0_454;
   wire n_0_0_455;
   wire n_0_0_456;
   wire n_0_0_457;
   wire n_0_0_458;
   wire n_0_0_459;
   wire n_0_0_460;
   wire n_0_0_461;
   wire n_0_0_462;
   wire n_0_0_463;
   wire n_0_257;
   wire n_0_258;
   wire n_0_259;
   wire n_0_260;
   wire n_0_261;
   wire n_0_262;
   wire n_0_263;
   wire n_0_264;
   wire n_0_265;
   wire n_0_266;
   wire n_0_267;
   wire n_0_268;
   wire n_0_269;
   wire n_0_270;
   wire n_0_271;
   wire n_0_272;
   wire n_0_273;
   wire n_0_274;
   wire n_0_275;
   wire n_0_276;
   wire n_0_277;
   wire n_0_278;
   wire n_0_0_464;
   wire n_0_0_465;
   wire n_0_0_466;
   wire n_0_0_467;
   wire n_0_0_468;
   wire n_0_0_469;
   wire n_0_0_470;
   wire n_0_0_471;
   wire n_0_0_472;
   wire n_0_0_473;
   wire n_0_0_474;
   wire n_0_0_475;
   wire n_0_0_476;
   wire n_0_0_477;
   wire n_0_0_478;
   wire n_0_0_479;
   wire n_0_0_480;
   wire n_0_0_481;
   wire n_0_0_482;
   wire n_0_0_483;
   wire n_0_0_484;
   wire n_0_0_485;
   wire n_0_0_486;
   wire n_0_0_487;
   wire n_0_0_488;
   wire n_0_0_489;
   wire n_0_0_490;
   wire n_0_0_491;
   wire n_0_0_492;
   wire n_0_0_493;
   wire n_0_0_494;
   wire n_0_0_495;
   wire n_0_212;
   wire n_0_213;
   wire n_0_214;
   wire n_0_215;
   wire n_0_216;
   wire n_0_217;
   wire n_0_218;
   wire n_0_219;
   wire n_0_220;
   wire n_0_221;
   wire n_0_222;
   wire n_0_223;
   wire n_0_224;
   wire n_0_225;
   wire n_0_226;
   wire n_0_227;
   wire n_0_228;
   wire n_0_229;
   wire n_0_230;
   wire n_0_231;
   wire n_0_232;
   wire n_0_233;
   wire n_0_0_496;
   wire n_0_0_497;
   wire n_0_0_498;
   wire n_0_0_499;
   wire n_0_0_500;
   wire n_0_0_501;
   wire n_0_0_502;
   wire n_0_0_503;
   wire n_0_0_504;
   wire n_0_0_505;
   wire n_0_0_506;
   wire n_0_0_507;
   wire n_0_0_508;
   wire n_0_0_509;
   wire n_0_0_510;
   wire n_0_0_511;
   wire n_0_0_512;
   wire n_0_0_513;
   wire n_0_0_514;
   wire n_0_0_515;
   wire n_0_0_516;
   wire n_0_0_517;
   wire n_0_0_518;
   wire n_0_0_519;
   wire n_0_0_520;
   wire n_0_0_521;
   wire n_0_0_522;
   wire n_0_0_523;
   wire n_0_0_524;
   wire n_0_0_525;
   wire n_0_0_526;
   wire n_0_0_527;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_180;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_0_528;
   wire n_0_0_529;
   wire n_0_0_530;
   wire n_0_0_531;
   wire n_0_0_532;
   wire n_0_0_533;
   wire n_0_0_534;
   wire n_0_0_535;
   wire n_0_0_536;
   wire n_0_0_537;
   wire n_0_0_538;
   wire n_0_0_539;
   wire n_0_0_540;
   wire n_0_0_541;
   wire n_0_0_542;
   wire n_0_0_543;
   wire n_0_0_544;
   wire n_0_0_545;
   wire n_0_0_546;
   wire n_0_0_547;
   wire n_0_0_548;
   wire n_0_0_549;
   wire n_0_0_550;
   wire n_0_0_551;
   wire n_0_0_552;
   wire n_0_0_553;
   wire n_0_0_554;
   wire n_0_0_555;
   wire n_0_0_556;
   wire n_0_0_557;
   wire n_0_0_558;
   wire n_0_0_559;
   wire n_0_0_560;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_0_561;
   wire n_0_0_562;
   wire n_0_0_563;
   wire n_0_0_564;
   wire n_0_0_565;
   wire n_0_0_566;
   wire n_0_0_567;
   wire n_0_0_568;
   wire n_0_0_569;
   wire n_0_0_570;
   wire n_0_0_571;
   wire n_0_0_572;
   wire n_0_0_573;
   wire n_0_0_574;
   wire n_0_0_575;
   wire n_0_0_576;
   wire n_0_0_577;
   wire n_0_0_578;
   wire n_0_0_579;
   wire n_0_0_580;
   wire n_0_0_581;
   wire n_0_0_582;
   wire n_0_0_583;
   wire n_0_0_584;
   wire n_0_0_585;
   wire n_0_0_586;
   wire n_0_0_587;
   wire n_0_0_588;
   wire n_0_0_589;
   wire n_0_0_590;
   wire n_0_0_591;
   wire n_0_0_592;
   wire n_0_0_593;
   wire n_0_0_594;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_0_595;
   wire n_0_0_596;
   wire n_0_0_597;
   wire n_0_0_598;
   wire n_0_0_599;
   wire n_0_0_600;
   wire n_0_0_601;
   wire n_0_0_602;
   wire n_0_0_603;
   wire n_0_0_604;
   wire n_0_973;
   wire n_0_974;
   wire n_0_975;
   wire n_0_976;
   wire n_0_977;
   wire n_0_978;
   wire n_0_979;
   wire n_0_980;
   wire n_0_981;
   wire n_0_982;
   wire n_0_983;
   wire n_0_984;
   wire n_0_985;
   wire n_0_986;
   wire n_0_987;
   wire n_0_988;
   wire n_0_989;
   wire n_0_990;
   wire n_0_991;
   wire n_0_992;
   wire n_0_993;
   wire n_0_994;
   wire n_0_1068;
   wire n_0_0_605;
   wire n_0_0_606;
   wire n_0_0_607;
   wire n_0_0_608;
   wire n_0_0_609;
   wire n_0_0_610;
   wire n_0_0_611;
   wire n_0_0_612;
   wire n_0_0_613;
   wire n_0_0_614;
   wire n_0_0_615;
   wire n_0_0_616;
   wire n_0_0_617;
   wire n_0_0_618;
   wire n_0_0_619;
   wire n_0_0_620;
   wire n_0_0_621;
   wire n_0_0_622;
   wire n_0_0_623;
   wire n_0_0_624;
   wire n_0_0_625;
   wire n_0_0_626;
   wire n_0_0_627;
   wire n_0_0_628;
   wire n_0_0_629;
   wire n_0_0_630;
   wire n_0_0_631;
   wire n_0_0_632;
   wire n_0_0_633;
   wire n_0_0_634;
   wire n_0_0_635;
   wire n_0_0_636;
   wire n_0_929;
   wire n_0_930;
   wire n_0_931;
   wire n_0_932;
   wire n_0_933;
   wire n_0_934;
   wire n_0_935;
   wire n_0_936;
   wire n_0_937;
   wire n_0_938;
   wire n_0_939;
   wire n_0_940;
   wire n_0_941;
   wire n_0_942;
   wire n_0_943;
   wire n_0_944;
   wire n_0_945;
   wire n_0_946;
   wire n_0_947;
   wire n_0_948;
   wire n_0_949;
   wire n_0_950;
   wire n_0_1069;
   wire n_0_0_637;
   wire n_0_0_638;
   wire n_0_0_639;
   wire n_0_0_640;
   wire n_0_0_641;
   wire n_0_0_642;
   wire n_0_0_643;
   wire n_0_0_644;
   wire n_0_0_645;
   wire n_0_0_646;
   wire n_0_0_647;
   wire n_0_0_648;
   wire n_0_0_649;
   wire n_0_0_650;
   wire n_0_0_651;
   wire n_0_0_652;
   wire n_0_0_653;
   wire n_0_0_654;
   wire n_0_0_655;
   wire n_0_0_656;
   wire n_0_0_657;
   wire n_0_0_658;
   wire n_0_0_659;
   wire n_0_0_660;
   wire n_0_0_661;
   wire n_0_0_662;
   wire n_0_0_663;
   wire n_0_0_664;
   wire n_0_0_665;
   wire n_0_885;
   wire n_0_886;
   wire n_0_887;
   wire n_0_888;
   wire n_0_889;
   wire n_0_890;
   wire n_0_891;
   wire n_0_892;
   wire n_0_893;
   wire n_0_894;
   wire n_0_895;
   wire n_0_896;
   wire n_0_897;
   wire n_0_898;
   wire n_0_899;
   wire n_0_900;
   wire n_0_901;
   wire n_0_902;
   wire n_0_903;
   wire n_0_904;
   wire n_0_905;
   wire n_0_906;
   wire n_0_0_666;
   wire n_0_1070;
   wire n_0_0_667;
   wire n_0_0_668;
   wire n_0_0_669;
   wire n_0_0_670;
   wire n_0_0_671;
   wire n_0_0_672;
   wire n_0_0_673;
   wire n_0_0_674;
   wire n_0_0_675;
   wire n_0_0_676;
   wire n_0_0_677;
   wire n_0_0_678;
   wire n_0_0_679;
   wire n_0_0_680;
   wire n_0_0_681;
   wire n_0_0_682;
   wire n_0_0_683;
   wire n_0_0_684;
   wire n_0_0_685;
   wire n_0_0_686;
   wire n_0_0_687;
   wire n_0_0_688;
   wire n_0_0_689;
   wire n_0_0_690;
   wire n_0_0_691;
   wire n_0_0_692;
   wire n_0_0_693;
   wire n_0_0_694;
   wire n_0_0_695;
   wire n_0_841;
   wire n_0_842;
   wire n_0_843;
   wire n_0_844;
   wire n_0_845;
   wire n_0_846;
   wire n_0_847;
   wire n_0_848;
   wire n_0_849;
   wire n_0_850;
   wire n_0_851;
   wire n_0_852;
   wire n_0_853;
   wire n_0_854;
   wire n_0_855;
   wire n_0_856;
   wire n_0_857;
   wire n_0_858;
   wire n_0_859;
   wire n_0_860;
   wire n_0_861;
   wire n_0_862;
   wire n_0_0_696;
   wire n_0_1071;
   wire n_0_0_697;
   wire n_0_0_698;
   wire n_0_0_699;
   wire n_0_0_700;
   wire n_0_0_701;
   wire n_0_0_702;
   wire n_0_0_703;
   wire n_0_0_704;
   wire n_0_0_705;
   wire n_0_0_706;
   wire n_0_0_707;
   wire n_0_0_708;
   wire n_0_0_709;
   wire n_0_0_710;
   wire n_0_0_711;
   wire n_0_0_712;
   wire n_0_0_713;
   wire n_0_0_714;
   wire n_0_0_715;
   wire n_0_0_716;
   wire n_0_0_717;
   wire n_0_0_718;
   wire n_0_0_719;
   wire n_0_0_720;
   wire n_0_0_721;
   wire n_0_0_722;
   wire n_0_0_723;
   wire n_0_0_724;
   wire n_0_0_725;
   wire n_0_797;
   wire n_0_798;
   wire n_0_799;
   wire n_0_800;
   wire n_0_801;
   wire n_0_802;
   wire n_0_803;
   wire n_0_804;
   wire n_0_805;
   wire n_0_806;
   wire n_0_807;
   wire n_0_808;
   wire n_0_809;
   wire n_0_810;
   wire n_0_811;
   wire n_0_812;
   wire n_0_813;
   wire n_0_814;
   wire n_0_815;
   wire n_0_816;
   wire n_0_817;
   wire n_0_818;
   wire n_0_1072;
   wire n_0_0_726;
   wire n_0_0_727;
   wire n_0_0_728;
   wire n_0_0_729;
   wire n_0_0_730;
   wire n_0_0_731;
   wire n_0_0_732;
   wire n_0_0_733;
   wire n_0_0_734;
   wire n_0_0_735;
   wire n_0_0_736;
   wire n_0_0_737;
   wire n_0_0_738;
   wire n_0_0_739;
   wire n_0_0_740;
   wire n_0_0_741;
   wire n_0_0_742;
   wire n_0_0_743;
   wire n_0_0_744;
   wire n_0_0_745;
   wire n_0_0_746;
   wire n_0_0_747;
   wire n_0_0_748;
   wire n_0_0_749;
   wire n_0_0_750;
   wire n_0_0_751;
   wire n_0_0_752;
   wire n_0_0_753;
   wire n_0_0_754;
   wire n_0_0_755;
   wire n_0_0_756;
   wire n_0_0_757;
   wire n_0_0_758;
   wire n_0_0_759;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_0_760;
   wire n_0_74;
   wire n_0_0_761;
   wire n_0_0_762;
   wire n_0_75;
   wire n_0_76;
   wire n_0_0_763;
   wire n_0_77;
   wire n_0_121;
   wire n_0_166;
   wire n_0_211;
   wire n_0_256;
   wire n_0_0_764;
   wire n_0_301;
   wire n_0_0_765;
   wire n_0_0_766;
   wire n_0_346;
   wire n_0_0_767;
   wire n_0_0_768;
   wire n_0_0_769;
   wire n_0_0_770;
   wire n_0_0_771;
   wire n_0_0_772;
   wire n_0_0_773;
   wire n_0_0_774;
   wire n_0_0_775;
   wire n_0_0_776;
   wire n_0_0_777;
   wire n_0_0_778;
   wire n_0_0_779;
   wire n_0_0_780;
   wire n_0_0_781;
   wire n_0_0_782;
   wire n_0_0_783;
   wire n_0_0_784;
   wire n_0_0_785;
   wire n_0_0_786;
   wire n_0_0_787;
   wire n_0_0_788;
   wire n_0_0_789;
   wire n_0_0_790;
   wire n_0_391;
   wire n_0_0_791;
   wire n_0_0_792;
   wire n_0_436;
   wire n_0_0_793;
   wire n_0_0_794;
   wire n_0_481;
   wire n_0_0_795;
   wire n_0_0_796;
   wire n_0_526;
   wire n_0_0_797;
   wire n_0_0_798;
   wire n_0_571;
   wire n_0_0_799;
   wire n_0_0_800;
   wire n_0_616;
   wire n_0_0_801;
   wire n_0_0_802;
   wire n_0_661;
   wire n_0_0_803;
   wire n_0_0_804;
   wire n_0_706;
   wire n_0_0_805;
   wire n_0_0_806;
   wire n_0_751;
   wire n_0_0_807;
   wire n_0_0_808;
   wire n_0_796;
   wire n_0_0_809;
   wire n_0_0_810;
   wire n_0_840;
   wire n_0_0_811;
   wire n_0_0_812;
   wire n_0_884;
   wire n_0_0_813;
   wire n_0_0_814;
   wire n_0_928;
   wire n_0_0_815;
   wire n_0_0_816;
   wire n_0_972;
   wire n_0_0_817;
   wire n_0_0_818;
   wire n_0_1016;
   wire n_0_0_819;
   wire n_0_0_820;
   wire n_0_1017;
   wire n_0_0_821;
   wire n_0_0_822;
   wire n_0_1060;
   wire n_0_0_823;
   wire n_0_0_824;
   wire n_0_1061;
   wire n_0_0_825;
   wire n_0_0_826;
   wire n_0_1062;
   wire n_0_0_827;
   wire n_0_0_828;
   wire n_0_1063;
   wire n_0_0_829;
   wire n_0_0_830;
   wire n_0_1064;
   wire n_0_0_831;
   wire n_0_0_832;
   wire n_0_39;
   wire n_0_0_833;
   wire n_0_0_834;
   wire n_0_0_835;
   wire n_0_0_836;
   wire n_0_0_837;
   wire n_0_0_838;
   wire n_0_0_839;
   wire n_0_0_840;
   wire n_0_0_841;
   wire n_0_0_842;
   wire n_0_0_843;
   wire n_0_0_844;
   wire n_0_0_845;
   wire n_0_0_846;
   wire n_0_0_847;
   wire n_0_0_848;
   wire n_0_0_849;
   wire n_0_0_850;
   wire n_0_0_851;
   wire n_0_0_852;
   wire n_0_0_853;
   wire n_0_0_854;
   wire n_0_0_855;
   wire n_0_0_856;
   wire n_0_0_857;
   wire n_0_0_858;
   wire n_0_0_859;
   wire n_0_0_860;
   wire n_0_0_861;
   wire n_0_0_862;

   assign out_c[63] = out_c[16];
   assign out_c[62] = out_c[16];
   assign out_c[61] = out_c[16];
   assign out_c[60] = out_c[16];
   assign out_c[59] = out_c[16];
   assign out_c[58] = out_c[16];
   assign out_c[57] = out_c[16];
   assign out_c[56] = out_c[16];
   assign out_c[55] = out_c[16];
   assign out_c[54] = out_c[16];
   assign out_c[53] = out_c[16];
   assign out_c[52] = out_c[16];
   assign out_c[51] = out_c[16];
   assign out_c[50] = out_c[16];
   assign out_c[49] = out_c[16];
   assign out_c[48] = out_c[16];
   assign out_c[47] = out_c[16];
   assign out_c[46] = out_c[16];
   assign out_c[45] = out_c[16];
   assign out_c[44] = out_c[16];
   assign out_c[43] = out_c[16];
   assign out_c[42] = out_c[16];
   assign out_c[41] = out_c[16];
   assign out_c[40] = out_c[16];
   assign out_c[39] = out_c[16];
   assign out_c[38] = out_c[16];
   assign out_c[37] = out_c[16];
   assign out_c[36] = out_c[16];
   assign out_c[35] = out_c[16];
   assign out_c[34] = out_c[16];
   assign out_c[33] = out_c[16];
   assign out_c[32] = out_c[16];
   assign out_c[31] = out_c[16];
   assign out_c[30] = out_c[16];
   assign out_c[29] = out_c[16];
   assign out_c[28] = out_c[16];
   assign out_c[27] = out_c[16];
   assign out_c[26] = out_c[16];
   assign out_c[25] = out_c[16];
   assign out_c[24] = out_c[16];
   assign out_c[23] = out_c[16];
   assign out_c[22] = out_c[16];
   assign out_c[21] = out_c[16];
   assign out_c[20] = out_c[16];
   assign out_c[19] = out_c[16];
   assign out_c[18] = out_c[16];
   assign out_c[17] = out_c[16];

   DFFR_X1 posv_flag_reg (.D(n_0_42), .RN(n_0_39), .CK(n_0_38), .Q(posv), .QN());
   datapath i_0_1 (.in_b({in_b[22], in_b[21], in_b[20], in_b[19], in_b[18], 
      in_b[17], in_b[16], in_b[15], in_b[14], in_b[13], in_b[12], in_b[11], 
      in_b[10], in_b[9], in_b[8], in_b[7], in_b[6], in_b[5], in_b[4], in_b[3], 
      in_b[2], in_b[1], in_b[0]}), .p_0({n_0_22, n_0_21, n_0_20, n_0_19, n_0_18, 
      n_0_17, n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, n_0_11, n_0_10, n_0_9, 
      n_0_8, n_0_7, n_0_6, n_0_5, n_0_4, n_0_3, n_0_2, n_0_1, uc_0}));
   datapath__0_7 i_0_9 (.p_0({uc_1, n_0_1064, n_0_1063, n_0_1062, n_0_1061, 
      n_0_1060, n_0_1017, n_0_1016, n_0_972, n_0_928, n_0_884, n_0_840, n_0_796, 
      n_0_751, n_0_706, n_0_661, n_0_616, n_0_571, n_0_526, n_0_481, n_0_436, 
      n_0_391, in_b[0]}), .p_1({uc_2, n_0_98, n_0_97, n_0_96, n_0_95, n_0_94, 
      n_0_93, n_0_92, n_0_91, n_0_90, n_0_89, n_0_88, n_0_87, n_0_86, n_0_85, 
      n_0_84, n_0_83, n_0_82, n_0_81, n_0_80, n_0_79, n_0_78, uc_3}));
   datapath__0_9 i_0_11 (.p_0({uc_4, n_0_120, n_0_119, n_0_118, n_0_117, n_0_116, 
      n_0_115, n_0_114, n_0_113, n_0_112, n_0_111, n_0_110, n_0_109, n_0_108, 
      n_0_107, n_0_106, n_0_105, n_0_104, n_0_103, n_0_102, n_0_101, n_0_100, 
      n_0_99}), .p_1({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      n_0_346}), .divider({uc_5, divider[21], divider[20], divider[19], 
      divider[18], divider[17], divider[16], divider[15], divider[14], 
      divider[13], divider[12], divider[11], divider[10], divider[9], divider[8], 
      divider[7], divider[6], divider[5], divider[4], divider[3], divider[2], 
      divider[1], divider[0]}));
   datapath__0_13 i_0_14 (.p_0({uc_6, n_0_143, n_0_142, n_0_141, n_0_140, 
      n_0_139, n_0_138, n_0_137, n_0_136, n_0_135, n_0_134, n_0_133, n_0_132, 
      n_0_131, n_0_130, n_0_129, n_0_128, n_0_127, n_0_126, n_0_125, n_0_124, 
      n_0_123, n_0_122}), .p_1({uc_7, divider[20], divider[19], divider[18], 
      divider[17], divider[16], divider[15], divider[14], divider[13], 
      divider[12], divider[11], divider[10], divider[9], divider[8], divider[7], 
      divider[6], divider[5], divider[4], divider[3], divider[2], divider[1], 
      divider[0], n_0_301}), .divider({uc_8, n_0_165, n_0_164, n_0_163, n_0_162, 
      n_0_161, n_0_160, n_0_159, n_0_158, n_0_157, n_0_156, n_0_155, n_0_154, 
      n_0_153, n_0_152, n_0_151, n_0_150, n_0_149, n_0_148, n_0_147, n_0_146, 
      n_0_145, n_0_144}));
   datapath__0_17 i_0_17 (.p_0({uc_9, n_0_188, n_0_187, n_0_186, n_0_185, 
      n_0_184, n_0_183, n_0_182, n_0_181, n_0_180, n_0_179, n_0_178, n_0_177, 
      n_0_176, n_0_175, n_0_174, n_0_173, n_0_172, n_0_171, n_0_170, n_0_169, 
      n_0_168, n_0_167}), .p_1({uc_10, n_0_164, n_0_163, n_0_162, n_0_161, 
      n_0_160, n_0_159, n_0_158, n_0_157, n_0_156, n_0_155, n_0_154, n_0_153, 
      n_0_152, n_0_151, n_0_150, n_0_149, n_0_148, n_0_147, n_0_146, n_0_145, 
      n_0_144, n_0_256}), .divider({uc_11, n_0_210, n_0_209, n_0_208, n_0_207, 
      n_0_206, n_0_205, n_0_204, n_0_203, n_0_202, n_0_201, n_0_200, n_0_199, 
      n_0_198, n_0_197, n_0_196, n_0_195, n_0_194, n_0_193, n_0_192, n_0_191, 
      n_0_190, n_0_189}));
   datapath__0_21 i_0_20 (.p_0({uc_12, n_0_233, n_0_232, n_0_231, n_0_230, 
      n_0_229, n_0_228, n_0_227, n_0_226, n_0_225, n_0_224, n_0_223, n_0_222, 
      n_0_221, n_0_220, n_0_219, n_0_218, n_0_217, n_0_216, n_0_215, n_0_214, 
      n_0_213, n_0_212}), .p_1({uc_13, n_0_209, n_0_208, n_0_207, n_0_206, 
      n_0_205, n_0_204, n_0_203, n_0_202, n_0_201, n_0_200, n_0_199, n_0_198, 
      n_0_197, n_0_196, n_0_195, n_0_194, n_0_193, n_0_192, n_0_191, n_0_190, 
      n_0_189, n_0_211}), .divider({uc_14, n_0_255, n_0_254, n_0_253, n_0_252, 
      n_0_251, n_0_250, n_0_249, n_0_248, n_0_247, n_0_246, n_0_245, n_0_244, 
      n_0_243, n_0_242, n_0_241, n_0_240, n_0_239, n_0_238, n_0_237, n_0_236, 
      n_0_235, n_0_234}));
   datapath__0_25 i_0_23 (.p_0({uc_15, n_0_278, n_0_277, n_0_276, n_0_275, 
      n_0_274, n_0_273, n_0_272, n_0_271, n_0_270, n_0_269, n_0_268, n_0_267, 
      n_0_266, n_0_265, n_0_264, n_0_263, n_0_262, n_0_261, n_0_260, n_0_259, 
      n_0_258, n_0_257}), .p_1({uc_16, n_0_254, n_0_253, n_0_252, n_0_251, 
      n_0_250, n_0_249, n_0_248, n_0_247, n_0_246, n_0_245, n_0_244, n_0_243, 
      n_0_242, n_0_241, n_0_240, n_0_239, n_0_238, n_0_237, n_0_236, n_0_235, 
      n_0_234, n_0_166}), .divider({uc_17, n_0_300, n_0_299, n_0_298, n_0_297, 
      n_0_296, n_0_295, n_0_294, n_0_293, n_0_292, n_0_291, n_0_290, n_0_289, 
      n_0_288, n_0_287, n_0_286, n_0_285, n_0_284, n_0_283, n_0_282, n_0_281, 
      n_0_280, n_0_279}));
   datapath__0_29 i_0_26 (.p_0({uc_18, n_0_323, n_0_322, n_0_321, n_0_320, 
      n_0_319, n_0_318, n_0_317, n_0_316, n_0_315, n_0_314, n_0_313, n_0_312, 
      n_0_311, n_0_310, n_0_309, n_0_308, n_0_307, n_0_306, n_0_305, n_0_304, 
      n_0_303, n_0_302}), .p_1({uc_19, n_0_299, n_0_298, n_0_297, n_0_296, 
      n_0_295, n_0_294, n_0_293, n_0_292, n_0_291, n_0_290, n_0_289, n_0_288, 
      n_0_287, n_0_286, n_0_285, n_0_284, n_0_283, n_0_282, n_0_281, n_0_280, 
      n_0_279, n_0_121}), .divider({uc_20, n_0_345, n_0_344, n_0_343, n_0_342, 
      n_0_341, n_0_340, n_0_339, n_0_338, n_0_337, n_0_336, n_0_335, n_0_334, 
      n_0_333, n_0_332, n_0_331, n_0_330, n_0_329, n_0_328, n_0_327, n_0_326, 
      n_0_325, n_0_324}));
   datapath__0_33 i_0_29 (.p_0({uc_21, n_0_368, n_0_367, n_0_366, n_0_365, 
      n_0_364, n_0_363, n_0_362, n_0_361, n_0_360, n_0_359, n_0_358, n_0_357, 
      n_0_356, n_0_355, n_0_354, n_0_353, n_0_352, n_0_351, n_0_350, n_0_349, 
      n_0_348, n_0_347}), .p_1({uc_22, n_0_344, n_0_343, n_0_342, n_0_341, 
      n_0_340, n_0_339, n_0_338, n_0_337, n_0_336, n_0_335, n_0_334, n_0_333, 
      n_0_332, n_0_331, n_0_330, n_0_329, n_0_328, n_0_327, n_0_326, n_0_325, 
      n_0_324, n_0_77}), .divider({uc_23, n_0_390, n_0_389, n_0_388, n_0_387, 
      n_0_386, n_0_385, n_0_384, n_0_383, n_0_382, n_0_381, n_0_380, n_0_379, 
      n_0_378, n_0_377, n_0_376, n_0_375, n_0_374, n_0_373, n_0_372, n_0_371, 
      n_0_370, n_0_369}));
   datapath__0_37 i_0_32 (.p_0({uc_24, n_0_413, n_0_412, n_0_411, n_0_410, 
      n_0_409, n_0_408, n_0_407, n_0_406, n_0_405, n_0_404, n_0_403, n_0_402, 
      n_0_401, n_0_400, n_0_399, n_0_398, n_0_397, n_0_396, n_0_395, n_0_394, 
      n_0_393, n_0_392}), .p_1({uc_25, n_0_389, n_0_388, n_0_387, n_0_386, 
      n_0_385, n_0_384, n_0_383, n_0_382, n_0_381, n_0_380, n_0_379, n_0_378, 
      n_0_377, n_0_376, n_0_375, n_0_374, n_0_373, n_0_372, n_0_371, n_0_370, 
      n_0_369, n_0_76}), .divider({uc_26, n_0_435, n_0_434, n_0_433, n_0_432, 
      n_0_431, n_0_430, n_0_429, n_0_428, n_0_427, n_0_426, n_0_425, n_0_424, 
      n_0_423, n_0_422, n_0_421, n_0_420, n_0_419, n_0_418, n_0_417, n_0_416, 
      n_0_415, n_0_414}));
   datapath__0_41 i_0_35 (.p_0({uc_27, n_0_458, n_0_457, n_0_456, n_0_455, 
      n_0_454, n_0_453, n_0_452, n_0_451, n_0_450, n_0_449, n_0_448, n_0_447, 
      n_0_446, n_0_445, n_0_444, n_0_443, n_0_442, n_0_441, n_0_440, n_0_439, 
      n_0_438, n_0_437}), .p_1({uc_28, n_0_434, n_0_433, n_0_432, n_0_431, 
      n_0_430, n_0_429, n_0_428, n_0_427, n_0_426, n_0_425, n_0_424, n_0_423, 
      n_0_422, n_0_421, n_0_420, n_0_419, n_0_418, n_0_417, n_0_416, n_0_415, 
      n_0_414, n_0_75}), .divider({uc_29, n_0_480, n_0_479, n_0_478, n_0_477, 
      n_0_476, n_0_475, n_0_474, n_0_473, n_0_472, n_0_471, n_0_470, n_0_469, 
      n_0_468, n_0_467, n_0_466, n_0_465, n_0_464, n_0_463, n_0_462, n_0_461, 
      n_0_460, n_0_459}));
   datapath__0_45 i_0_38 (.p_0({uc_30, n_0_503, n_0_502, n_0_501, n_0_500, 
      n_0_499, n_0_498, n_0_497, n_0_496, n_0_495, n_0_494, n_0_493, n_0_492, 
      n_0_491, n_0_490, n_0_489, n_0_488, n_0_487, n_0_486, n_0_485, n_0_484, 
      n_0_483, n_0_482}), .p_1({uc_31, n_0_479, n_0_478, n_0_477, n_0_476, 
      n_0_475, n_0_474, n_0_473, n_0_472, n_0_471, n_0_470, n_0_469, n_0_468, 
      n_0_467, n_0_466, n_0_465, n_0_464, n_0_463, n_0_462, n_0_461, n_0_460, 
      n_0_459, n_0_74}), .divider({uc_32, n_0_525, n_0_524, n_0_523, n_0_522, 
      n_0_521, n_0_520, n_0_519, n_0_518, n_0_517, n_0_516, n_0_515, n_0_514, 
      n_0_513, n_0_512, n_0_511, n_0_510, n_0_509, n_0_508, n_0_507, n_0_506, 
      n_0_505, n_0_504}));
   datapath__0_49 i_0_41 (.p_0({uc_33, n_0_548, n_0_547, n_0_546, n_0_545, 
      n_0_544, n_0_543, n_0_542, n_0_541, n_0_540, n_0_539, n_0_538, n_0_537, 
      n_0_536, n_0_535, n_0_534, n_0_533, n_0_532, n_0_531, n_0_530, n_0_529, 
      n_0_528, n_0_527}), .p_1({uc_34, n_0_524, n_0_523, n_0_522, n_0_521, 
      n_0_520, n_0_519, n_0_518, n_0_517, n_0_516, n_0_515, n_0_514, n_0_513, 
      n_0_512, n_0_511, n_0_510, n_0_509, n_0_508, n_0_507, n_0_506, n_0_505, 
      n_0_504, n_0_73}), .divider({uc_35, n_0_570, n_0_569, n_0_568, n_0_567, 
      n_0_566, n_0_565, n_0_564, n_0_563, n_0_562, n_0_561, n_0_560, n_0_559, 
      n_0_558, n_0_557, n_0_556, n_0_555, n_0_554, n_0_553, n_0_552, n_0_551, 
      n_0_550, n_0_549}));
   datapath__0_53 i_0_44 (.p_0({uc_36, n_0_593, n_0_592, n_0_591, n_0_590, 
      n_0_589, n_0_588, n_0_587, n_0_586, n_0_585, n_0_584, n_0_583, n_0_582, 
      n_0_581, n_0_580, n_0_579, n_0_578, n_0_577, n_0_576, n_0_575, n_0_574, 
      n_0_573, n_0_572}), .p_1({uc_37, n_0_569, n_0_568, n_0_567, n_0_566, 
      n_0_565, n_0_564, n_0_563, n_0_562, n_0_561, n_0_560, n_0_559, n_0_558, 
      n_0_557, n_0_556, n_0_555, n_0_554, n_0_553, n_0_552, n_0_551, n_0_550, 
      n_0_549, n_0_72}), .divider({uc_38, n_0_615, n_0_614, n_0_613, n_0_612, 
      n_0_611, n_0_610, n_0_609, n_0_608, n_0_607, n_0_606, n_0_605, n_0_604, 
      n_0_603, n_0_602, n_0_601, n_0_600, n_0_599, n_0_598, n_0_597, n_0_596, 
      n_0_595, n_0_594}));
   datapath__0_57 i_0_47 (.p_0({uc_39, n_0_638, n_0_637, n_0_636, n_0_635, 
      n_0_634, n_0_633, n_0_632, n_0_631, n_0_630, n_0_629, n_0_628, n_0_627, 
      n_0_626, n_0_625, n_0_624, n_0_623, n_0_622, n_0_621, n_0_620, n_0_619, 
      n_0_618, n_0_617}), .p_1({uc_40, n_0_614, n_0_613, n_0_612, n_0_611, 
      n_0_610, n_0_609, n_0_608, n_0_607, n_0_606, n_0_605, n_0_604, n_0_603, 
      n_0_602, n_0_601, n_0_600, n_0_599, n_0_598, n_0_597, n_0_596, n_0_595, 
      n_0_594, n_0_71}), .divider({uc_41, n_0_660, n_0_659, n_0_658, n_0_657, 
      n_0_656, n_0_655, n_0_654, n_0_653, n_0_652, n_0_651, n_0_650, n_0_649, 
      n_0_648, n_0_647, n_0_646, n_0_645, n_0_644, n_0_643, n_0_642, n_0_641, 
      n_0_640, n_0_639}));
   datapath__0_61 i_0_50 (.p_0({uc_42, n_0_683, n_0_682, n_0_681, n_0_680, 
      n_0_679, n_0_678, n_0_677, n_0_676, n_0_675, n_0_674, n_0_673, n_0_672, 
      n_0_671, n_0_670, n_0_669, n_0_668, n_0_667, n_0_666, n_0_665, n_0_664, 
      n_0_663, n_0_662}), .p_1({uc_43, n_0_659, n_0_658, n_0_657, n_0_656, 
      n_0_655, n_0_654, n_0_653, n_0_652, n_0_651, n_0_650, n_0_649, n_0_648, 
      n_0_647, n_0_646, n_0_645, n_0_644, n_0_643, n_0_642, n_0_641, n_0_640, 
      n_0_639, n_0_70}), .divider({uc_44, n_0_705, n_0_704, n_0_703, n_0_702, 
      n_0_701, n_0_700, n_0_699, n_0_698, n_0_697, n_0_696, n_0_695, n_0_694, 
      n_0_693, n_0_692, n_0_691, n_0_690, n_0_689, n_0_688, n_0_687, n_0_686, 
      n_0_685, n_0_684}));
   datapath__0_65 i_0_53 (.p_0({uc_45, n_0_728, n_0_727, n_0_726, n_0_725, 
      n_0_724, n_0_723, n_0_722, n_0_721, n_0_720, n_0_719, n_0_718, n_0_717, 
      n_0_716, n_0_715, n_0_714, n_0_713, n_0_712, n_0_711, n_0_710, n_0_709, 
      n_0_708, n_0_707}), .p_1({uc_46, n_0_704, n_0_703, n_0_702, n_0_701, 
      n_0_700, n_0_699, n_0_698, n_0_697, n_0_696, n_0_695, n_0_694, n_0_693, 
      n_0_692, n_0_691, n_0_690, n_0_689, n_0_688, n_0_687, n_0_686, n_0_685, 
      n_0_684, n_0_69}), .divider({uc_47, n_0_750, n_0_749, n_0_748, n_0_747, 
      n_0_746, n_0_745, n_0_744, n_0_743, n_0_742, n_0_741, n_0_740, n_0_739, 
      n_0_738, n_0_737, n_0_736, n_0_735, n_0_734, n_0_733, n_0_732, n_0_731, 
      n_0_730, n_0_729}));
   datapath__0_69 i_0_56 (.p_0({uc_48, n_0_773, n_0_772, n_0_771, n_0_770, 
      n_0_769, n_0_768, n_0_767, n_0_766, n_0_765, n_0_764, n_0_763, n_0_762, 
      n_0_761, n_0_760, n_0_759, n_0_758, n_0_757, n_0_756, n_0_755, n_0_754, 
      n_0_753, n_0_752}), .p_1({uc_49, n_0_749, n_0_748, n_0_747, n_0_746, 
      n_0_745, n_0_744, n_0_743, n_0_742, n_0_741, n_0_740, n_0_739, n_0_738, 
      n_0_737, n_0_736, n_0_735, n_0_734, n_0_733, n_0_732, n_0_731, n_0_730, 
      n_0_729, in_a[0]}), .divider({uc_50, n_0_795, n_0_794, n_0_793, n_0_792, 
      n_0_791, n_0_790, n_0_789, n_0_788, n_0_787, n_0_786, n_0_785, n_0_784, 
      n_0_783, n_0_782, n_0_781, n_0_780, n_0_779, n_0_778, n_0_777, n_0_776, 
      n_0_775, n_0_774}));
   datapath__0_73 i_0_59 (.p_0({uc_51, n_0_818, n_0_817, n_0_816, n_0_815, 
      n_0_814, n_0_813, n_0_812, n_0_811, n_0_810, n_0_809, n_0_808, n_0_807, 
      n_0_806, n_0_805, n_0_804, n_0_803, n_0_802, n_0_801, n_0_800, n_0_799, 
      n_0_798, uc_52}), .p_1({uc_53, n_0_794, n_0_793, n_0_792, n_0_791, n_0_790, 
      n_0_789, n_0_788, n_0_787, n_0_786, n_0_785, n_0_784, n_0_783, n_0_782, 
      n_0_781, n_0_780, n_0_779, n_0_778, n_0_777, n_0_776, n_0_775, n_0_774, 
      1'b0}), .divider({uc_54, n_0_839, n_0_838, n_0_837, n_0_836, n_0_835, 
      n_0_834, n_0_833, n_0_832, n_0_831, n_0_830, n_0_829, n_0_828, n_0_827, 
      n_0_826, n_0_825, n_0_824, n_0_823, n_0_822, n_0_821, n_0_820, n_0_819, 
      uc_55}));
   datapath__0_77 i_0_62 (.p_0({uc_56, n_0_862, n_0_861, n_0_860, n_0_859, 
      n_0_858, n_0_857, n_0_856, n_0_855, n_0_854, n_0_853, n_0_852, n_0_851, 
      n_0_850, n_0_849, n_0_848, n_0_847, n_0_846, n_0_845, n_0_844, n_0_843, 
      n_0_842, uc_57}), .p_1({uc_58, n_0_838, n_0_837, n_0_836, n_0_835, n_0_834, 
      n_0_833, n_0_832, n_0_831, n_0_830, n_0_829, n_0_828, n_0_827, n_0_826, 
      n_0_825, n_0_824, n_0_823, n_0_822, n_0_821, n_0_820, n_0_819, n_0_797, 
      1'b0}), .divider({uc_59, n_0_883, n_0_882, n_0_881, n_0_880, n_0_879, 
      n_0_878, n_0_877, n_0_876, n_0_875, n_0_874, n_0_873, n_0_872, n_0_871, 
      n_0_870, n_0_869, n_0_868, n_0_867, n_0_866, n_0_865, n_0_864, n_0_863, 
      uc_60}));
   datapath__0_81 i_0_65 (.p_0({uc_61, n_0_906, n_0_905, n_0_904, n_0_903, 
      n_0_902, n_0_901, n_0_900, n_0_899, n_0_898, n_0_897, n_0_896, n_0_895, 
      n_0_894, n_0_893, n_0_892, n_0_891, n_0_890, n_0_889, n_0_888, n_0_887, 
      n_0_886, uc_62}), .p_1({uc_63, n_0_882, n_0_881, n_0_880, n_0_879, n_0_878, 
      n_0_877, n_0_876, n_0_875, n_0_874, n_0_873, n_0_872, n_0_871, n_0_870, 
      n_0_869, n_0_868, n_0_867, n_0_866, n_0_865, n_0_864, n_0_863, n_0_841, 
      1'b0}), .divider({uc_64, n_0_927, n_0_926, n_0_925, n_0_924, n_0_923, 
      n_0_922, n_0_921, n_0_920, n_0_919, n_0_918, n_0_917, n_0_916, n_0_915, 
      n_0_914, n_0_913, n_0_912, n_0_911, n_0_910, n_0_909, n_0_908, n_0_907, 
      uc_65}));
   datapath__0_85 i_0_68 (.p_0({uc_66, n_0_950, n_0_949, n_0_948, n_0_947, 
      n_0_946, n_0_945, n_0_944, n_0_943, n_0_942, n_0_941, n_0_940, n_0_939, 
      n_0_938, n_0_937, n_0_936, n_0_935, n_0_934, n_0_933, n_0_932, n_0_931, 
      n_0_930, uc_67}), .p_1({uc_68, n_0_926, n_0_925, n_0_924, n_0_923, n_0_922, 
      n_0_921, n_0_920, n_0_919, n_0_918, n_0_917, n_0_916, n_0_915, n_0_914, 
      n_0_913, n_0_912, n_0_911, n_0_910, n_0_909, n_0_908, n_0_907, n_0_885, 
      1'b0}), .divider({uc_69, n_0_971, n_0_970, n_0_969, n_0_968, n_0_967, 
      n_0_966, n_0_965, n_0_964, n_0_963, n_0_962, n_0_961, n_0_960, n_0_959, 
      n_0_958, n_0_957, n_0_956, n_0_955, n_0_954, n_0_953, n_0_952, n_0_951, 
      uc_70}));
   datapath__0_89 i_0_71 (.p_0({uc_71, n_0_994, n_0_993, n_0_992, n_0_991, 
      n_0_990, n_0_989, n_0_988, n_0_987, n_0_986, n_0_985, n_0_984, n_0_983, 
      n_0_982, n_0_981, n_0_980, n_0_979, n_0_978, n_0_977, n_0_976, n_0_975, 
      n_0_974, uc_72}), .p_1({uc_73, n_0_970, n_0_969, n_0_968, n_0_967, n_0_966, 
      n_0_965, n_0_964, n_0_963, n_0_962, n_0_961, n_0_960, n_0_959, n_0_958, 
      n_0_957, n_0_956, n_0_955, n_0_954, n_0_953, n_0_952, n_0_951, n_0_929, 
      1'b0}), .divider({uc_74, n_0_1015, n_0_1014, n_0_1013, n_0_1012, n_0_1011, 
      n_0_1010, n_0_1009, n_0_1008, n_0_1007, n_0_1006, n_0_1005, n_0_1004, 
      n_0_1003, n_0_1002, n_0_1001, n_0_1000, n_0_999, n_0_998, n_0_997, n_0_996, 
      n_0_995, uc_75}));
   datapath__0_93 i_0_74 (.p_0({uc_76, n_0_1038, n_0_1037, n_0_1036, n_0_1035, 
      n_0_1034, n_0_1033, n_0_1032, n_0_1031, n_0_1030, n_0_1029, n_0_1028, 
      n_0_1027, n_0_1026, n_0_1025, n_0_1024, n_0_1023, n_0_1022, n_0_1021, 
      n_0_1020, n_0_1019, n_0_1018, uc_77}), .p_1({uc_78, n_0_1014, n_0_1013, 
      n_0_1012, n_0_1011, n_0_1010, n_0_1009, n_0_1008, n_0_1007, n_0_1006, 
      n_0_1005, n_0_1004, n_0_1003, n_0_1002, n_0_1001, n_0_1000, n_0_999, 
      n_0_998, n_0_997, n_0_996, n_0_995, n_0_973, 1'b0}), .divider({uc_79, 
      n_0_1059, n_0_1058, n_0_1057, n_0_1056, n_0_1055, n_0_1054, n_0_1053, 
      n_0_1052, n_0_1051, n_0_1050, n_0_1049, n_0_1048, n_0_1047, n_0_1046, 
      n_0_1045, n_0_1044, n_0_1043, n_0_1042, n_0_1041, n_0_1040, n_0_1039, 
      uc_80}));
   datapath__0_103 i_0_83 (.plus({n_0_37, uc_81, uc_82, uc_83, uc_84, uc_85, 
      uc_86, uc_87, uc_88, uc_89, uc_90, uc_91, uc_92, uc_93, uc_94, uc_95, 
      uc_96, uc_97, uc_98, uc_99, uc_100, uc_101, uc_102, uc_103, uc_104, uc_105, 
      uc_106, uc_107, uc_108, uc_109, uc_110, uc_111, uc_112, uc_113, uc_114, 
      uc_115, uc_116, uc_117, uc_118, uc_119, uc_120, uc_121, uc_122, uc_123, 
      uc_124, uc_125, uc_126, uc_127, n_0_36, n_0_35, n_0_34, n_0_33, n_0_32, 
      n_0_31, n_0_30, n_0_29, n_0_28, n_0_27, n_0_26, n_0_25, n_0_24, n_0_23, 
      n_0_0, uc_128}), .p_0({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
      1'b0, 1'b0, 1'b0, 1'b0, n_0_68, n_0_67, n_0_66, n_0_65, n_0_64, n_0_63, 
      n_0_62, n_0_61, n_0_60, n_0_1072, n_0_1071, n_0_1070, n_0_1069, n_0_1068, 
      n_0_1067, n_0_1066}));
   DFFR_X1 zero_flag_reg (.D(n_0_43), .RN(n_0_39), .CK(n_0_38), .Q(zero), .QN());
   DFFR_X1 ovfl_flag_reg (.D(n_0_41), .RN(n_0_39), .CK(n_0_38), .Q(ovfl_flag), 
      .QN());
   DFFR_X1 divide_by_zero_error_reg (.D(n_0_1065), .RN(n_0_39), .CK(clk), 
      .Q(divide_by_zero_error), .QN());
   OR2_X1 divide_by_zero_error_reg_enable_mux_0 (.A1(n_0_40), .A2(
      divide_by_zero_error), .ZN(n_0_1065));
   DFFR_X1 ready_reg (.D(1'b1), .RN(n_0_39), .CK(n_0_38), .Q(done), .QN());
   DFFR_X1 \out64_reg[63]  (.D(n_0_59), .RN(n_0_39), .CK(n_0_38), .Q(out_c[16]), 
      .QN());
   DFFR_X1 \out64_reg[15]  (.D(n_0_58), .RN(n_0_39), .CK(n_0_38), .Q(out_c[15]), 
      .QN());
   DFFR_X1 \out64_reg[14]  (.D(n_0_57), .RN(n_0_39), .CK(n_0_38), .Q(out_c[14]), 
      .QN());
   DFFR_X1 \out64_reg[13]  (.D(n_0_56), .RN(n_0_39), .CK(n_0_38), .Q(out_c[13]), 
      .QN());
   DFFR_X1 \out64_reg[12]  (.D(n_0_55), .RN(n_0_39), .CK(n_0_38), .Q(out_c[12]), 
      .QN());
   DFFR_X1 \out64_reg[11]  (.D(n_0_54), .RN(n_0_39), .CK(n_0_38), .Q(out_c[11]), 
      .QN());
   DFFR_X1 \out64_reg[10]  (.D(n_0_53), .RN(n_0_39), .CK(n_0_38), .Q(out_c[10]), 
      .QN());
   DFFR_X1 \out64_reg[9]  (.D(n_0_52), .RN(n_0_39), .CK(n_0_38), .Q(out_c[9]), 
      .QN());
   DFFR_X1 \out64_reg[8]  (.D(n_0_51), .RN(n_0_39), .CK(n_0_38), .Q(out_c[8]), 
      .QN());
   DFFR_X1 \out64_reg[7]  (.D(n_0_50), .RN(n_0_39), .CK(n_0_38), .Q(out_c[7]), 
      .QN());
   DFFR_X1 \out64_reg[6]  (.D(n_0_49), .RN(n_0_39), .CK(n_0_38), .Q(out_c[6]), 
      .QN());
   DFFR_X1 \out64_reg[5]  (.D(n_0_48), .RN(n_0_39), .CK(n_0_38), .Q(out_c[5]), 
      .QN());
   DFFR_X1 \out64_reg[4]  (.D(n_0_47), .RN(n_0_39), .CK(n_0_38), .Q(out_c[4]), 
      .QN());
   DFFR_X1 \out64_reg[3]  (.D(n_0_46), .RN(n_0_39), .CK(n_0_38), .Q(out_c[3]), 
      .QN());
   DFFR_X1 \out64_reg[2]  (.D(n_0_45), .RN(n_0_39), .CK(n_0_38), .Q(out_c[2]), 
      .QN());
   DFFR_X1 \out64_reg[1]  (.D(n_0_44), .RN(n_0_39), .CK(n_0_38), .Q(out_c[1]), 
      .QN());
   DFFR_X1 \out64_reg[0]  (.D(n_0_1066), .RN(n_0_39), .CK(n_0_38), .Q(out_c[0]), 
      .QN());
   CLKGATETST_X1 clk_gate_ovfl_flag_reg (.CK(clk), .E(enbl), .SE(1'b0), .GCK(
      n_0_38));
   NOR4_X1 i_0_0_0 (.A1(n_0_0_14), .A2(n_0_0_10), .A3(n_0_0_5), .A4(n_0_0_0), 
      .ZN(n_0_40));
   NAND4_X1 i_0_0_1 (.A1(n_0_0_4), .A2(n_0_0_3), .A3(n_0_0_2), .A4(n_0_0_1), 
      .ZN(n_0_0_0));
   NOR4_X1 i_0_0_2 (.A1(in_b[34]), .A2(in_b[33]), .A3(in_b[32]), .A4(in_b[31]), 
      .ZN(n_0_0_1));
   NOR4_X1 i_0_0_3 (.A1(in_b[30]), .A2(in_b[29]), .A3(in_b[28]), .A4(in_b[27]), 
      .ZN(n_0_0_2));
   NOR4_X1 i_0_0_4 (.A1(in_b[42]), .A2(in_b[41]), .A3(in_b[40]), .A4(in_b[39]), 
      .ZN(n_0_0_3));
   NOR4_X1 i_0_0_5 (.A1(in_b[38]), .A2(in_b[37]), .A3(in_b[36]), .A4(in_b[35]), 
      .ZN(n_0_0_4));
   NAND4_X1 i_0_0_6 (.A1(n_0_0_9), .A2(n_0_0_8), .A3(n_0_0_7), .A4(n_0_0_6), 
      .ZN(n_0_0_5));
   NOR4_X1 i_0_0_7 (.A1(in_b[18]), .A2(in_b[17]), .A3(in_b[16]), .A4(in_b[15]), 
      .ZN(n_0_0_6));
   NOR4_X1 i_0_0_8 (.A1(in_b[14]), .A2(in_b[13]), .A3(in_b[12]), .A4(in_b[11]), 
      .ZN(n_0_0_7));
   NOR4_X1 i_0_0_9 (.A1(in_b[26]), .A2(in_b[23]), .A3(in_b[21]), .A4(in_b[20]), 
      .ZN(n_0_0_8));
   NOR4_X1 i_0_0_10 (.A1(in_b[25]), .A2(in_b[24]), .A3(in_b[22]), .A4(in_b[19]), 
      .ZN(n_0_0_9));
   NAND3_X1 i_0_0_11 (.A1(n_0_0_13), .A2(n_0_0_12), .A3(n_0_0_11), .ZN(n_0_0_10));
   NOR4_X1 i_0_0_12 (.A1(in_b[10]), .A2(in_b[9]), .A3(in_b[8]), .A4(in_b[7]), 
      .ZN(n_0_0_11));
   NOR4_X1 i_0_0_13 (.A1(in_b[6]), .A2(in_b[5]), .A3(in_b[4]), .A4(in_b[3]), 
      .ZN(n_0_0_12));
   NOR3_X1 i_0_0_14 (.A1(in_b[2]), .A2(in_b[1]), .A3(in_b[0]), .ZN(n_0_0_13));
   NAND4_X1 i_0_0_15 (.A1(enbl), .A2(n_0_0_15), .A3(n_0_0_862), .A4(n_0_0_20), 
      .ZN(n_0_0_14));
   AND4_X1 i_0_0_16 (.A1(n_0_0_19), .A2(n_0_0_18), .A3(n_0_0_17), .A4(n_0_0_16), 
      .ZN(n_0_0_15));
   NOR4_X1 i_0_0_17 (.A1(in_b[50]), .A2(in_b[49]), .A3(in_b[48]), .A4(in_b[47]), 
      .ZN(n_0_0_16));
   NOR4_X1 i_0_0_18 (.A1(in_b[46]), .A2(in_b[45]), .A3(in_b[44]), .A4(in_b[43]), 
      .ZN(n_0_0_17));
   NOR4_X1 i_0_0_19 (.A1(in_b[58]), .A2(in_b[57]), .A3(in_b[56]), .A4(in_b[55]), 
      .ZN(n_0_0_18));
   NOR4_X1 i_0_0_20 (.A1(in_b[54]), .A2(in_b[53]), .A3(in_b[52]), .A4(in_b[51]), 
      .ZN(n_0_0_19));
   NOR4_X1 i_0_0_21 (.A1(in_b[62]), .A2(in_b[61]), .A3(in_b[60]), .A4(in_b[59]), 
      .ZN(n_0_0_20));
   OR4_X1 i_0_0_22 (.A1(n_0_0_561), .A2(n_0_0_528), .A3(n_0_0_496), .A4(n_0_0_21), 
      .ZN(n_0_41));
   OR4_X1 i_0_0_23 (.A1(n_0_0_464), .A2(n_0_0_432), .A3(n_0_0_400), .A4(
      n_0_0_595), .ZN(n_0_0_21));
   OAI22_X1 i_0_0_24 (.A1(n_0_0_29), .A2(n_0_0_38), .B1(n_0_0_40), .B2(n_0_0_23), 
      .ZN(n_0_42));
   NAND2_X1 i_0_0_25 (.A1(n_0_0_28), .A2(n_0_0_22), .ZN(n_0_43));
   NAND3_X1 i_0_0_26 (.A1(n_0_0_23), .A2(n_0_0_41), .A3(n_0_0_833), .ZN(n_0_0_22));
   NOR3_X1 i_0_0_27 (.A1(n_0_0_24), .A2(n_0_32), .A3(n_0_33), .ZN(n_0_0_23));
   NAND3_X1 i_0_0_28 (.A1(n_0_0_27), .A2(n_0_0_26), .A3(n_0_0_25), .ZN(n_0_0_24));
   NOR2_X1 i_0_0_29 (.A1(n_0_34), .A2(n_0_31), .ZN(n_0_0_25));
   NOR3_X1 i_0_0_30 (.A1(n_0_30), .A2(n_0_29), .A3(n_0_28), .ZN(n_0_0_26));
   NOR2_X1 i_0_0_31 (.A1(n_0_37), .A2(n_0_35), .ZN(n_0_0_27));
   NAND2_X1 i_0_0_32 (.A1(n_0_0_39), .A2(n_0_0_29), .ZN(n_0_0_28));
   NOR3_X1 i_0_0_33 (.A1(n_0_67), .A2(n_0_66), .A3(n_0_0_30), .ZN(n_0_0_29));
   NAND4_X1 i_0_0_34 (.A1(n_0_0_270), .A2(n_0_0_238), .A3(n_0_0_206), .A4(
      n_0_0_31), .ZN(n_0_0_30));
   NOR3_X1 i_0_0_35 (.A1(n_0_62), .A2(n_0_61), .A3(n_0_60), .ZN(n_0_0_31));
   MUX2_X1 i_0_0_36 (.A(n_0_1067), .B(n_0_0), .S(n_0_0_41), .Z(n_0_44));
   MUX2_X1 i_0_0_37 (.A(n_0_1068), .B(n_0_23), .S(n_0_0_41), .Z(n_0_45));
   MUX2_X1 i_0_0_38 (.A(n_0_1069), .B(n_0_24), .S(n_0_0_41), .Z(n_0_46));
   OAI21_X1 i_0_0_39 (.A(n_0_0_32), .B1(n_0_0_666), .B2(n_0_0_41), .ZN(n_0_47));
   NAND2_X1 i_0_0_40 (.A1(n_0_0_41), .A2(n_0_25), .ZN(n_0_0_32));
   OAI21_X1 i_0_0_41 (.A(n_0_0_33), .B1(n_0_0_696), .B2(n_0_0_41), .ZN(n_0_48));
   NAND2_X1 i_0_0_42 (.A1(n_0_0_41), .A2(n_0_26), .ZN(n_0_0_33));
   MUX2_X1 i_0_0_43 (.A(n_0_1072), .B(n_0_27), .S(n_0_0_41), .Z(n_0_49));
   MUX2_X1 i_0_0_44 (.A(n_0_60), .B(n_0_28), .S(n_0_0_41), .Z(n_0_50));
   OAI21_X1 i_0_0_45 (.A(n_0_0_34), .B1(n_0_0_139), .B2(n_0_0_41), .ZN(n_0_51));
   NAND2_X1 i_0_0_46 (.A1(n_0_0_41), .A2(n_0_29), .ZN(n_0_0_34));
   MUX2_X1 i_0_0_47 (.A(n_0_62), .B(n_0_30), .S(n_0_0_41), .Z(n_0_52));
   OAI21_X1 i_0_0_48 (.A(n_0_0_35), .B1(n_0_0_206), .B2(n_0_0_41), .ZN(n_0_53));
   NAND2_X1 i_0_0_49 (.A1(n_0_0_41), .A2(n_0_31), .ZN(n_0_0_35));
   OAI21_X1 i_0_0_50 (.A(n_0_0_36), .B1(n_0_0_238), .B2(n_0_0_41), .ZN(n_0_54));
   NAND2_X1 i_0_0_51 (.A1(n_0_0_41), .A2(n_0_32), .ZN(n_0_0_36));
   OAI21_X1 i_0_0_52 (.A(n_0_0_37), .B1(n_0_0_270), .B2(n_0_0_41), .ZN(n_0_55));
   NAND2_X1 i_0_0_53 (.A1(n_0_0_41), .A2(n_0_33), .ZN(n_0_0_37));
   MUX2_X1 i_0_0_54 (.A(n_0_66), .B(n_0_34), .S(n_0_0_41), .Z(n_0_56));
   MUX2_X1 i_0_0_55 (.A(n_0_67), .B(n_0_35), .S(n_0_0_41), .Z(n_0_57));
   AOI21_X1 i_0_0_56 (.A(n_0_0_39), .B1(n_0_0_41), .B2(n_0_0_833), .ZN(n_0_58));
   INV_X1 i_0_0_57 (.A(n_0_0_39), .ZN(n_0_0_38));
   NOR2_X1 i_0_0_58 (.A1(n_0_68), .A2(n_0_0_41), .ZN(n_0_0_39));
   NAND2_X1 i_0_0_59 (.A1(n_0_0_833), .A2(n_0_0_41), .ZN(n_0_0_40));
   AND2_X1 i_0_0_60 (.A1(n_0_0_41), .A2(n_0_37), .ZN(n_0_59));
   XOR2_X1 i_0_0_61 (.A(in_b[15]), .B(in_a[15]), .Z(n_0_0_41));
   AOI21_X1 i_0_0_62 (.A(n_0_0_72), .B1(n_0_0_43), .B2(n_0_0_42), .ZN(n_0_1066));
   AOI22_X1 i_0_0_63 (.A1(n_0_1058), .A2(n_0_0_831), .B1(n_0_0_758), .B2(
      n_0_1059), .ZN(n_0_0_42));
   OAI221_X1 i_0_0_64 (.A(n_0_0_44), .B1(n_0_0_829), .B2(n_0_1057), .C1(n_0_1058), 
      .C2(n_0_0_831), .ZN(n_0_0_43));
   OAI21_X1 i_0_0_65 (.A(n_0_0_45), .B1(n_0_0_47), .B2(n_0_0_46), .ZN(n_0_0_44));
   AOI22_X1 i_0_0_66 (.A1(n_0_1057), .A2(n_0_0_829), .B1(n_0_0_827), .B2(
      n_0_1056), .ZN(n_0_0_45));
   OAI22_X1 i_0_0_67 (.A1(n_0_1056), .A2(n_0_0_827), .B1(n_0_0_825), .B2(
      n_0_1055), .ZN(n_0_0_46));
   AOI221_X1 i_0_0_68 (.A(n_0_0_48), .B1(n_0_0_823), .B2(n_0_1054), .C1(n_0_1055), 
      .C2(n_0_0_825), .ZN(n_0_0_47));
   INV_X1 i_0_0_69 (.A(n_0_0_49), .ZN(n_0_0_48));
   OAI221_X1 i_0_0_70 (.A(n_0_0_50), .B1(n_0_0_821), .B2(n_0_1053), .C1(n_0_1054), 
      .C2(n_0_0_823), .ZN(n_0_0_49));
   NAND3_X1 i_0_0_71 (.A1(n_0_0_71), .A2(n_0_0_52), .A3(n_0_0_51), .ZN(n_0_0_50));
   OAI221_X1 i_0_0_72 (.A(n_0_0_53), .B1(n_0_0_817), .B2(n_0_1051), .C1(n_0_1052), 
      .C2(n_0_0_819), .ZN(n_0_0_51));
   NAND2_X1 i_0_0_73 (.A1(n_0_0_819), .A2(n_0_1052), .ZN(n_0_0_52));
   OAI21_X1 i_0_0_74 (.A(n_0_0_54), .B1(n_0_0_56), .B2(n_0_0_55), .ZN(n_0_0_53));
   AOI22_X1 i_0_0_75 (.A1(n_0_1051), .A2(n_0_0_817), .B1(n_0_0_815), .B2(
      n_0_1050), .ZN(n_0_0_54));
   OAI22_X1 i_0_0_76 (.A1(n_0_1050), .A2(n_0_0_815), .B1(n_0_0_813), .B2(
      n_0_1049), .ZN(n_0_0_55));
   AOI221_X1 i_0_0_77 (.A(n_0_0_57), .B1(n_0_0_811), .B2(n_0_1048), .C1(n_0_1049), 
      .C2(n_0_0_813), .ZN(n_0_0_56));
   AOI21_X1 i_0_0_78 (.A(n_0_0_58), .B1(n_0_0_60), .B2(n_0_0_59), .ZN(n_0_0_57));
   OAI22_X1 i_0_0_79 (.A1(n_0_1048), .A2(n_0_0_811), .B1(n_0_0_809), .B2(
      n_0_1047), .ZN(n_0_0_58));
   AOI22_X1 i_0_0_80 (.A1(n_0_1047), .A2(n_0_0_809), .B1(n_0_0_807), .B2(
      n_0_1046), .ZN(n_0_0_59));
   OAI221_X1 i_0_0_81 (.A(n_0_0_61), .B1(n_0_0_805), .B2(n_0_1045), .C1(n_0_1046), 
      .C2(n_0_0_807), .ZN(n_0_0_60));
   OAI21_X1 i_0_0_82 (.A(n_0_0_62), .B1(n_0_0_64), .B2(n_0_0_63), .ZN(n_0_0_61));
   AOI22_X1 i_0_0_83 (.A1(n_0_1045), .A2(n_0_0_805), .B1(n_0_0_803), .B2(
      n_0_1044), .ZN(n_0_0_62));
   OAI22_X1 i_0_0_84 (.A1(n_0_1044), .A2(n_0_0_803), .B1(n_0_0_801), .B2(
      n_0_1043), .ZN(n_0_0_63));
   AOI21_X1 i_0_0_85 (.A(n_0_0_65), .B1(n_0_0_801), .B2(n_0_1043), .ZN(n_0_0_64));
   AOI21_X1 i_0_0_86 (.A(n_0_0_66), .B1(n_0_571), .B2(n_0_0_856), .ZN(n_0_0_65));
   AOI221_X1 i_0_0_87 (.A(n_0_0_67), .B1(n_0_0_797), .B2(n_0_1041), .C1(n_0_1042), 
      .C2(n_0_0_799), .ZN(n_0_0_66));
   AOI21_X1 i_0_0_88 (.A(n_0_0_68), .B1(n_0_0_70), .B2(n_0_0_69), .ZN(n_0_0_67));
   OAI22_X1 i_0_0_89 (.A1(n_0_1041), .A2(n_0_0_797), .B1(n_0_0_795), .B2(
      n_0_1040), .ZN(n_0_0_68));
   AOI22_X1 i_0_0_90 (.A1(n_0_1040), .A2(n_0_0_795), .B1(n_0_0_793), .B2(
      n_0_1039), .ZN(n_0_0_69));
   OAI221_X1 i_0_0_91 (.A(n_0_0_791), .B1(n_0_0_793), .B2(n_0_1039), .C1(
      n_0_1067), .C2(n_0_0_861), .ZN(n_0_0_70));
   NAND2_X1 i_0_0_92 (.A1(n_0_1053), .A2(n_0_0_821), .ZN(n_0_0_71));
   NOR2_X1 i_0_0_93 (.A1(n_0_1059), .A2(n_0_0_758), .ZN(n_0_0_72));
   NOR3_X1 i_0_0_94 (.A1(n_0_0_73), .A2(n_0_0_834), .A3(n_0_0_106), .ZN(n_0_1018));
   NOR3_X1 i_0_0_95 (.A1(n_0_0_73), .A2(n_0_0_835), .A3(n_0_0_106), .ZN(n_0_1019));
   NOR3_X1 i_0_0_96 (.A1(n_0_0_73), .A2(n_0_0_836), .A3(n_0_0_106), .ZN(n_0_1020));
   NOR3_X1 i_0_0_97 (.A1(n_0_0_73), .A2(n_0_0_837), .A3(n_0_0_106), .ZN(n_0_1021));
   NOR3_X1 i_0_0_98 (.A1(n_0_0_73), .A2(n_0_0_838), .A3(n_0_0_106), .ZN(n_0_1022));
   NOR3_X1 i_0_0_99 (.A1(n_0_0_73), .A2(n_0_0_839), .A3(n_0_0_106), .ZN(n_0_1023));
   NOR3_X1 i_0_0_100 (.A1(n_0_0_73), .A2(n_0_0_840), .A3(n_0_0_106), .ZN(
      n_0_1024));
   NOR3_X1 i_0_0_101 (.A1(n_0_0_73), .A2(n_0_0_841), .A3(n_0_0_106), .ZN(
      n_0_1025));
   NOR3_X1 i_0_0_102 (.A1(n_0_0_73), .A2(n_0_0_842), .A3(n_0_0_106), .ZN(
      n_0_1026));
   NOR3_X1 i_0_0_103 (.A1(n_0_0_73), .A2(n_0_0_843), .A3(n_0_0_106), .ZN(
      n_0_1027));
   NOR3_X1 i_0_0_104 (.A1(n_0_0_73), .A2(n_0_0_844), .A3(n_0_0_106), .ZN(
      n_0_1028));
   NOR3_X1 i_0_0_105 (.A1(n_0_0_73), .A2(n_0_0_845), .A3(n_0_0_106), .ZN(
      n_0_1029));
   NOR3_X1 i_0_0_106 (.A1(n_0_0_73), .A2(n_0_0_846), .A3(n_0_0_106), .ZN(
      n_0_1030));
   NOR3_X1 i_0_0_107 (.A1(n_0_0_73), .A2(n_0_0_847), .A3(n_0_0_106), .ZN(
      n_0_1031));
   NOR3_X1 i_0_0_108 (.A1(n_0_0_73), .A2(n_0_0_848), .A3(n_0_0_106), .ZN(
      n_0_1032));
   NOR3_X1 i_0_0_109 (.A1(n_0_0_73), .A2(n_0_0_849), .A3(n_0_0_106), .ZN(
      n_0_1033));
   NOR3_X1 i_0_0_110 (.A1(n_0_0_73), .A2(n_0_0_850), .A3(n_0_0_106), .ZN(
      n_0_1034));
   NOR3_X1 i_0_0_111 (.A1(n_0_0_73), .A2(n_0_0_851), .A3(n_0_0_106), .ZN(
      n_0_1035));
   NOR3_X1 i_0_0_112 (.A1(n_0_0_73), .A2(n_0_0_852), .A3(n_0_0_106), .ZN(
      n_0_1036));
   NOR3_X1 i_0_0_113 (.A1(n_0_0_73), .A2(n_0_0_853), .A3(n_0_0_106), .ZN(
      n_0_1037));
   NOR3_X1 i_0_0_114 (.A1(n_0_0_73), .A2(n_0_0_854), .A3(n_0_0_106), .ZN(
      n_0_1038));
   NOR2_X1 i_0_0_115 (.A1(n_0_0_106), .A2(n_0_0_73), .ZN(n_0_1067));
   AOI221_X1 i_0_0_116 (.A(n_0_0_74), .B1(n_0_0_831), .B2(n_0_1014), .C1(
      n_0_1015), .C2(n_0_0_758), .ZN(n_0_0_73));
   NOR2_X1 i_0_0_117 (.A1(n_0_0_76), .A2(n_0_0_75), .ZN(n_0_0_74));
   OAI22_X1 i_0_0_118 (.A1(n_0_1014), .A2(n_0_0_831), .B1(n_0_0_829), .B2(
      n_0_1013), .ZN(n_0_0_75));
   AOI221_X1 i_0_0_119 (.A(n_0_0_77), .B1(n_0_0_827), .B2(n_0_1012), .C1(
      n_0_1013), .C2(n_0_0_829), .ZN(n_0_0_76));
   NOR3_X1 i_0_0_120 (.A1(n_0_0_105), .A2(n_0_0_104), .A3(n_0_0_78), .ZN(
      n_0_0_77));
   AOI221_X1 i_0_0_121 (.A(n_0_0_79), .B1(n_0_0_823), .B2(n_0_1010), .C1(
      n_0_1011), .C2(n_0_0_825), .ZN(n_0_0_78));
   AOI21_X1 i_0_0_122 (.A(n_0_0_103), .B1(n_0_0_102), .B2(n_0_0_80), .ZN(
      n_0_0_79));
   OAI221_X1 i_0_0_123 (.A(n_0_0_81), .B1(n_0_0_819), .B2(n_0_1008), .C1(
      n_0_1009), .C2(n_0_0_821), .ZN(n_0_0_80));
   NAND2_X1 i_0_0_124 (.A1(n_0_0_83), .A2(n_0_0_82), .ZN(n_0_0_81));
   AOI22_X1 i_0_0_125 (.A1(n_0_1007), .A2(n_0_0_817), .B1(n_0_0_819), .B2(
      n_0_1008), .ZN(n_0_0_82));
   OAI221_X1 i_0_0_126 (.A(n_0_0_84), .B1(n_0_0_815), .B2(n_0_1006), .C1(
      n_0_1007), .C2(n_0_0_817), .ZN(n_0_0_83));
   OAI21_X1 i_0_0_127 (.A(n_0_0_85), .B1(n_0_0_87), .B2(n_0_0_86), .ZN(n_0_0_84));
   AOI22_X1 i_0_0_128 (.A1(n_0_1006), .A2(n_0_0_815), .B1(n_0_0_813), .B2(
      n_0_1005), .ZN(n_0_0_85));
   OAI22_X1 i_0_0_129 (.A1(n_0_1005), .A2(n_0_0_813), .B1(n_0_0_811), .B2(
      n_0_1004), .ZN(n_0_0_86));
   AOI21_X1 i_0_0_130 (.A(n_0_0_88), .B1(n_0_0_811), .B2(n_0_1004), .ZN(n_0_0_87));
   AOI21_X1 i_0_0_131 (.A(n_0_0_101), .B1(n_0_0_90), .B2(n_0_0_89), .ZN(n_0_0_88));
   AOI22_X1 i_0_0_132 (.A1(n_0_1003), .A2(n_0_0_809), .B1(n_0_0_807), .B2(
      n_0_1002), .ZN(n_0_0_89));
   OAI221_X1 i_0_0_133 (.A(n_0_0_91), .B1(n_0_0_805), .B2(n_0_1001), .C1(
      n_0_1002), .C2(n_0_0_807), .ZN(n_0_0_90));
   OAI21_X1 i_0_0_134 (.A(n_0_0_92), .B1(n_0_0_94), .B2(n_0_0_93), .ZN(n_0_0_91));
   AOI22_X1 i_0_0_135 (.A1(n_0_1001), .A2(n_0_0_805), .B1(n_0_0_803), .B2(
      n_0_1000), .ZN(n_0_0_92));
   OAI22_X1 i_0_0_136 (.A1(n_0_1000), .A2(n_0_0_803), .B1(n_0_0_801), .B2(
      n_0_999), .ZN(n_0_0_93));
   AOI21_X1 i_0_0_137 (.A(n_0_0_95), .B1(n_0_0_801), .B2(n_0_999), .ZN(n_0_0_94));
   AOI21_X1 i_0_0_138 (.A(n_0_0_96), .B1(n_0_571), .B2(n_0_0_857), .ZN(n_0_0_95));
   AOI221_X1 i_0_0_139 (.A(n_0_0_97), .B1(n_0_0_797), .B2(n_0_997), .C1(n_0_998), 
      .C2(n_0_0_799), .ZN(n_0_0_96));
   AOI21_X1 i_0_0_140 (.A(n_0_0_98), .B1(n_0_0_100), .B2(n_0_0_99), .ZN(n_0_0_97));
   OAI22_X1 i_0_0_141 (.A1(n_0_997), .A2(n_0_0_797), .B1(n_0_0_795), .B2(n_0_996), 
      .ZN(n_0_0_98));
   AOI22_X1 i_0_0_142 (.A1(n_0_996), .A2(n_0_0_795), .B1(n_0_0_793), .B2(n_0_995), 
      .ZN(n_0_0_99));
   OAI221_X1 i_0_0_143 (.A(n_0_0_791), .B1(n_0_0_793), .B2(n_0_995), .C1(
      n_0_1068), .C2(n_0_0_861), .ZN(n_0_0_100));
   NOR2_X1 i_0_0_144 (.A1(n_0_1003), .A2(n_0_0_809), .ZN(n_0_0_101));
   NAND2_X1 i_0_0_145 (.A1(n_0_1009), .A2(n_0_0_821), .ZN(n_0_0_102));
   NOR2_X1 i_0_0_146 (.A1(n_0_1010), .A2(n_0_0_823), .ZN(n_0_0_103));
   NOR2_X1 i_0_0_147 (.A1(n_0_1011), .A2(n_0_0_825), .ZN(n_0_0_104));
   NOR2_X1 i_0_0_148 (.A1(n_0_1012), .A2(n_0_0_827), .ZN(n_0_0_105));
   NOR2_X1 i_0_0_149 (.A1(n_0_1015), .A2(n_0_0_758), .ZN(n_0_0_106));
   AND2_X1 i_0_0_150 (.A1(n_0_60), .A2(in_b[0]), .ZN(n_0_752));
   AND2_X1 i_0_0_151 (.A1(n_0_60), .A2(n_0_78), .ZN(n_0_753));
   AND2_X1 i_0_0_152 (.A1(n_0_60), .A2(n_0_79), .ZN(n_0_754));
   AND2_X1 i_0_0_153 (.A1(n_0_60), .A2(n_0_80), .ZN(n_0_755));
   AND2_X1 i_0_0_154 (.A1(n_0_60), .A2(n_0_81), .ZN(n_0_756));
   AND2_X1 i_0_0_155 (.A1(n_0_60), .A2(n_0_82), .ZN(n_0_757));
   AND2_X1 i_0_0_156 (.A1(n_0_60), .A2(n_0_83), .ZN(n_0_758));
   AND2_X1 i_0_0_157 (.A1(n_0_60), .A2(n_0_84), .ZN(n_0_759));
   AND2_X1 i_0_0_158 (.A1(n_0_60), .A2(n_0_85), .ZN(n_0_760));
   AND2_X1 i_0_0_159 (.A1(n_0_60), .A2(n_0_86), .ZN(n_0_761));
   AND2_X1 i_0_0_160 (.A1(n_0_60), .A2(n_0_87), .ZN(n_0_762));
   AND2_X1 i_0_0_161 (.A1(n_0_60), .A2(n_0_88), .ZN(n_0_763));
   AND2_X1 i_0_0_162 (.A1(n_0_60), .A2(n_0_89), .ZN(n_0_764));
   AND2_X1 i_0_0_163 (.A1(n_0_60), .A2(n_0_90), .ZN(n_0_765));
   AND2_X1 i_0_0_164 (.A1(n_0_60), .A2(n_0_91), .ZN(n_0_766));
   AND2_X1 i_0_0_165 (.A1(n_0_60), .A2(n_0_92), .ZN(n_0_767));
   AND2_X1 i_0_0_166 (.A1(n_0_60), .A2(n_0_93), .ZN(n_0_768));
   AND2_X1 i_0_0_167 (.A1(n_0_60), .A2(n_0_94), .ZN(n_0_769));
   AND2_X1 i_0_0_168 (.A1(n_0_60), .A2(n_0_95), .ZN(n_0_770));
   AND2_X1 i_0_0_169 (.A1(n_0_60), .A2(n_0_96), .ZN(n_0_771));
   AND2_X1 i_0_0_170 (.A1(n_0_60), .A2(n_0_97), .ZN(n_0_772));
   AND2_X1 i_0_0_171 (.A1(n_0_60), .A2(n_0_98), .ZN(n_0_773));
   NAND2_X1 i_0_0_172 (.A1(n_0_0_138), .A2(n_0_0_107), .ZN(n_0_60));
   OAI221_X1 i_0_0_173 (.A(n_0_0_108), .B1(n_0_0_831), .B2(n_0_749), .C1(n_0_750), 
      .C2(n_0_0_758), .ZN(n_0_0_107));
   NAND2_X1 i_0_0_174 (.A1(n_0_0_110), .A2(n_0_0_109), .ZN(n_0_0_108));
   AOI22_X1 i_0_0_175 (.A1(n_0_749), .A2(n_0_0_831), .B1(n_0_0_829), .B2(n_0_748), 
      .ZN(n_0_0_109));
   OAI221_X1 i_0_0_176 (.A(n_0_0_111), .B1(n_0_0_827), .B2(n_0_747), .C1(n_0_748), 
      .C2(n_0_0_829), .ZN(n_0_0_110));
   NAND2_X1 i_0_0_177 (.A1(n_0_0_113), .A2(n_0_0_112), .ZN(n_0_0_111));
   AOI22_X1 i_0_0_178 (.A1(n_0_747), .A2(n_0_0_827), .B1(n_0_0_825), .B2(n_0_746), 
      .ZN(n_0_0_112));
   OAI221_X1 i_0_0_179 (.A(n_0_0_114), .B1(n_0_0_823), .B2(n_0_745), .C1(n_0_746), 
      .C2(n_0_0_825), .ZN(n_0_0_113));
   NAND2_X1 i_0_0_180 (.A1(n_0_0_116), .A2(n_0_0_115), .ZN(n_0_0_114));
   AOI22_X1 i_0_0_181 (.A1(n_0_745), .A2(n_0_0_823), .B1(n_0_0_821), .B2(n_0_744), 
      .ZN(n_0_0_115));
   OAI221_X1 i_0_0_182 (.A(n_0_0_117), .B1(n_0_0_819), .B2(n_0_743), .C1(n_0_744), 
      .C2(n_0_0_821), .ZN(n_0_0_116));
   OAI21_X1 i_0_0_183 (.A(n_0_0_118), .B1(n_0_0_120), .B2(n_0_0_119), .ZN(
      n_0_0_117));
   AOI22_X1 i_0_0_184 (.A1(n_0_742), .A2(n_0_0_817), .B1(n_0_0_819), .B2(n_0_743), 
      .ZN(n_0_0_118));
   OAI22_X1 i_0_0_185 (.A1(n_0_742), .A2(n_0_0_817), .B1(n_0_0_815), .B2(n_0_741), 
      .ZN(n_0_0_119));
   AOI221_X1 i_0_0_186 (.A(n_0_0_121), .B1(n_0_0_813), .B2(n_0_740), .C1(n_0_741), 
      .C2(n_0_0_815), .ZN(n_0_0_120));
   AOI21_X1 i_0_0_187 (.A(n_0_0_122), .B1(n_0_0_124), .B2(n_0_0_123), .ZN(
      n_0_0_121));
   OAI22_X1 i_0_0_188 (.A1(n_0_740), .A2(n_0_0_813), .B1(n_0_0_811), .B2(n_0_739), 
      .ZN(n_0_0_122));
   AOI22_X1 i_0_0_189 (.A1(n_0_739), .A2(n_0_0_811), .B1(n_0_0_809), .B2(n_0_738), 
      .ZN(n_0_0_123));
   OAI221_X1 i_0_0_190 (.A(n_0_0_125), .B1(n_0_0_807), .B2(n_0_737), .C1(n_0_738), 
      .C2(n_0_0_809), .ZN(n_0_0_124));
   OAI21_X1 i_0_0_191 (.A(n_0_0_126), .B1(n_0_0_128), .B2(n_0_0_127), .ZN(
      n_0_0_125));
   AOI22_X1 i_0_0_192 (.A1(n_0_737), .A2(n_0_0_807), .B1(n_0_0_805), .B2(n_0_736), 
      .ZN(n_0_0_126));
   OAI22_X1 i_0_0_193 (.A1(n_0_736), .A2(n_0_0_805), .B1(n_0_0_803), .B2(n_0_735), 
      .ZN(n_0_0_127));
   AOI221_X1 i_0_0_194 (.A(n_0_0_129), .B1(n_0_0_801), .B2(n_0_734), .C1(n_0_735), 
      .C2(n_0_0_803), .ZN(n_0_0_128));
   AOI21_X1 i_0_0_195 (.A(n_0_0_130), .B1(n_0_0_132), .B2(n_0_0_131), .ZN(
      n_0_0_129));
   OAI22_X1 i_0_0_196 (.A1(n_0_734), .A2(n_0_0_801), .B1(n_0_0_799), .B2(n_0_733), 
      .ZN(n_0_0_130));
   AOI22_X1 i_0_0_197 (.A1(n_0_733), .A2(n_0_0_799), .B1(n_0_0_797), .B2(n_0_732), 
      .ZN(n_0_0_131));
   OAI22_X1 i_0_0_198 (.A1(n_0_732), .A2(n_0_0_797), .B1(n_0_0_137), .B2(
      n_0_0_133), .ZN(n_0_0_132));
   AOI21_X1 i_0_0_199 (.A(n_0_0_134), .B1(n_0_0_135), .B2(n_0_0_136), .ZN(
      n_0_0_133));
   OAI22_X1 i_0_0_200 (.A1(n_0_731), .A2(n_0_0_795), .B1(n_0_0_793), .B2(n_0_730), 
      .ZN(n_0_0_134));
   AOI22_X1 i_0_0_201 (.A1(n_0_730), .A2(n_0_0_793), .B1(n_0_0_791), .B2(n_0_729), 
      .ZN(n_0_0_135));
   OAI22_X1 i_0_0_202 (.A1(n_0_729), .A2(n_0_0_791), .B1(n_0_0_861), .B2(in_a[0]), 
      .ZN(n_0_0_136));
   AND2_X1 i_0_0_203 (.A1(n_0_731), .A2(n_0_0_795), .ZN(n_0_0_137));
   NAND2_X1 i_0_0_204 (.A1(n_0_750), .A2(n_0_0_758), .ZN(n_0_0_138));
   NOR2_X1 i_0_0_205 (.A1(n_0_0_139), .A2(n_0_0_861), .ZN(n_0_707));
   NOR2_X1 i_0_0_206 (.A1(n_0_0_139), .A2(n_0_0_834), .ZN(n_0_708));
   NOR2_X1 i_0_0_207 (.A1(n_0_0_139), .A2(n_0_0_835), .ZN(n_0_709));
   NOR2_X1 i_0_0_208 (.A1(n_0_0_139), .A2(n_0_0_836), .ZN(n_0_710));
   NOR2_X1 i_0_0_209 (.A1(n_0_0_139), .A2(n_0_0_837), .ZN(n_0_711));
   NOR2_X1 i_0_0_210 (.A1(n_0_0_139), .A2(n_0_0_838), .ZN(n_0_712));
   NOR2_X1 i_0_0_211 (.A1(n_0_0_139), .A2(n_0_0_839), .ZN(n_0_713));
   NOR2_X1 i_0_0_212 (.A1(n_0_0_139), .A2(n_0_0_840), .ZN(n_0_714));
   NOR2_X1 i_0_0_213 (.A1(n_0_0_139), .A2(n_0_0_841), .ZN(n_0_715));
   NOR2_X1 i_0_0_214 (.A1(n_0_0_139), .A2(n_0_0_842), .ZN(n_0_716));
   NOR2_X1 i_0_0_215 (.A1(n_0_0_139), .A2(n_0_0_843), .ZN(n_0_717));
   NOR2_X1 i_0_0_216 (.A1(n_0_0_139), .A2(n_0_0_844), .ZN(n_0_718));
   NOR2_X1 i_0_0_217 (.A1(n_0_0_139), .A2(n_0_0_845), .ZN(n_0_719));
   NOR2_X1 i_0_0_218 (.A1(n_0_0_139), .A2(n_0_0_846), .ZN(n_0_720));
   NOR2_X1 i_0_0_219 (.A1(n_0_0_139), .A2(n_0_0_847), .ZN(n_0_721));
   NOR2_X1 i_0_0_220 (.A1(n_0_0_139), .A2(n_0_0_848), .ZN(n_0_722));
   NOR2_X1 i_0_0_221 (.A1(n_0_0_139), .A2(n_0_0_849), .ZN(n_0_723));
   NOR2_X1 i_0_0_222 (.A1(n_0_0_139), .A2(n_0_0_850), .ZN(n_0_724));
   NOR2_X1 i_0_0_223 (.A1(n_0_0_139), .A2(n_0_0_851), .ZN(n_0_725));
   NOR2_X1 i_0_0_224 (.A1(n_0_0_139), .A2(n_0_0_852), .ZN(n_0_726));
   NOR2_X1 i_0_0_225 (.A1(n_0_0_139), .A2(n_0_0_853), .ZN(n_0_727));
   NOR2_X1 i_0_0_226 (.A1(n_0_0_139), .A2(n_0_0_854), .ZN(n_0_728));
   INV_X1 i_0_0_227 (.A(n_0_0_139), .ZN(n_0_61));
   AOI21_X1 i_0_0_228 (.A(n_0_0_140), .B1(n_0_0_758), .B2(n_0_705), .ZN(
      n_0_0_139));
   AOI21_X1 i_0_0_229 (.A(n_0_0_141), .B1(n_0_0_143), .B2(n_0_0_142), .ZN(
      n_0_0_140));
   OAI22_X1 i_0_0_230 (.A1(n_0_704), .A2(n_0_0_831), .B1(n_0_0_758), .B2(n_0_705), 
      .ZN(n_0_0_141));
   AOI22_X1 i_0_0_231 (.A1(n_0_704), .A2(n_0_0_831), .B1(n_0_0_829), .B2(n_0_703), 
      .ZN(n_0_0_142));
   OAI21_X1 i_0_0_232 (.A(n_0_0_144), .B1(n_0_0_829), .B2(n_0_703), .ZN(
      n_0_0_143));
   OAI21_X1 i_0_0_233 (.A(n_0_0_172), .B1(n_0_0_146), .B2(n_0_0_145), .ZN(
      n_0_0_144));
   OAI22_X1 i_0_0_234 (.A1(n_0_702), .A2(n_0_0_827), .B1(n_0_0_825), .B2(n_0_701), 
      .ZN(n_0_0_145));
   AOI221_X1 i_0_0_235 (.A(n_0_0_147), .B1(n_0_0_823), .B2(n_0_700), .C1(n_0_701), 
      .C2(n_0_0_825), .ZN(n_0_0_146));
   AOI21_X1 i_0_0_236 (.A(n_0_0_148), .B1(n_0_0_150), .B2(n_0_0_149), .ZN(
      n_0_0_147));
   OAI22_X1 i_0_0_237 (.A1(n_0_700), .A2(n_0_0_823), .B1(n_0_0_821), .B2(n_0_699), 
      .ZN(n_0_0_148));
   AOI22_X1 i_0_0_238 (.A1(n_0_699), .A2(n_0_0_821), .B1(n_0_0_819), .B2(n_0_698), 
      .ZN(n_0_0_149));
   OAI221_X1 i_0_0_239 (.A(n_0_0_151), .B1(n_0_0_817), .B2(n_0_697), .C1(n_0_698), 
      .C2(n_0_0_819), .ZN(n_0_0_150));
   OAI21_X1 i_0_0_240 (.A(n_0_0_152), .B1(n_0_0_154), .B2(n_0_0_153), .ZN(
      n_0_0_151));
   AOI22_X1 i_0_0_241 (.A1(n_0_697), .A2(n_0_0_817), .B1(n_0_0_815), .B2(n_0_696), 
      .ZN(n_0_0_152));
   OAI22_X1 i_0_0_242 (.A1(n_0_696), .A2(n_0_0_815), .B1(n_0_0_813), .B2(n_0_695), 
      .ZN(n_0_0_153));
   AOI221_X1 i_0_0_243 (.A(n_0_0_155), .B1(n_0_0_811), .B2(n_0_694), .C1(n_0_695), 
      .C2(n_0_0_813), .ZN(n_0_0_154));
   AOI21_X1 i_0_0_244 (.A(n_0_0_156), .B1(n_0_0_158), .B2(n_0_0_157), .ZN(
      n_0_0_155));
   OAI22_X1 i_0_0_245 (.A1(n_0_694), .A2(n_0_0_811), .B1(n_0_0_809), .B2(n_0_693), 
      .ZN(n_0_0_156));
   AOI22_X1 i_0_0_246 (.A1(n_0_693), .A2(n_0_0_809), .B1(n_0_0_807), .B2(n_0_692), 
      .ZN(n_0_0_157));
   OAI221_X1 i_0_0_247 (.A(n_0_0_159), .B1(n_0_0_805), .B2(n_0_691), .C1(n_0_692), 
      .C2(n_0_0_807), .ZN(n_0_0_158));
   OAI21_X1 i_0_0_248 (.A(n_0_0_160), .B1(n_0_0_162), .B2(n_0_0_161), .ZN(
      n_0_0_159));
   AOI22_X1 i_0_0_249 (.A1(n_0_691), .A2(n_0_0_805), .B1(n_0_0_803), .B2(n_0_690), 
      .ZN(n_0_0_160));
   OAI22_X1 i_0_0_250 (.A1(n_0_690), .A2(n_0_0_803), .B1(n_0_0_801), .B2(n_0_689), 
      .ZN(n_0_0_161));
   AOI221_X1 i_0_0_251 (.A(n_0_0_163), .B1(n_0_0_799), .B2(n_0_688), .C1(n_0_689), 
      .C2(n_0_0_801), .ZN(n_0_0_162));
   AOI21_X1 i_0_0_252 (.A(n_0_0_164), .B1(n_0_0_165), .B2(n_0_0_171), .ZN(
      n_0_0_163));
   OAI22_X1 i_0_0_253 (.A1(n_0_688), .A2(n_0_0_799), .B1(n_0_0_797), .B2(n_0_687), 
      .ZN(n_0_0_164));
   OAI21_X1 i_0_0_254 (.A(n_0_0_166), .B1(n_0_0_795), .B2(n_0_686), .ZN(
      n_0_0_165));
   INV_X1 i_0_0_255 (.A(n_0_0_167), .ZN(n_0_0_166));
   AOI221_X1 i_0_0_256 (.A(n_0_0_168), .B1(n_0_0_793), .B2(n_0_685), .C1(n_0_686), 
      .C2(n_0_0_795), .ZN(n_0_0_167));
   AOI21_X1 i_0_0_257 (.A(n_0_0_169), .B1(n_0_0_170), .B2(in_b[0]), .ZN(
      n_0_0_168));
   OAI22_X1 i_0_0_258 (.A1(n_0_685), .A2(n_0_0_793), .B1(n_0_0_791), .B2(n_0_684), 
      .ZN(n_0_0_169));
   AOI21_X1 i_0_0_259 (.A(n_0_69), .B1(n_0_0_791), .B2(n_0_684), .ZN(n_0_0_170));
   NAND2_X1 i_0_0_260 (.A1(n_0_687), .A2(n_0_0_797), .ZN(n_0_0_171));
   NAND2_X1 i_0_0_261 (.A1(n_0_702), .A2(n_0_0_827), .ZN(n_0_0_172));
   AND2_X1 i_0_0_262 (.A1(n_0_62), .A2(in_b[0]), .ZN(n_0_662));
   AND2_X1 i_0_0_263 (.A1(n_0_62), .A2(n_0_78), .ZN(n_0_663));
   AND2_X1 i_0_0_264 (.A1(n_0_62), .A2(n_0_79), .ZN(n_0_664));
   AND2_X1 i_0_0_265 (.A1(n_0_62), .A2(n_0_80), .ZN(n_0_665));
   AND2_X1 i_0_0_266 (.A1(n_0_62), .A2(n_0_81), .ZN(n_0_666));
   AND2_X1 i_0_0_267 (.A1(n_0_62), .A2(n_0_82), .ZN(n_0_667));
   AND2_X1 i_0_0_268 (.A1(n_0_62), .A2(n_0_83), .ZN(n_0_668));
   AND2_X1 i_0_0_269 (.A1(n_0_62), .A2(n_0_84), .ZN(n_0_669));
   AND2_X1 i_0_0_270 (.A1(n_0_62), .A2(n_0_85), .ZN(n_0_670));
   AND2_X1 i_0_0_271 (.A1(n_0_62), .A2(n_0_86), .ZN(n_0_671));
   AND2_X1 i_0_0_272 (.A1(n_0_62), .A2(n_0_87), .ZN(n_0_672));
   AND2_X1 i_0_0_273 (.A1(n_0_62), .A2(n_0_88), .ZN(n_0_673));
   AND2_X1 i_0_0_274 (.A1(n_0_62), .A2(n_0_89), .ZN(n_0_674));
   AND2_X1 i_0_0_275 (.A1(n_0_62), .A2(n_0_90), .ZN(n_0_675));
   AND2_X1 i_0_0_276 (.A1(n_0_62), .A2(n_0_91), .ZN(n_0_676));
   AND2_X1 i_0_0_277 (.A1(n_0_62), .A2(n_0_92), .ZN(n_0_677));
   AND2_X1 i_0_0_278 (.A1(n_0_62), .A2(n_0_93), .ZN(n_0_678));
   AND2_X1 i_0_0_279 (.A1(n_0_62), .A2(n_0_94), .ZN(n_0_679));
   AND2_X1 i_0_0_280 (.A1(n_0_62), .A2(n_0_95), .ZN(n_0_680));
   AND2_X1 i_0_0_281 (.A1(n_0_62), .A2(n_0_96), .ZN(n_0_681));
   AND2_X1 i_0_0_282 (.A1(n_0_62), .A2(n_0_97), .ZN(n_0_682));
   AND2_X1 i_0_0_283 (.A1(n_0_62), .A2(n_0_98), .ZN(n_0_683));
   NAND2_X1 i_0_0_284 (.A1(n_0_0_205), .A2(n_0_0_173), .ZN(n_0_62));
   OAI221_X1 i_0_0_285 (.A(n_0_0_174), .B1(n_0_0_831), .B2(n_0_659), .C1(n_0_660), 
      .C2(n_0_0_758), .ZN(n_0_0_173));
   NAND2_X1 i_0_0_286 (.A1(n_0_0_176), .A2(n_0_0_175), .ZN(n_0_0_174));
   AOI22_X1 i_0_0_287 (.A1(n_0_659), .A2(n_0_0_831), .B1(n_0_0_829), .B2(n_0_658), 
      .ZN(n_0_0_175));
   OAI221_X1 i_0_0_288 (.A(n_0_0_177), .B1(n_0_0_827), .B2(n_0_657), .C1(n_0_658), 
      .C2(n_0_0_829), .ZN(n_0_0_176));
   NAND2_X1 i_0_0_289 (.A1(n_0_0_179), .A2(n_0_0_178), .ZN(n_0_0_177));
   AOI22_X1 i_0_0_290 (.A1(n_0_657), .A2(n_0_0_827), .B1(n_0_0_825), .B2(n_0_656), 
      .ZN(n_0_0_178));
   OAI221_X1 i_0_0_291 (.A(n_0_0_180), .B1(n_0_0_823), .B2(n_0_655), .C1(n_0_656), 
      .C2(n_0_0_825), .ZN(n_0_0_179));
   NAND2_X1 i_0_0_292 (.A1(n_0_0_182), .A2(n_0_0_181), .ZN(n_0_0_180));
   AOI22_X1 i_0_0_293 (.A1(n_0_655), .A2(n_0_0_823), .B1(n_0_0_821), .B2(n_0_654), 
      .ZN(n_0_0_181));
   OAI221_X1 i_0_0_294 (.A(n_0_0_183), .B1(n_0_0_819), .B2(n_0_653), .C1(n_0_654), 
      .C2(n_0_0_821), .ZN(n_0_0_182));
   OAI21_X1 i_0_0_295 (.A(n_0_0_184), .B1(n_0_0_186), .B2(n_0_0_185), .ZN(
      n_0_0_183));
   AOI22_X1 i_0_0_296 (.A1(n_0_652), .A2(n_0_0_817), .B1(n_0_0_819), .B2(n_0_653), 
      .ZN(n_0_0_184));
   OAI22_X1 i_0_0_297 (.A1(n_0_652), .A2(n_0_0_817), .B1(n_0_0_815), .B2(n_0_651), 
      .ZN(n_0_0_185));
   AOI221_X1 i_0_0_298 (.A(n_0_0_187), .B1(n_0_0_813), .B2(n_0_650), .C1(n_0_651), 
      .C2(n_0_0_815), .ZN(n_0_0_186));
   AOI21_X1 i_0_0_299 (.A(n_0_0_188), .B1(n_0_0_190), .B2(n_0_0_189), .ZN(
      n_0_0_187));
   OAI22_X1 i_0_0_300 (.A1(n_0_650), .A2(n_0_0_813), .B1(n_0_0_811), .B2(n_0_649), 
      .ZN(n_0_0_188));
   AOI22_X1 i_0_0_301 (.A1(n_0_649), .A2(n_0_0_811), .B1(n_0_0_809), .B2(n_0_648), 
      .ZN(n_0_0_189));
   OAI221_X1 i_0_0_302 (.A(n_0_0_191), .B1(n_0_0_807), .B2(n_0_647), .C1(n_0_648), 
      .C2(n_0_0_809), .ZN(n_0_0_190));
   OAI21_X1 i_0_0_303 (.A(n_0_0_192), .B1(n_0_0_194), .B2(n_0_0_193), .ZN(
      n_0_0_191));
   AOI22_X1 i_0_0_304 (.A1(n_0_647), .A2(n_0_0_807), .B1(n_0_0_805), .B2(n_0_646), 
      .ZN(n_0_0_192));
   OAI22_X1 i_0_0_305 (.A1(n_0_646), .A2(n_0_0_805), .B1(n_0_0_803), .B2(n_0_645), 
      .ZN(n_0_0_193));
   AOI221_X1 i_0_0_306 (.A(n_0_0_195), .B1(n_0_0_801), .B2(n_0_644), .C1(n_0_645), 
      .C2(n_0_0_803), .ZN(n_0_0_194));
   AOI21_X1 i_0_0_307 (.A(n_0_0_196), .B1(n_0_0_198), .B2(n_0_0_197), .ZN(
      n_0_0_195));
   OAI22_X1 i_0_0_308 (.A1(n_0_644), .A2(n_0_0_801), .B1(n_0_0_799), .B2(n_0_643), 
      .ZN(n_0_0_196));
   AOI22_X1 i_0_0_309 (.A1(n_0_643), .A2(n_0_0_799), .B1(n_0_0_797), .B2(n_0_642), 
      .ZN(n_0_0_197));
   OAI22_X1 i_0_0_310 (.A1(n_0_642), .A2(n_0_0_797), .B1(n_0_0_203), .B2(
      n_0_0_199), .ZN(n_0_0_198));
   AOI21_X1 i_0_0_311 (.A(n_0_0_200), .B1(n_0_0_202), .B2(n_0_0_201), .ZN(
      n_0_0_199));
   OAI22_X1 i_0_0_312 (.A1(n_0_641), .A2(n_0_0_795), .B1(n_0_0_793), .B2(n_0_640), 
      .ZN(n_0_0_200));
   AOI22_X1 i_0_0_313 (.A1(n_0_640), .A2(n_0_0_793), .B1(n_0_0_791), .B2(n_0_639), 
      .ZN(n_0_0_201));
   OAI22_X1 i_0_0_314 (.A1(n_0_0_861), .A2(n_0_70), .B1(n_0_0_791), .B2(n_0_639), 
      .ZN(n_0_0_202));
   INV_X1 i_0_0_315 (.A(n_0_0_204), .ZN(n_0_0_203));
   NAND2_X1 i_0_0_316 (.A1(n_0_641), .A2(n_0_0_795), .ZN(n_0_0_204));
   NAND2_X1 i_0_0_317 (.A1(n_0_660), .A2(n_0_0_758), .ZN(n_0_0_205));
   NOR2_X1 i_0_0_318 (.A1(n_0_0_206), .A2(n_0_0_861), .ZN(n_0_617));
   NOR2_X1 i_0_0_319 (.A1(n_0_0_206), .A2(n_0_0_834), .ZN(n_0_618));
   NOR2_X1 i_0_0_320 (.A1(n_0_0_206), .A2(n_0_0_835), .ZN(n_0_619));
   NOR2_X1 i_0_0_321 (.A1(n_0_0_206), .A2(n_0_0_836), .ZN(n_0_620));
   NOR2_X1 i_0_0_322 (.A1(n_0_0_206), .A2(n_0_0_837), .ZN(n_0_621));
   NOR2_X1 i_0_0_323 (.A1(n_0_0_206), .A2(n_0_0_838), .ZN(n_0_622));
   NOR2_X1 i_0_0_324 (.A1(n_0_0_206), .A2(n_0_0_839), .ZN(n_0_623));
   NOR2_X1 i_0_0_325 (.A1(n_0_0_206), .A2(n_0_0_840), .ZN(n_0_624));
   NOR2_X1 i_0_0_326 (.A1(n_0_0_206), .A2(n_0_0_841), .ZN(n_0_625));
   NOR2_X1 i_0_0_327 (.A1(n_0_0_206), .A2(n_0_0_842), .ZN(n_0_626));
   NOR2_X1 i_0_0_328 (.A1(n_0_0_206), .A2(n_0_0_843), .ZN(n_0_627));
   NOR2_X1 i_0_0_329 (.A1(n_0_0_206), .A2(n_0_0_844), .ZN(n_0_628));
   NOR2_X1 i_0_0_330 (.A1(n_0_0_206), .A2(n_0_0_845), .ZN(n_0_629));
   NOR2_X1 i_0_0_331 (.A1(n_0_0_206), .A2(n_0_0_846), .ZN(n_0_630));
   NOR2_X1 i_0_0_332 (.A1(n_0_0_206), .A2(n_0_0_847), .ZN(n_0_631));
   NOR2_X1 i_0_0_333 (.A1(n_0_0_206), .A2(n_0_0_848), .ZN(n_0_632));
   NOR2_X1 i_0_0_334 (.A1(n_0_0_206), .A2(n_0_0_849), .ZN(n_0_633));
   NOR2_X1 i_0_0_335 (.A1(n_0_0_206), .A2(n_0_0_850), .ZN(n_0_634));
   NOR2_X1 i_0_0_336 (.A1(n_0_0_206), .A2(n_0_0_851), .ZN(n_0_635));
   NOR2_X1 i_0_0_337 (.A1(n_0_0_206), .A2(n_0_0_852), .ZN(n_0_636));
   NOR2_X1 i_0_0_338 (.A1(n_0_0_206), .A2(n_0_0_853), .ZN(n_0_637));
   NOR2_X1 i_0_0_339 (.A1(n_0_0_206), .A2(n_0_0_854), .ZN(n_0_638));
   INV_X1 i_0_0_340 (.A(n_0_0_206), .ZN(n_0_63));
   AOI21_X1 i_0_0_341 (.A(n_0_0_207), .B1(n_0_0_758), .B2(n_0_615), .ZN(
      n_0_0_206));
   AOI21_X1 i_0_0_342 (.A(n_0_0_208), .B1(n_0_0_210), .B2(n_0_0_209), .ZN(
      n_0_0_207));
   OAI22_X1 i_0_0_343 (.A1(n_0_614), .A2(n_0_0_831), .B1(n_0_0_758), .B2(n_0_615), 
      .ZN(n_0_0_208));
   AOI22_X1 i_0_0_344 (.A1(n_0_614), .A2(n_0_0_831), .B1(n_0_0_829), .B2(n_0_613), 
      .ZN(n_0_0_209));
   OAI221_X1 i_0_0_345 (.A(n_0_0_211), .B1(n_0_0_827), .B2(n_0_612), .C1(n_0_613), 
      .C2(n_0_0_829), .ZN(n_0_0_210));
   OAI21_X1 i_0_0_346 (.A(n_0_0_212), .B1(n_0_0_214), .B2(n_0_0_213), .ZN(
      n_0_0_211));
   AOI22_X1 i_0_0_347 (.A1(n_0_612), .A2(n_0_0_827), .B1(n_0_0_825), .B2(n_0_611), 
      .ZN(n_0_0_212));
   OAI22_X1 i_0_0_348 (.A1(n_0_611), .A2(n_0_0_825), .B1(n_0_0_823), .B2(n_0_610), 
      .ZN(n_0_0_213));
   AOI221_X1 i_0_0_349 (.A(n_0_0_215), .B1(n_0_0_821), .B2(n_0_609), .C1(n_0_610), 
      .C2(n_0_0_823), .ZN(n_0_0_214));
   AOI21_X1 i_0_0_350 (.A(n_0_0_216), .B1(n_0_0_218), .B2(n_0_0_217), .ZN(
      n_0_0_215));
   OAI22_X1 i_0_0_351 (.A1(n_0_609), .A2(n_0_0_821), .B1(n_0_0_819), .B2(n_0_608), 
      .ZN(n_0_0_216));
   AOI22_X1 i_0_0_352 (.A1(n_0_607), .A2(n_0_0_817), .B1(n_0_0_819), .B2(n_0_608), 
      .ZN(n_0_0_217));
   OAI221_X1 i_0_0_353 (.A(n_0_0_219), .B1(n_0_0_815), .B2(n_0_606), .C1(n_0_607), 
      .C2(n_0_0_817), .ZN(n_0_0_218));
   OAI21_X1 i_0_0_354 (.A(n_0_0_220), .B1(n_0_0_222), .B2(n_0_0_221), .ZN(
      n_0_0_219));
   AOI22_X1 i_0_0_355 (.A1(n_0_606), .A2(n_0_0_815), .B1(n_0_0_813), .B2(n_0_605), 
      .ZN(n_0_0_220));
   OAI22_X1 i_0_0_356 (.A1(n_0_605), .A2(n_0_0_813), .B1(n_0_0_811), .B2(n_0_604), 
      .ZN(n_0_0_221));
   AOI221_X1 i_0_0_357 (.A(n_0_0_223), .B1(n_0_0_809), .B2(n_0_603), .C1(n_0_604), 
      .C2(n_0_0_811), .ZN(n_0_0_222));
   NOR2_X1 i_0_0_358 (.A1(n_0_0_225), .A2(n_0_0_224), .ZN(n_0_0_223));
   OAI22_X1 i_0_0_359 (.A1(n_0_603), .A2(n_0_0_809), .B1(n_0_0_807), .B2(n_0_602), 
      .ZN(n_0_0_224));
   AOI221_X1 i_0_0_360 (.A(n_0_0_226), .B1(n_0_0_805), .B2(n_0_601), .C1(n_0_602), 
      .C2(n_0_0_807), .ZN(n_0_0_225));
   AOI21_X1 i_0_0_361 (.A(n_0_0_227), .B1(n_0_0_229), .B2(n_0_0_228), .ZN(
      n_0_0_226));
   OAI22_X1 i_0_0_362 (.A1(n_0_601), .A2(n_0_0_805), .B1(n_0_0_803), .B2(n_0_600), 
      .ZN(n_0_0_227));
   AOI22_X1 i_0_0_363 (.A1(n_0_600), .A2(n_0_0_803), .B1(n_0_0_801), .B2(n_0_599), 
      .ZN(n_0_0_228));
   OAI221_X1 i_0_0_364 (.A(n_0_0_230), .B1(n_0_0_799), .B2(n_0_598), .C1(n_0_599), 
      .C2(n_0_0_801), .ZN(n_0_0_229));
   OAI21_X1 i_0_0_365 (.A(n_0_0_231), .B1(n_0_0_233), .B2(n_0_0_232), .ZN(
      n_0_0_230));
   AOI22_X1 i_0_0_366 (.A1(n_0_598), .A2(n_0_0_799), .B1(n_0_0_797), .B2(n_0_597), 
      .ZN(n_0_0_231));
   OAI22_X1 i_0_0_367 (.A1(n_0_597), .A2(n_0_0_797), .B1(n_0_0_795), .B2(n_0_596), 
      .ZN(n_0_0_232));
   AOI21_X1 i_0_0_368 (.A(n_0_0_234), .B1(n_0_0_795), .B2(n_0_596), .ZN(
      n_0_0_233));
   AOI21_X1 i_0_0_369 (.A(n_0_0_237), .B1(n_0_0_236), .B2(n_0_0_235), .ZN(
      n_0_0_234));
   AOI22_X1 i_0_0_370 (.A1(n_0_595), .A2(n_0_0_793), .B1(n_0_0_791), .B2(n_0_594), 
      .ZN(n_0_0_235));
   OAI22_X1 i_0_0_371 (.A1(n_0_0_861), .A2(n_0_71), .B1(n_0_0_791), .B2(n_0_594), 
      .ZN(n_0_0_236));
   NOR2_X1 i_0_0_372 (.A1(n_0_595), .A2(n_0_0_793), .ZN(n_0_0_237));
   NOR2_X1 i_0_0_373 (.A1(n_0_0_238), .A2(n_0_0_861), .ZN(n_0_572));
   NOR2_X1 i_0_0_374 (.A1(n_0_0_238), .A2(n_0_0_834), .ZN(n_0_573));
   NOR2_X1 i_0_0_375 (.A1(n_0_0_238), .A2(n_0_0_835), .ZN(n_0_574));
   NOR2_X1 i_0_0_376 (.A1(n_0_0_238), .A2(n_0_0_836), .ZN(n_0_575));
   NOR2_X1 i_0_0_377 (.A1(n_0_0_238), .A2(n_0_0_837), .ZN(n_0_576));
   NOR2_X1 i_0_0_378 (.A1(n_0_0_238), .A2(n_0_0_838), .ZN(n_0_577));
   NOR2_X1 i_0_0_379 (.A1(n_0_0_238), .A2(n_0_0_839), .ZN(n_0_578));
   NOR2_X1 i_0_0_380 (.A1(n_0_0_238), .A2(n_0_0_840), .ZN(n_0_579));
   NOR2_X1 i_0_0_381 (.A1(n_0_0_238), .A2(n_0_0_841), .ZN(n_0_580));
   NOR2_X1 i_0_0_382 (.A1(n_0_0_238), .A2(n_0_0_842), .ZN(n_0_581));
   NOR2_X1 i_0_0_383 (.A1(n_0_0_238), .A2(n_0_0_843), .ZN(n_0_582));
   NOR2_X1 i_0_0_384 (.A1(n_0_0_238), .A2(n_0_0_844), .ZN(n_0_583));
   NOR2_X1 i_0_0_385 (.A1(n_0_0_238), .A2(n_0_0_845), .ZN(n_0_584));
   NOR2_X1 i_0_0_386 (.A1(n_0_0_238), .A2(n_0_0_846), .ZN(n_0_585));
   NOR2_X1 i_0_0_387 (.A1(n_0_0_238), .A2(n_0_0_847), .ZN(n_0_586));
   NOR2_X1 i_0_0_388 (.A1(n_0_0_238), .A2(n_0_0_848), .ZN(n_0_587));
   NOR2_X1 i_0_0_389 (.A1(n_0_0_238), .A2(n_0_0_849), .ZN(n_0_588));
   NOR2_X1 i_0_0_390 (.A1(n_0_0_238), .A2(n_0_0_850), .ZN(n_0_589));
   NOR2_X1 i_0_0_391 (.A1(n_0_0_238), .A2(n_0_0_851), .ZN(n_0_590));
   NOR2_X1 i_0_0_392 (.A1(n_0_0_238), .A2(n_0_0_852), .ZN(n_0_591));
   NOR2_X1 i_0_0_393 (.A1(n_0_0_238), .A2(n_0_0_853), .ZN(n_0_592));
   NOR2_X1 i_0_0_394 (.A1(n_0_0_238), .A2(n_0_0_854), .ZN(n_0_593));
   INV_X1 i_0_0_395 (.A(n_0_64), .ZN(n_0_0_238));
   OAI21_X1 i_0_0_396 (.A(n_0_0_269), .B1(n_0_0_240), .B2(n_0_0_239), .ZN(n_0_64));
   OAI22_X1 i_0_0_397 (.A1(n_0_569), .A2(n_0_0_831), .B1(n_0_0_758), .B2(n_0_570), 
      .ZN(n_0_0_239));
   AOI221_X1 i_0_0_398 (.A(n_0_0_241), .B1(n_0_0_829), .B2(n_0_568), .C1(n_0_569), 
      .C2(n_0_0_831), .ZN(n_0_0_240));
   AOI21_X1 i_0_0_399 (.A(n_0_0_242), .B1(n_0_0_244), .B2(n_0_0_243), .ZN(
      n_0_0_241));
   OAI22_X1 i_0_0_400 (.A1(n_0_568), .A2(n_0_0_829), .B1(n_0_0_827), .B2(n_0_567), 
      .ZN(n_0_0_242));
   AOI22_X1 i_0_0_401 (.A1(n_0_567), .A2(n_0_0_827), .B1(n_0_0_825), .B2(n_0_566), 
      .ZN(n_0_0_243));
   OAI221_X1 i_0_0_402 (.A(n_0_0_245), .B1(n_0_0_823), .B2(n_0_565), .C1(n_0_566), 
      .C2(n_0_0_825), .ZN(n_0_0_244));
   OAI21_X1 i_0_0_403 (.A(n_0_0_246), .B1(n_0_0_248), .B2(n_0_0_247), .ZN(
      n_0_0_245));
   AOI22_X1 i_0_0_404 (.A1(n_0_565), .A2(n_0_0_823), .B1(n_0_0_821), .B2(n_0_564), 
      .ZN(n_0_0_246));
   OAI22_X1 i_0_0_405 (.A1(n_0_564), .A2(n_0_0_821), .B1(n_0_0_819), .B2(n_0_563), 
      .ZN(n_0_0_247));
   AOI221_X1 i_0_0_406 (.A(n_0_0_249), .B1(n_0_0_817), .B2(n_0_562), .C1(n_0_563), 
      .C2(n_0_0_819), .ZN(n_0_0_248));
   AOI21_X1 i_0_0_407 (.A(n_0_0_250), .B1(n_0_0_252), .B2(n_0_0_251), .ZN(
      n_0_0_249));
   OAI22_X1 i_0_0_408 (.A1(n_0_562), .A2(n_0_0_817), .B1(n_0_0_815), .B2(n_0_561), 
      .ZN(n_0_0_250));
   AOI22_X1 i_0_0_409 (.A1(n_0_561), .A2(n_0_0_815), .B1(n_0_0_813), .B2(n_0_560), 
      .ZN(n_0_0_251));
   OAI221_X1 i_0_0_410 (.A(n_0_0_253), .B1(n_0_0_811), .B2(n_0_559), .C1(n_0_560), 
      .C2(n_0_0_813), .ZN(n_0_0_252));
   OAI21_X1 i_0_0_411 (.A(n_0_0_254), .B1(n_0_0_256), .B2(n_0_0_255), .ZN(
      n_0_0_253));
   AOI22_X1 i_0_0_412 (.A1(n_0_559), .A2(n_0_0_811), .B1(n_0_0_809), .B2(n_0_558), 
      .ZN(n_0_0_254));
   OAI22_X1 i_0_0_413 (.A1(n_0_558), .A2(n_0_0_809), .B1(n_0_0_807), .B2(n_0_557), 
      .ZN(n_0_0_255));
   AOI221_X1 i_0_0_414 (.A(n_0_0_257), .B1(n_0_0_805), .B2(n_0_556), .C1(n_0_557), 
      .C2(n_0_0_807), .ZN(n_0_0_256));
   AOI21_X1 i_0_0_415 (.A(n_0_0_258), .B1(n_0_0_260), .B2(n_0_0_259), .ZN(
      n_0_0_257));
   OAI22_X1 i_0_0_416 (.A1(n_0_556), .A2(n_0_0_805), .B1(n_0_0_803), .B2(n_0_555), 
      .ZN(n_0_0_258));
   AOI22_X1 i_0_0_417 (.A1(n_0_555), .A2(n_0_0_803), .B1(n_0_0_801), .B2(n_0_554), 
      .ZN(n_0_0_259));
   OAI221_X1 i_0_0_418 (.A(n_0_0_261), .B1(n_0_0_799), .B2(n_0_553), .C1(n_0_554), 
      .C2(n_0_0_801), .ZN(n_0_0_260));
   OAI21_X1 i_0_0_419 (.A(n_0_0_262), .B1(n_0_0_263), .B2(n_0_0_264), .ZN(
      n_0_0_261));
   AOI22_X1 i_0_0_420 (.A1(n_0_553), .A2(n_0_0_799), .B1(n_0_0_797), .B2(n_0_552), 
      .ZN(n_0_0_262));
   NOR2_X1 i_0_0_421 (.A1(n_0_552), .A2(n_0_0_797), .ZN(n_0_0_263));
   AOI21_X1 i_0_0_422 (.A(n_0_0_265), .B1(n_0_0_795), .B2(n_0_551), .ZN(
      n_0_0_264));
   AOI21_X1 i_0_0_423 (.A(n_0_0_266), .B1(n_0_0_268), .B2(n_0_0_267), .ZN(
      n_0_0_265));
   OAI22_X1 i_0_0_424 (.A1(n_0_551), .A2(n_0_0_795), .B1(n_0_0_793), .B2(n_0_550), 
      .ZN(n_0_0_266));
   AOI22_X1 i_0_0_425 (.A1(n_0_550), .A2(n_0_0_793), .B1(n_0_0_791), .B2(n_0_549), 
      .ZN(n_0_0_267));
   OAI22_X1 i_0_0_426 (.A1(n_0_72), .A2(n_0_0_861), .B1(n_0_549), .B2(n_0_0_791), 
      .ZN(n_0_0_268));
   NAND2_X1 i_0_0_427 (.A1(n_0_570), .A2(n_0_0_758), .ZN(n_0_0_269));
   NOR2_X1 i_0_0_428 (.A1(n_0_0_270), .A2(n_0_0_861), .ZN(n_0_527));
   NOR2_X1 i_0_0_429 (.A1(n_0_0_270), .A2(n_0_0_834), .ZN(n_0_528));
   NOR2_X1 i_0_0_430 (.A1(n_0_0_270), .A2(n_0_0_835), .ZN(n_0_529));
   NOR2_X1 i_0_0_431 (.A1(n_0_0_270), .A2(n_0_0_836), .ZN(n_0_530));
   NOR2_X1 i_0_0_432 (.A1(n_0_0_270), .A2(n_0_0_837), .ZN(n_0_531));
   NOR2_X1 i_0_0_433 (.A1(n_0_0_270), .A2(n_0_0_838), .ZN(n_0_532));
   NOR2_X1 i_0_0_434 (.A1(n_0_0_270), .A2(n_0_0_839), .ZN(n_0_533));
   NOR2_X1 i_0_0_435 (.A1(n_0_0_270), .A2(n_0_0_840), .ZN(n_0_534));
   NOR2_X1 i_0_0_436 (.A1(n_0_0_270), .A2(n_0_0_841), .ZN(n_0_535));
   NOR2_X1 i_0_0_437 (.A1(n_0_0_270), .A2(n_0_0_842), .ZN(n_0_536));
   NOR2_X1 i_0_0_438 (.A1(n_0_0_270), .A2(n_0_0_843), .ZN(n_0_537));
   NOR2_X1 i_0_0_439 (.A1(n_0_0_270), .A2(n_0_0_844), .ZN(n_0_538));
   NOR2_X1 i_0_0_440 (.A1(n_0_0_270), .A2(n_0_0_845), .ZN(n_0_539));
   NOR2_X1 i_0_0_441 (.A1(n_0_0_270), .A2(n_0_0_846), .ZN(n_0_540));
   NOR2_X1 i_0_0_442 (.A1(n_0_0_270), .A2(n_0_0_847), .ZN(n_0_541));
   NOR2_X1 i_0_0_443 (.A1(n_0_0_270), .A2(n_0_0_848), .ZN(n_0_542));
   NOR2_X1 i_0_0_444 (.A1(n_0_0_270), .A2(n_0_0_849), .ZN(n_0_543));
   NOR2_X1 i_0_0_445 (.A1(n_0_0_270), .A2(n_0_0_850), .ZN(n_0_544));
   NOR2_X1 i_0_0_446 (.A1(n_0_0_270), .A2(n_0_0_851), .ZN(n_0_545));
   NOR2_X1 i_0_0_447 (.A1(n_0_0_270), .A2(n_0_0_852), .ZN(n_0_546));
   NOR2_X1 i_0_0_448 (.A1(n_0_0_270), .A2(n_0_0_853), .ZN(n_0_547));
   NOR2_X1 i_0_0_449 (.A1(n_0_0_270), .A2(n_0_0_854), .ZN(n_0_548));
   INV_X1 i_0_0_450 (.A(n_0_0_270), .ZN(n_0_65));
   AOI22_X1 i_0_0_451 (.A1(n_0_0_273), .A2(n_0_0_271), .B1(n_0_525), .B2(
      n_0_0_758), .ZN(n_0_0_270));
   INV_X1 i_0_0_452 (.A(n_0_0_272), .ZN(n_0_0_271));
   OAI22_X1 i_0_0_453 (.A1(n_0_524), .A2(n_0_0_831), .B1(n_0_0_758), .B2(n_0_525), 
      .ZN(n_0_0_272));
   OAI21_X1 i_0_0_454 (.A(n_0_0_274), .B1(n_0_0_276), .B2(n_0_0_275), .ZN(
      n_0_0_273));
   AOI22_X1 i_0_0_455 (.A1(n_0_524), .A2(n_0_0_831), .B1(n_0_0_829), .B2(n_0_523), 
      .ZN(n_0_0_274));
   OAI22_X1 i_0_0_456 (.A1(n_0_523), .A2(n_0_0_829), .B1(n_0_0_827), .B2(n_0_522), 
      .ZN(n_0_0_275));
   AOI221_X1 i_0_0_457 (.A(n_0_0_277), .B1(n_0_0_825), .B2(n_0_521), .C1(n_0_522), 
      .C2(n_0_0_827), .ZN(n_0_0_276));
   AOI21_X1 i_0_0_458 (.A(n_0_0_278), .B1(n_0_0_280), .B2(n_0_0_279), .ZN(
      n_0_0_277));
   OAI22_X1 i_0_0_459 (.A1(n_0_521), .A2(n_0_0_825), .B1(n_0_0_823), .B2(n_0_520), 
      .ZN(n_0_0_278));
   AOI22_X1 i_0_0_460 (.A1(n_0_520), .A2(n_0_0_823), .B1(n_0_0_821), .B2(n_0_519), 
      .ZN(n_0_0_279));
   OAI221_X1 i_0_0_461 (.A(n_0_0_281), .B1(n_0_0_819), .B2(n_0_518), .C1(n_0_519), 
      .C2(n_0_0_821), .ZN(n_0_0_280));
   OAI21_X1 i_0_0_462 (.A(n_0_0_282), .B1(n_0_0_284), .B2(n_0_0_283), .ZN(
      n_0_0_281));
   AOI22_X1 i_0_0_463 (.A1(n_0_517), .A2(n_0_0_817), .B1(n_0_0_819), .B2(n_0_518), 
      .ZN(n_0_0_282));
   OAI22_X1 i_0_0_464 (.A1(n_0_517), .A2(n_0_0_817), .B1(n_0_0_815), .B2(n_0_516), 
      .ZN(n_0_0_283));
   AOI221_X1 i_0_0_465 (.A(n_0_0_285), .B1(n_0_0_813), .B2(n_0_515), .C1(n_0_516), 
      .C2(n_0_0_815), .ZN(n_0_0_284));
   AOI21_X1 i_0_0_466 (.A(n_0_0_286), .B1(n_0_0_288), .B2(n_0_0_287), .ZN(
      n_0_0_285));
   OAI22_X1 i_0_0_467 (.A1(n_0_515), .A2(n_0_0_813), .B1(n_0_0_811), .B2(n_0_514), 
      .ZN(n_0_0_286));
   AOI22_X1 i_0_0_468 (.A1(n_0_514), .A2(n_0_0_811), .B1(n_0_0_809), .B2(n_0_513), 
      .ZN(n_0_0_287));
   OAI221_X1 i_0_0_469 (.A(n_0_0_289), .B1(n_0_0_807), .B2(n_0_512), .C1(n_0_513), 
      .C2(n_0_0_809), .ZN(n_0_0_288));
   OAI21_X1 i_0_0_470 (.A(n_0_0_290), .B1(n_0_0_292), .B2(n_0_0_291), .ZN(
      n_0_0_289));
   AOI22_X1 i_0_0_471 (.A1(n_0_512), .A2(n_0_0_807), .B1(n_0_0_805), .B2(n_0_511), 
      .ZN(n_0_0_290));
   OAI22_X1 i_0_0_472 (.A1(n_0_511), .A2(n_0_0_805), .B1(n_0_0_803), .B2(n_0_510), 
      .ZN(n_0_0_291));
   AOI221_X1 i_0_0_473 (.A(n_0_0_293), .B1(n_0_0_801), .B2(n_0_509), .C1(n_0_510), 
      .C2(n_0_0_803), .ZN(n_0_0_292));
   AOI21_X1 i_0_0_474 (.A(n_0_0_294), .B1(n_0_0_296), .B2(n_0_0_295), .ZN(
      n_0_0_293));
   OAI22_X1 i_0_0_475 (.A1(n_0_509), .A2(n_0_0_801), .B1(n_0_0_799), .B2(n_0_508), 
      .ZN(n_0_0_294));
   AOI22_X1 i_0_0_476 (.A1(n_0_508), .A2(n_0_0_799), .B1(n_0_0_797), .B2(n_0_507), 
      .ZN(n_0_0_295));
   OAI21_X1 i_0_0_477 (.A(n_0_0_297), .B1(n_0_0_797), .B2(n_0_507), .ZN(
      n_0_0_296));
   OAI21_X1 i_0_0_478 (.A(n_0_0_302), .B1(n_0_0_299), .B2(n_0_0_298), .ZN(
      n_0_0_297));
   OAI22_X1 i_0_0_479 (.A1(n_0_506), .A2(n_0_0_795), .B1(n_0_0_793), .B2(n_0_505), 
      .ZN(n_0_0_298));
   AOI221_X1 i_0_0_480 (.A(n_0_0_300), .B1(n_0_0_791), .B2(n_0_504), .C1(n_0_505), 
      .C2(n_0_0_793), .ZN(n_0_0_299));
   AOI21_X1 i_0_0_481 (.A(n_0_0_301), .B1(n_0_0_760), .B2(in_b[0]), .ZN(
      n_0_0_300));
   NOR2_X1 i_0_0_482 (.A1(n_0_504), .A2(n_0_0_791), .ZN(n_0_0_301));
   NAND2_X1 i_0_0_483 (.A1(n_0_506), .A2(n_0_0_795), .ZN(n_0_0_302));
   AND2_X1 i_0_0_484 (.A1(n_0_66), .A2(in_b[0]), .ZN(n_0_482));
   AND2_X1 i_0_0_485 (.A1(n_0_66), .A2(n_0_78), .ZN(n_0_483));
   AND2_X1 i_0_0_486 (.A1(n_0_66), .A2(n_0_79), .ZN(n_0_484));
   AND2_X1 i_0_0_487 (.A1(n_0_66), .A2(n_0_80), .ZN(n_0_485));
   AND2_X1 i_0_0_488 (.A1(n_0_66), .A2(n_0_81), .ZN(n_0_486));
   AND2_X1 i_0_0_489 (.A1(n_0_66), .A2(n_0_82), .ZN(n_0_487));
   AND2_X1 i_0_0_490 (.A1(n_0_66), .A2(n_0_83), .ZN(n_0_488));
   AND2_X1 i_0_0_491 (.A1(n_0_66), .A2(n_0_84), .ZN(n_0_489));
   AND2_X1 i_0_0_492 (.A1(n_0_66), .A2(n_0_85), .ZN(n_0_490));
   AND2_X1 i_0_0_493 (.A1(n_0_66), .A2(n_0_86), .ZN(n_0_491));
   AND2_X1 i_0_0_494 (.A1(n_0_66), .A2(n_0_87), .ZN(n_0_492));
   AND2_X1 i_0_0_495 (.A1(n_0_66), .A2(n_0_88), .ZN(n_0_493));
   AND2_X1 i_0_0_496 (.A1(n_0_66), .A2(n_0_89), .ZN(n_0_494));
   AND2_X1 i_0_0_497 (.A1(n_0_66), .A2(n_0_90), .ZN(n_0_495));
   AND2_X1 i_0_0_498 (.A1(n_0_66), .A2(n_0_91), .ZN(n_0_496));
   AND2_X1 i_0_0_499 (.A1(n_0_66), .A2(n_0_92), .ZN(n_0_497));
   AND2_X1 i_0_0_500 (.A1(n_0_66), .A2(n_0_93), .ZN(n_0_498));
   AND2_X1 i_0_0_501 (.A1(n_0_66), .A2(n_0_94), .ZN(n_0_499));
   AND2_X1 i_0_0_502 (.A1(n_0_66), .A2(n_0_95), .ZN(n_0_500));
   AND2_X1 i_0_0_503 (.A1(n_0_66), .A2(n_0_96), .ZN(n_0_501));
   AND2_X1 i_0_0_504 (.A1(n_0_66), .A2(n_0_97), .ZN(n_0_502));
   AND2_X1 i_0_0_505 (.A1(n_0_66), .A2(n_0_98), .ZN(n_0_503));
   NAND2_X1 i_0_0_506 (.A1(n_0_0_335), .A2(n_0_0_303), .ZN(n_0_66));
   OAI221_X1 i_0_0_507 (.A(n_0_0_304), .B1(n_0_0_831), .B2(n_0_479), .C1(n_0_480), 
      .C2(n_0_0_758), .ZN(n_0_0_303));
   NAND2_X1 i_0_0_508 (.A1(n_0_0_306), .A2(n_0_0_305), .ZN(n_0_0_304));
   AOI22_X1 i_0_0_509 (.A1(n_0_479), .A2(n_0_0_831), .B1(n_0_0_829), .B2(n_0_478), 
      .ZN(n_0_0_305));
   OAI221_X1 i_0_0_510 (.A(n_0_0_307), .B1(n_0_0_827), .B2(n_0_477), .C1(n_0_478), 
      .C2(n_0_0_829), .ZN(n_0_0_306));
   NAND2_X1 i_0_0_511 (.A1(n_0_0_309), .A2(n_0_0_308), .ZN(n_0_0_307));
   AOI22_X1 i_0_0_512 (.A1(n_0_477), .A2(n_0_0_827), .B1(n_0_0_825), .B2(n_0_476), 
      .ZN(n_0_0_308));
   OAI221_X1 i_0_0_513 (.A(n_0_0_310), .B1(n_0_0_823), .B2(n_0_475), .C1(n_0_476), 
      .C2(n_0_0_825), .ZN(n_0_0_309));
   OAI21_X1 i_0_0_514 (.A(n_0_0_311), .B1(n_0_0_313), .B2(n_0_0_312), .ZN(
      n_0_0_310));
   AOI22_X1 i_0_0_515 (.A1(n_0_475), .A2(n_0_0_823), .B1(n_0_0_821), .B2(n_0_474), 
      .ZN(n_0_0_311));
   OAI22_X1 i_0_0_516 (.A1(n_0_474), .A2(n_0_0_821), .B1(n_0_0_819), .B2(n_0_473), 
      .ZN(n_0_0_312));
   AOI221_X1 i_0_0_517 (.A(n_0_0_314), .B1(n_0_0_817), .B2(n_0_472), .C1(n_0_473), 
      .C2(n_0_0_819), .ZN(n_0_0_313));
   AOI21_X1 i_0_0_518 (.A(n_0_0_315), .B1(n_0_0_317), .B2(n_0_0_316), .ZN(
      n_0_0_314));
   OAI22_X1 i_0_0_519 (.A1(n_0_472), .A2(n_0_0_817), .B1(n_0_0_815), .B2(n_0_471), 
      .ZN(n_0_0_315));
   AOI22_X1 i_0_0_520 (.A1(n_0_471), .A2(n_0_0_815), .B1(n_0_0_813), .B2(n_0_470), 
      .ZN(n_0_0_316));
   OAI221_X1 i_0_0_521 (.A(n_0_0_318), .B1(n_0_0_811), .B2(n_0_469), .C1(n_0_470), 
      .C2(n_0_0_813), .ZN(n_0_0_317));
   NAND2_X1 i_0_0_522 (.A1(n_0_0_320), .A2(n_0_0_319), .ZN(n_0_0_318));
   AOI22_X1 i_0_0_523 (.A1(n_0_469), .A2(n_0_0_811), .B1(n_0_0_809), .B2(n_0_468), 
      .ZN(n_0_0_319));
   OAI221_X1 i_0_0_524 (.A(n_0_0_321), .B1(n_0_0_807), .B2(n_0_467), .C1(n_0_468), 
      .C2(n_0_0_809), .ZN(n_0_0_320));
   OAI21_X1 i_0_0_525 (.A(n_0_0_322), .B1(n_0_0_324), .B2(n_0_0_323), .ZN(
      n_0_0_321));
   AOI22_X1 i_0_0_526 (.A1(n_0_467), .A2(n_0_0_807), .B1(n_0_0_805), .B2(n_0_466), 
      .ZN(n_0_0_322));
   OAI22_X1 i_0_0_527 (.A1(n_0_466), .A2(n_0_0_805), .B1(n_0_0_803), .B2(n_0_465), 
      .ZN(n_0_0_323));
   AOI221_X1 i_0_0_528 (.A(n_0_0_325), .B1(n_0_0_801), .B2(n_0_464), .C1(n_0_465), 
      .C2(n_0_0_803), .ZN(n_0_0_324));
   AOI21_X1 i_0_0_529 (.A(n_0_0_326), .B1(n_0_0_328), .B2(n_0_0_327), .ZN(
      n_0_0_325));
   OAI22_X1 i_0_0_530 (.A1(n_0_464), .A2(n_0_0_801), .B1(n_0_0_799), .B2(n_0_463), 
      .ZN(n_0_0_326));
   AOI22_X1 i_0_0_531 (.A1(n_0_463), .A2(n_0_0_799), .B1(n_0_0_797), .B2(n_0_462), 
      .ZN(n_0_0_327));
   OAI21_X1 i_0_0_532 (.A(n_0_0_329), .B1(n_0_0_797), .B2(n_0_462), .ZN(
      n_0_0_328));
   OAI21_X1 i_0_0_533 (.A(n_0_0_334), .B1(n_0_0_331), .B2(n_0_0_330), .ZN(
      n_0_0_329));
   OAI22_X1 i_0_0_534 (.A1(n_0_461), .A2(n_0_0_795), .B1(n_0_0_793), .B2(n_0_460), 
      .ZN(n_0_0_330));
   AOI221_X1 i_0_0_535 (.A(n_0_0_332), .B1(n_0_0_791), .B2(n_0_459), .C1(n_0_460), 
      .C2(n_0_0_793), .ZN(n_0_0_331));
   AOI21_X1 i_0_0_536 (.A(n_0_0_333), .B1(n_0_0_761), .B2(in_b[0]), .ZN(
      n_0_0_332));
   NOR2_X1 i_0_0_537 (.A1(n_0_459), .A2(n_0_0_791), .ZN(n_0_0_333));
   NAND2_X1 i_0_0_538 (.A1(n_0_461), .A2(n_0_0_795), .ZN(n_0_0_334));
   NAND2_X1 i_0_0_539 (.A1(n_0_480), .A2(n_0_0_758), .ZN(n_0_0_335));
   NOR3_X1 i_0_0_540 (.A1(n_0_0_336), .A2(n_0_0_861), .A3(n_0_0_338), .ZN(
      n_0_437));
   NOR3_X1 i_0_0_541 (.A1(n_0_0_336), .A2(n_0_0_834), .A3(n_0_0_338), .ZN(
      n_0_438));
   NOR3_X1 i_0_0_542 (.A1(n_0_0_336), .A2(n_0_0_835), .A3(n_0_0_338), .ZN(
      n_0_439));
   NOR3_X1 i_0_0_543 (.A1(n_0_0_336), .A2(n_0_0_836), .A3(n_0_0_338), .ZN(
      n_0_440));
   NOR3_X1 i_0_0_544 (.A1(n_0_0_336), .A2(n_0_0_837), .A3(n_0_0_338), .ZN(
      n_0_441));
   NOR3_X1 i_0_0_545 (.A1(n_0_0_336), .A2(n_0_0_838), .A3(n_0_0_338), .ZN(
      n_0_442));
   NOR3_X1 i_0_0_546 (.A1(n_0_0_336), .A2(n_0_0_839), .A3(n_0_0_338), .ZN(
      n_0_443));
   NOR3_X1 i_0_0_547 (.A1(n_0_0_336), .A2(n_0_0_840), .A3(n_0_0_338), .ZN(
      n_0_444));
   NOR3_X1 i_0_0_548 (.A1(n_0_0_336), .A2(n_0_0_841), .A3(n_0_0_338), .ZN(
      n_0_445));
   NOR3_X1 i_0_0_549 (.A1(n_0_0_336), .A2(n_0_0_842), .A3(n_0_0_338), .ZN(
      n_0_446));
   NOR3_X1 i_0_0_550 (.A1(n_0_0_336), .A2(n_0_0_843), .A3(n_0_0_338), .ZN(
      n_0_447));
   NOR3_X1 i_0_0_551 (.A1(n_0_0_336), .A2(n_0_0_844), .A3(n_0_0_338), .ZN(
      n_0_448));
   NOR3_X1 i_0_0_552 (.A1(n_0_0_336), .A2(n_0_0_845), .A3(n_0_0_338), .ZN(
      n_0_449));
   NOR3_X1 i_0_0_553 (.A1(n_0_0_336), .A2(n_0_0_846), .A3(n_0_0_338), .ZN(
      n_0_450));
   NOR3_X1 i_0_0_554 (.A1(n_0_0_336), .A2(n_0_0_847), .A3(n_0_0_338), .ZN(
      n_0_451));
   NOR3_X1 i_0_0_555 (.A1(n_0_0_336), .A2(n_0_0_848), .A3(n_0_0_338), .ZN(
      n_0_452));
   NOR3_X1 i_0_0_556 (.A1(n_0_0_336), .A2(n_0_0_849), .A3(n_0_0_338), .ZN(
      n_0_453));
   NOR3_X1 i_0_0_557 (.A1(n_0_0_336), .A2(n_0_0_850), .A3(n_0_0_338), .ZN(
      n_0_454));
   NOR3_X1 i_0_0_558 (.A1(n_0_0_336), .A2(n_0_0_851), .A3(n_0_0_338), .ZN(
      n_0_455));
   NOR3_X1 i_0_0_559 (.A1(n_0_0_336), .A2(n_0_0_852), .A3(n_0_0_338), .ZN(
      n_0_456));
   NOR3_X1 i_0_0_560 (.A1(n_0_0_336), .A2(n_0_0_853), .A3(n_0_0_338), .ZN(
      n_0_457));
   NOR3_X1 i_0_0_561 (.A1(n_0_0_336), .A2(n_0_0_854), .A3(n_0_0_338), .ZN(
      n_0_458));
   NOR2_X1 i_0_0_562 (.A1(n_0_0_338), .A2(n_0_0_336), .ZN(n_0_67));
   AOI22_X1 i_0_0_563 (.A1(n_0_0_339), .A2(n_0_0_337), .B1(n_0_435), .B2(
      n_0_0_758), .ZN(n_0_0_336));
   OR2_X1 i_0_0_564 (.A1(n_0_434), .A2(n_0_0_831), .ZN(n_0_0_337));
   NOR2_X1 i_0_0_565 (.A1(n_0_435), .A2(n_0_0_758), .ZN(n_0_0_338));
   OAI21_X1 i_0_0_566 (.A(n_0_0_340), .B1(n_0_0_342), .B2(n_0_0_341), .ZN(
      n_0_0_339));
   AOI22_X1 i_0_0_567 (.A1(n_0_434), .A2(n_0_0_831), .B1(n_0_0_829), .B2(n_0_433), 
      .ZN(n_0_0_340));
   OAI22_X1 i_0_0_568 (.A1(n_0_433), .A2(n_0_0_829), .B1(n_0_0_827), .B2(n_0_432), 
      .ZN(n_0_0_341));
   AOI221_X1 i_0_0_569 (.A(n_0_0_343), .B1(n_0_0_825), .B2(n_0_431), .C1(n_0_432), 
      .C2(n_0_0_827), .ZN(n_0_0_342));
   AOI21_X1 i_0_0_570 (.A(n_0_0_344), .B1(n_0_0_346), .B2(n_0_0_345), .ZN(
      n_0_0_343));
   OAI22_X1 i_0_0_571 (.A1(n_0_431), .A2(n_0_0_825), .B1(n_0_0_823), .B2(n_0_430), 
      .ZN(n_0_0_344));
   AOI22_X1 i_0_0_572 (.A1(n_0_430), .A2(n_0_0_823), .B1(n_0_0_821), .B2(n_0_429), 
      .ZN(n_0_0_345));
   OAI221_X1 i_0_0_573 (.A(n_0_0_347), .B1(n_0_0_819), .B2(n_0_428), .C1(n_0_429), 
      .C2(n_0_0_821), .ZN(n_0_0_346));
   OAI21_X1 i_0_0_574 (.A(n_0_0_348), .B1(n_0_0_350), .B2(n_0_0_349), .ZN(
      n_0_0_347));
   AOI22_X1 i_0_0_575 (.A1(n_0_427), .A2(n_0_0_817), .B1(n_0_0_819), .B2(n_0_428), 
      .ZN(n_0_0_348));
   OAI22_X1 i_0_0_576 (.A1(n_0_427), .A2(n_0_0_817), .B1(n_0_0_815), .B2(n_0_426), 
      .ZN(n_0_0_349));
   AOI221_X1 i_0_0_577 (.A(n_0_0_351), .B1(n_0_0_813), .B2(n_0_425), .C1(n_0_426), 
      .C2(n_0_0_815), .ZN(n_0_0_350));
   AOI21_X1 i_0_0_578 (.A(n_0_0_352), .B1(n_0_0_354), .B2(n_0_0_353), .ZN(
      n_0_0_351));
   OAI22_X1 i_0_0_579 (.A1(n_0_425), .A2(n_0_0_813), .B1(n_0_0_811), .B2(n_0_424), 
      .ZN(n_0_0_352));
   AOI22_X1 i_0_0_580 (.A1(n_0_424), .A2(n_0_0_811), .B1(n_0_0_809), .B2(n_0_423), 
      .ZN(n_0_0_353));
   OAI221_X1 i_0_0_581 (.A(n_0_0_355), .B1(n_0_0_807), .B2(n_0_422), .C1(n_0_423), 
      .C2(n_0_0_809), .ZN(n_0_0_354));
   OAI21_X1 i_0_0_582 (.A(n_0_0_356), .B1(n_0_0_358), .B2(n_0_0_357), .ZN(
      n_0_0_355));
   AOI22_X1 i_0_0_583 (.A1(n_0_422), .A2(n_0_0_807), .B1(n_0_0_805), .B2(n_0_421), 
      .ZN(n_0_0_356));
   OAI22_X1 i_0_0_584 (.A1(n_0_421), .A2(n_0_0_805), .B1(n_0_0_803), .B2(n_0_420), 
      .ZN(n_0_0_357));
   AOI221_X1 i_0_0_585 (.A(n_0_0_359), .B1(n_0_0_801), .B2(n_0_419), .C1(n_0_420), 
      .C2(n_0_0_803), .ZN(n_0_0_358));
   AOI21_X1 i_0_0_586 (.A(n_0_0_360), .B1(n_0_0_362), .B2(n_0_0_361), .ZN(
      n_0_0_359));
   OAI22_X1 i_0_0_587 (.A1(n_0_419), .A2(n_0_0_801), .B1(n_0_0_799), .B2(n_0_418), 
      .ZN(n_0_0_360));
   AOI22_X1 i_0_0_588 (.A1(n_0_418), .A2(n_0_0_799), .B1(n_0_0_797), .B2(n_0_417), 
      .ZN(n_0_0_361));
   OAI22_X1 i_0_0_589 (.A1(n_0_417), .A2(n_0_0_797), .B1(n_0_0_367), .B2(
      n_0_0_363), .ZN(n_0_0_362));
   AOI21_X1 i_0_0_590 (.A(n_0_0_364), .B1(n_0_0_366), .B2(n_0_0_365), .ZN(
      n_0_0_363));
   OAI22_X1 i_0_0_591 (.A1(n_0_416), .A2(n_0_0_795), .B1(n_0_0_793), .B2(n_0_415), 
      .ZN(n_0_0_364));
   AOI22_X1 i_0_0_592 (.A1(n_0_415), .A2(n_0_0_793), .B1(n_0_0_791), .B2(n_0_414), 
      .ZN(n_0_0_365));
   OAI22_X1 i_0_0_593 (.A1(n_0_0_861), .A2(n_0_75), .B1(n_0_0_791), .B2(n_0_414), 
      .ZN(n_0_0_366));
   AND2_X1 i_0_0_594 (.A1(n_0_416), .A2(n_0_0_795), .ZN(n_0_0_367));
   AND2_X1 i_0_0_595 (.A1(in_b[0]), .A2(n_0_68), .ZN(n_0_392));
   AND2_X1 i_0_0_596 (.A1(n_0_78), .A2(n_0_68), .ZN(n_0_393));
   AND2_X1 i_0_0_597 (.A1(n_0_79), .A2(n_0_68), .ZN(n_0_394));
   AND2_X1 i_0_0_598 (.A1(n_0_80), .A2(n_0_68), .ZN(n_0_395));
   AND2_X1 i_0_0_599 (.A1(n_0_81), .A2(n_0_68), .ZN(n_0_396));
   AND2_X1 i_0_0_600 (.A1(n_0_82), .A2(n_0_68), .ZN(n_0_397));
   AND2_X1 i_0_0_601 (.A1(n_0_83), .A2(n_0_68), .ZN(n_0_398));
   AND2_X1 i_0_0_602 (.A1(n_0_84), .A2(n_0_68), .ZN(n_0_399));
   AND2_X1 i_0_0_603 (.A1(n_0_85), .A2(n_0_68), .ZN(n_0_400));
   AND2_X1 i_0_0_604 (.A1(n_0_86), .A2(n_0_68), .ZN(n_0_401));
   AND2_X1 i_0_0_605 (.A1(n_0_87), .A2(n_0_68), .ZN(n_0_402));
   AND2_X1 i_0_0_606 (.A1(n_0_88), .A2(n_0_68), .ZN(n_0_403));
   AND2_X1 i_0_0_607 (.A1(n_0_89), .A2(n_0_68), .ZN(n_0_404));
   AND2_X1 i_0_0_608 (.A1(n_0_90), .A2(n_0_68), .ZN(n_0_405));
   AND2_X1 i_0_0_609 (.A1(n_0_91), .A2(n_0_68), .ZN(n_0_406));
   AND2_X1 i_0_0_610 (.A1(n_0_92), .A2(n_0_68), .ZN(n_0_407));
   AND2_X1 i_0_0_611 (.A1(n_0_93), .A2(n_0_68), .ZN(n_0_408));
   AND2_X1 i_0_0_612 (.A1(n_0_94), .A2(n_0_68), .ZN(n_0_409));
   AND2_X1 i_0_0_613 (.A1(n_0_95), .A2(n_0_68), .ZN(n_0_410));
   AND2_X1 i_0_0_614 (.A1(n_0_96), .A2(n_0_68), .ZN(n_0_411));
   AND2_X1 i_0_0_615 (.A1(n_0_97), .A2(n_0_68), .ZN(n_0_412));
   AND2_X1 i_0_0_616 (.A1(n_0_98), .A2(n_0_68), .ZN(n_0_413));
   OAI21_X1 i_0_0_617 (.A(n_0_0_399), .B1(n_0_0_369), .B2(n_0_0_368), .ZN(n_0_68));
   OAI22_X1 i_0_0_618 (.A1(n_0_389), .A2(n_0_0_831), .B1(n_0_0_758), .B2(n_0_390), 
      .ZN(n_0_0_368));
   AOI221_X1 i_0_0_619 (.A(n_0_0_370), .B1(n_0_0_829), .B2(n_0_388), .C1(n_0_389), 
      .C2(n_0_0_831), .ZN(n_0_0_369));
   AOI21_X1 i_0_0_620 (.A(n_0_0_371), .B1(n_0_0_373), .B2(n_0_0_372), .ZN(
      n_0_0_370));
   OAI22_X1 i_0_0_621 (.A1(n_0_388), .A2(n_0_0_829), .B1(n_0_0_827), .B2(n_0_387), 
      .ZN(n_0_0_371));
   AOI22_X1 i_0_0_622 (.A1(n_0_387), .A2(n_0_0_827), .B1(n_0_0_825), .B2(n_0_386), 
      .ZN(n_0_0_372));
   OAI221_X1 i_0_0_623 (.A(n_0_0_374), .B1(n_0_0_823), .B2(n_0_385), .C1(n_0_386), 
      .C2(n_0_0_825), .ZN(n_0_0_373));
   NAND2_X1 i_0_0_624 (.A1(n_0_0_376), .A2(n_0_0_375), .ZN(n_0_0_374));
   AOI22_X1 i_0_0_625 (.A1(n_0_385), .A2(n_0_0_823), .B1(n_0_0_821), .B2(n_0_384), 
      .ZN(n_0_0_375));
   OAI221_X1 i_0_0_626 (.A(n_0_0_377), .B1(n_0_0_819), .B2(n_0_383), .C1(n_0_384), 
      .C2(n_0_0_821), .ZN(n_0_0_376));
   OAI21_X1 i_0_0_627 (.A(n_0_0_378), .B1(n_0_0_380), .B2(n_0_0_379), .ZN(
      n_0_0_377));
   AOI22_X1 i_0_0_628 (.A1(n_0_382), .A2(n_0_0_817), .B1(n_0_0_819), .B2(n_0_383), 
      .ZN(n_0_0_378));
   OAI22_X1 i_0_0_629 (.A1(n_0_382), .A2(n_0_0_817), .B1(n_0_0_815), .B2(n_0_381), 
      .ZN(n_0_0_379));
   AOI221_X1 i_0_0_630 (.A(n_0_0_381), .B1(n_0_0_813), .B2(n_0_380), .C1(n_0_381), 
      .C2(n_0_0_815), .ZN(n_0_0_380));
   AOI21_X1 i_0_0_631 (.A(n_0_0_382), .B1(n_0_0_384), .B2(n_0_0_383), .ZN(
      n_0_0_381));
   OAI22_X1 i_0_0_632 (.A1(n_0_380), .A2(n_0_0_813), .B1(n_0_0_811), .B2(n_0_379), 
      .ZN(n_0_0_382));
   AOI22_X1 i_0_0_633 (.A1(n_0_379), .A2(n_0_0_811), .B1(n_0_0_809), .B2(n_0_378), 
      .ZN(n_0_0_383));
   OAI221_X1 i_0_0_634 (.A(n_0_0_385), .B1(n_0_0_807), .B2(n_0_377), .C1(n_0_378), 
      .C2(n_0_0_809), .ZN(n_0_0_384));
   OAI21_X1 i_0_0_635 (.A(n_0_0_386), .B1(n_0_0_388), .B2(n_0_0_387), .ZN(
      n_0_0_385));
   AOI22_X1 i_0_0_636 (.A1(n_0_377), .A2(n_0_0_807), .B1(n_0_0_805), .B2(n_0_376), 
      .ZN(n_0_0_386));
   OAI22_X1 i_0_0_637 (.A1(n_0_376), .A2(n_0_0_805), .B1(n_0_0_803), .B2(n_0_375), 
      .ZN(n_0_0_387));
   AOI221_X1 i_0_0_638 (.A(n_0_0_389), .B1(n_0_0_801), .B2(n_0_374), .C1(n_0_375), 
      .C2(n_0_0_803), .ZN(n_0_0_388));
   AOI21_X1 i_0_0_639 (.A(n_0_0_390), .B1(n_0_0_392), .B2(n_0_0_391), .ZN(
      n_0_0_389));
   OAI22_X1 i_0_0_640 (.A1(n_0_374), .A2(n_0_0_801), .B1(n_0_0_799), .B2(n_0_373), 
      .ZN(n_0_0_390));
   AOI22_X1 i_0_0_641 (.A1(n_0_373), .A2(n_0_0_799), .B1(n_0_0_797), .B2(n_0_372), 
      .ZN(n_0_0_391));
   OAI21_X1 i_0_0_642 (.A(n_0_0_393), .B1(n_0_0_797), .B2(n_0_372), .ZN(
      n_0_0_392));
   OAI21_X1 i_0_0_643 (.A(n_0_0_398), .B1(n_0_0_395), .B2(n_0_0_394), .ZN(
      n_0_0_393));
   OAI22_X1 i_0_0_644 (.A1(n_0_371), .A2(n_0_0_795), .B1(n_0_0_793), .B2(n_0_370), 
      .ZN(n_0_0_394));
   AOI221_X1 i_0_0_645 (.A(n_0_0_396), .B1(n_0_0_791), .B2(n_0_369), .C1(n_0_370), 
      .C2(n_0_0_793), .ZN(n_0_0_395));
   AOI21_X1 i_0_0_646 (.A(n_0_0_397), .B1(n_0_0_763), .B2(in_b[0]), .ZN(
      n_0_0_396));
   NOR2_X1 i_0_0_647 (.A1(n_0_369), .A2(n_0_0_791), .ZN(n_0_0_397));
   NAND2_X1 i_0_0_648 (.A1(n_0_371), .A2(n_0_0_795), .ZN(n_0_0_398));
   NAND2_X1 i_0_0_649 (.A1(n_0_390), .A2(n_0_0_758), .ZN(n_0_0_399));
   AND2_X1 i_0_0_650 (.A1(n_0_0_400), .A2(in_b[0]), .ZN(n_0_347));
   AND2_X1 i_0_0_651 (.A1(n_0_0_400), .A2(n_0_78), .ZN(n_0_348));
   AND2_X1 i_0_0_652 (.A1(n_0_0_400), .A2(n_0_79), .ZN(n_0_349));
   AND2_X1 i_0_0_653 (.A1(n_0_0_400), .A2(n_0_80), .ZN(n_0_350));
   AND2_X1 i_0_0_654 (.A1(n_0_0_400), .A2(n_0_81), .ZN(n_0_351));
   AND2_X1 i_0_0_655 (.A1(n_0_0_400), .A2(n_0_82), .ZN(n_0_352));
   AND2_X1 i_0_0_656 (.A1(n_0_0_400), .A2(n_0_83), .ZN(n_0_353));
   AND2_X1 i_0_0_657 (.A1(n_0_0_400), .A2(n_0_84), .ZN(n_0_354));
   AND2_X1 i_0_0_658 (.A1(n_0_0_400), .A2(n_0_85), .ZN(n_0_355));
   AND2_X1 i_0_0_659 (.A1(n_0_0_400), .A2(n_0_86), .ZN(n_0_356));
   AND2_X1 i_0_0_660 (.A1(n_0_0_400), .A2(n_0_87), .ZN(n_0_357));
   AND2_X1 i_0_0_661 (.A1(n_0_0_400), .A2(n_0_88), .ZN(n_0_358));
   AND2_X1 i_0_0_662 (.A1(n_0_0_400), .A2(n_0_89), .ZN(n_0_359));
   AND2_X1 i_0_0_663 (.A1(n_0_0_400), .A2(n_0_90), .ZN(n_0_360));
   AND2_X1 i_0_0_664 (.A1(n_0_0_400), .A2(n_0_91), .ZN(n_0_361));
   AND2_X1 i_0_0_665 (.A1(n_0_0_400), .A2(n_0_92), .ZN(n_0_362));
   AND2_X1 i_0_0_666 (.A1(n_0_0_400), .A2(n_0_93), .ZN(n_0_363));
   AND2_X1 i_0_0_667 (.A1(n_0_0_400), .A2(n_0_94), .ZN(n_0_364));
   AND2_X1 i_0_0_668 (.A1(n_0_0_400), .A2(n_0_95), .ZN(n_0_365));
   AND2_X1 i_0_0_669 (.A1(n_0_0_400), .A2(n_0_96), .ZN(n_0_366));
   AND2_X1 i_0_0_670 (.A1(n_0_0_400), .A2(n_0_97), .ZN(n_0_367));
   AND2_X1 i_0_0_671 (.A1(n_0_0_400), .A2(n_0_98), .ZN(n_0_368));
   OAI21_X1 i_0_0_672 (.A(n_0_0_431), .B1(n_0_0_402), .B2(n_0_0_401), .ZN(
      n_0_0_400));
   OAI22_X1 i_0_0_673 (.A1(n_0_344), .A2(n_0_0_831), .B1(n_0_0_758), .B2(n_0_345), 
      .ZN(n_0_0_401));
   AOI221_X1 i_0_0_674 (.A(n_0_0_403), .B1(n_0_0_829), .B2(n_0_343), .C1(n_0_344), 
      .C2(n_0_0_831), .ZN(n_0_0_402));
   AOI21_X1 i_0_0_675 (.A(n_0_0_404), .B1(n_0_0_406), .B2(n_0_0_405), .ZN(
      n_0_0_403));
   OAI22_X1 i_0_0_676 (.A1(n_0_343), .A2(n_0_0_829), .B1(n_0_0_827), .B2(n_0_342), 
      .ZN(n_0_0_404));
   AOI22_X1 i_0_0_677 (.A1(n_0_342), .A2(n_0_0_827), .B1(n_0_0_825), .B2(n_0_341), 
      .ZN(n_0_0_405));
   OAI221_X1 i_0_0_678 (.A(n_0_0_407), .B1(n_0_0_823), .B2(n_0_340), .C1(n_0_341), 
      .C2(n_0_0_825), .ZN(n_0_0_406));
   OAI21_X1 i_0_0_679 (.A(n_0_0_408), .B1(n_0_0_410), .B2(n_0_0_409), .ZN(
      n_0_0_407));
   AOI22_X1 i_0_0_680 (.A1(n_0_340), .A2(n_0_0_823), .B1(n_0_0_821), .B2(n_0_339), 
      .ZN(n_0_0_408));
   OAI22_X1 i_0_0_681 (.A1(n_0_339), .A2(n_0_0_821), .B1(n_0_0_819), .B2(n_0_338), 
      .ZN(n_0_0_409));
   AOI221_X1 i_0_0_682 (.A(n_0_0_411), .B1(n_0_0_817), .B2(n_0_337), .C1(n_0_338), 
      .C2(n_0_0_819), .ZN(n_0_0_410));
   INV_X1 i_0_0_683 (.A(n_0_0_412), .ZN(n_0_0_411));
   OAI221_X1 i_0_0_684 (.A(n_0_0_413), .B1(n_0_0_815), .B2(n_0_336), .C1(n_0_337), 
      .C2(n_0_0_817), .ZN(n_0_0_412));
   OAI21_X1 i_0_0_685 (.A(n_0_0_414), .B1(n_0_0_416), .B2(n_0_0_415), .ZN(
      n_0_0_413));
   AOI22_X1 i_0_0_686 (.A1(n_0_336), .A2(n_0_0_815), .B1(n_0_0_813), .B2(n_0_335), 
      .ZN(n_0_0_414));
   OAI22_X1 i_0_0_687 (.A1(n_0_335), .A2(n_0_0_813), .B1(n_0_0_811), .B2(n_0_334), 
      .ZN(n_0_0_415));
   AOI221_X1 i_0_0_688 (.A(n_0_0_417), .B1(n_0_0_809), .B2(n_0_333), .C1(n_0_334), 
      .C2(n_0_0_811), .ZN(n_0_0_416));
   AOI21_X1 i_0_0_689 (.A(n_0_0_418), .B1(n_0_0_420), .B2(n_0_0_419), .ZN(
      n_0_0_417));
   OAI22_X1 i_0_0_690 (.A1(n_0_333), .A2(n_0_0_809), .B1(n_0_0_807), .B2(n_0_332), 
      .ZN(n_0_0_418));
   AOI22_X1 i_0_0_691 (.A1(n_0_332), .A2(n_0_0_807), .B1(n_0_0_805), .B2(n_0_331), 
      .ZN(n_0_0_419));
   OAI221_X1 i_0_0_692 (.A(n_0_0_421), .B1(n_0_0_803), .B2(n_0_330), .C1(n_0_331), 
      .C2(n_0_0_805), .ZN(n_0_0_420));
   OAI21_X1 i_0_0_693 (.A(n_0_0_422), .B1(n_0_0_424), .B2(n_0_0_423), .ZN(
      n_0_0_421));
   AOI22_X1 i_0_0_694 (.A1(n_0_330), .A2(n_0_0_803), .B1(n_0_0_801), .B2(n_0_329), 
      .ZN(n_0_0_422));
   OAI22_X1 i_0_0_695 (.A1(n_0_329), .A2(n_0_0_801), .B1(n_0_0_799), .B2(n_0_328), 
      .ZN(n_0_0_423));
   AOI221_X1 i_0_0_696 (.A(n_0_0_425), .B1(n_0_0_797), .B2(n_0_327), .C1(n_0_328), 
      .C2(n_0_0_799), .ZN(n_0_0_424));
   AOI21_X1 i_0_0_697 (.A(n_0_0_426), .B1(n_0_526), .B2(n_0_0_858), .ZN(
      n_0_0_425));
   AOI21_X1 i_0_0_698 (.A(n_0_0_427), .B1(n_0_0_795), .B2(n_0_326), .ZN(
      n_0_0_426));
   AOI21_X1 i_0_0_699 (.A(n_0_0_428), .B1(n_0_0_430), .B2(n_0_0_429), .ZN(
      n_0_0_427));
   OAI22_X1 i_0_0_700 (.A1(n_0_326), .A2(n_0_0_795), .B1(n_0_0_793), .B2(n_0_325), 
      .ZN(n_0_0_428));
   AOI22_X1 i_0_0_701 (.A1(n_0_325), .A2(n_0_0_793), .B1(n_0_0_791), .B2(n_0_324), 
      .ZN(n_0_0_429));
   OAI22_X1 i_0_0_702 (.A1(n_0_77), .A2(n_0_0_861), .B1(n_0_324), .B2(n_0_0_791), 
      .ZN(n_0_0_430));
   NAND2_X1 i_0_0_703 (.A1(n_0_345), .A2(n_0_0_758), .ZN(n_0_0_431));
   AND2_X1 i_0_0_704 (.A1(n_0_0_432), .A2(in_b[0]), .ZN(n_0_302));
   AND2_X1 i_0_0_705 (.A1(n_0_0_432), .A2(n_0_78), .ZN(n_0_303));
   AND2_X1 i_0_0_706 (.A1(n_0_0_432), .A2(n_0_79), .ZN(n_0_304));
   AND2_X1 i_0_0_707 (.A1(n_0_0_432), .A2(n_0_80), .ZN(n_0_305));
   AND2_X1 i_0_0_708 (.A1(n_0_0_432), .A2(n_0_81), .ZN(n_0_306));
   AND2_X1 i_0_0_709 (.A1(n_0_0_432), .A2(n_0_82), .ZN(n_0_307));
   AND2_X1 i_0_0_710 (.A1(n_0_0_432), .A2(n_0_83), .ZN(n_0_308));
   AND2_X1 i_0_0_711 (.A1(n_0_0_432), .A2(n_0_84), .ZN(n_0_309));
   AND2_X1 i_0_0_712 (.A1(n_0_0_432), .A2(n_0_85), .ZN(n_0_310));
   AND2_X1 i_0_0_713 (.A1(n_0_0_432), .A2(n_0_86), .ZN(n_0_311));
   AND2_X1 i_0_0_714 (.A1(n_0_0_432), .A2(n_0_87), .ZN(n_0_312));
   AND2_X1 i_0_0_715 (.A1(n_0_0_432), .A2(n_0_88), .ZN(n_0_313));
   AND2_X1 i_0_0_716 (.A1(n_0_0_432), .A2(n_0_89), .ZN(n_0_314));
   AND2_X1 i_0_0_717 (.A1(n_0_0_432), .A2(n_0_90), .ZN(n_0_315));
   AND2_X1 i_0_0_718 (.A1(n_0_0_432), .A2(n_0_91), .ZN(n_0_316));
   AND2_X1 i_0_0_719 (.A1(n_0_0_432), .A2(n_0_92), .ZN(n_0_317));
   AND2_X1 i_0_0_720 (.A1(n_0_0_432), .A2(n_0_93), .ZN(n_0_318));
   AND2_X1 i_0_0_721 (.A1(n_0_0_432), .A2(n_0_94), .ZN(n_0_319));
   AND2_X1 i_0_0_722 (.A1(n_0_0_432), .A2(n_0_95), .ZN(n_0_320));
   AND2_X1 i_0_0_723 (.A1(n_0_0_432), .A2(n_0_96), .ZN(n_0_321));
   AND2_X1 i_0_0_724 (.A1(n_0_0_432), .A2(n_0_97), .ZN(n_0_322));
   AND2_X1 i_0_0_725 (.A1(n_0_0_432), .A2(n_0_98), .ZN(n_0_323));
   OAI21_X1 i_0_0_726 (.A(n_0_0_463), .B1(n_0_0_434), .B2(n_0_0_433), .ZN(
      n_0_0_432));
   OAI22_X1 i_0_0_727 (.A1(n_0_299), .A2(n_0_0_831), .B1(n_0_0_758), .B2(n_0_300), 
      .ZN(n_0_0_433));
   AOI221_X1 i_0_0_728 (.A(n_0_0_435), .B1(n_0_0_829), .B2(n_0_298), .C1(n_0_299), 
      .C2(n_0_0_831), .ZN(n_0_0_434));
   AOI21_X1 i_0_0_729 (.A(n_0_0_436), .B1(n_0_0_438), .B2(n_0_0_437), .ZN(
      n_0_0_435));
   OAI22_X1 i_0_0_730 (.A1(n_0_298), .A2(n_0_0_829), .B1(n_0_0_827), .B2(n_0_297), 
      .ZN(n_0_0_436));
   AOI22_X1 i_0_0_731 (.A1(n_0_297), .A2(n_0_0_827), .B1(n_0_0_825), .B2(n_0_296), 
      .ZN(n_0_0_437));
   OAI221_X1 i_0_0_732 (.A(n_0_0_439), .B1(n_0_0_823), .B2(n_0_295), .C1(n_0_296), 
      .C2(n_0_0_825), .ZN(n_0_0_438));
   NAND2_X1 i_0_0_733 (.A1(n_0_0_441), .A2(n_0_0_440), .ZN(n_0_0_439));
   AOI22_X1 i_0_0_734 (.A1(n_0_295), .A2(n_0_0_823), .B1(n_0_0_821), .B2(n_0_294), 
      .ZN(n_0_0_440));
   OAI221_X1 i_0_0_735 (.A(n_0_0_442), .B1(n_0_0_819), .B2(n_0_293), .C1(n_0_294), 
      .C2(n_0_0_821), .ZN(n_0_0_441));
   OAI21_X1 i_0_0_736 (.A(n_0_0_443), .B1(n_0_0_445), .B2(n_0_0_444), .ZN(
      n_0_0_442));
   AOI22_X1 i_0_0_737 (.A1(n_0_292), .A2(n_0_0_817), .B1(n_0_0_819), .B2(n_0_293), 
      .ZN(n_0_0_443));
   OAI22_X1 i_0_0_738 (.A1(n_0_292), .A2(n_0_0_817), .B1(n_0_0_815), .B2(n_0_291), 
      .ZN(n_0_0_444));
   AOI221_X1 i_0_0_739 (.A(n_0_0_446), .B1(n_0_0_813), .B2(n_0_290), .C1(n_0_291), 
      .C2(n_0_0_815), .ZN(n_0_0_445));
   NOR2_X1 i_0_0_740 (.A1(n_0_0_448), .A2(n_0_0_447), .ZN(n_0_0_446));
   OAI22_X1 i_0_0_741 (.A1(n_0_290), .A2(n_0_0_813), .B1(n_0_0_811), .B2(n_0_289), 
      .ZN(n_0_0_447));
   AOI221_X1 i_0_0_742 (.A(n_0_0_449), .B1(n_0_0_809), .B2(n_0_288), .C1(n_0_289), 
      .C2(n_0_0_811), .ZN(n_0_0_448));
   AOI21_X1 i_0_0_743 (.A(n_0_0_450), .B1(n_0_0_452), .B2(n_0_0_451), .ZN(
      n_0_0_449));
   OAI22_X1 i_0_0_744 (.A1(n_0_288), .A2(n_0_0_809), .B1(n_0_0_807), .B2(n_0_287), 
      .ZN(n_0_0_450));
   AOI22_X1 i_0_0_745 (.A1(n_0_287), .A2(n_0_0_807), .B1(n_0_0_805), .B2(n_0_286), 
      .ZN(n_0_0_451));
   OAI221_X1 i_0_0_746 (.A(n_0_0_453), .B1(n_0_0_803), .B2(n_0_285), .C1(n_0_286), 
      .C2(n_0_0_805), .ZN(n_0_0_452));
   OAI21_X1 i_0_0_747 (.A(n_0_0_454), .B1(n_0_0_456), .B2(n_0_0_455), .ZN(
      n_0_0_453));
   AOI22_X1 i_0_0_748 (.A1(n_0_285), .A2(n_0_0_803), .B1(n_0_0_801), .B2(n_0_284), 
      .ZN(n_0_0_454));
   OAI22_X1 i_0_0_749 (.A1(n_0_284), .A2(n_0_0_801), .B1(n_0_0_799), .B2(n_0_283), 
      .ZN(n_0_0_455));
   AOI221_X1 i_0_0_750 (.A(n_0_0_457), .B1(n_0_0_797), .B2(n_0_282), .C1(n_0_283), 
      .C2(n_0_0_799), .ZN(n_0_0_456));
   AOI21_X1 i_0_0_751 (.A(n_0_0_458), .B1(n_0_526), .B2(n_0_0_859), .ZN(
      n_0_0_457));
   AOI21_X1 i_0_0_752 (.A(n_0_0_459), .B1(n_0_0_795), .B2(n_0_281), .ZN(
      n_0_0_458));
   AOI21_X1 i_0_0_753 (.A(n_0_0_460), .B1(n_0_0_462), .B2(n_0_0_461), .ZN(
      n_0_0_459));
   OAI22_X1 i_0_0_754 (.A1(n_0_281), .A2(n_0_0_795), .B1(n_0_0_793), .B2(n_0_280), 
      .ZN(n_0_0_460));
   AOI22_X1 i_0_0_755 (.A1(n_0_280), .A2(n_0_0_793), .B1(n_0_0_791), .B2(n_0_279), 
      .ZN(n_0_0_461));
   OAI22_X1 i_0_0_756 (.A1(n_0_0_861), .A2(n_0_121), .B1(n_0_0_791), .B2(n_0_279), 
      .ZN(n_0_0_462));
   NAND2_X1 i_0_0_757 (.A1(n_0_300), .A2(n_0_0_758), .ZN(n_0_0_463));
   AND2_X1 i_0_0_758 (.A1(n_0_0_464), .A2(in_b[0]), .ZN(n_0_257));
   AND2_X1 i_0_0_759 (.A1(n_0_0_464), .A2(n_0_78), .ZN(n_0_258));
   AND2_X1 i_0_0_760 (.A1(n_0_0_464), .A2(n_0_79), .ZN(n_0_259));
   AND2_X1 i_0_0_761 (.A1(n_0_0_464), .A2(n_0_80), .ZN(n_0_260));
   AND2_X1 i_0_0_762 (.A1(n_0_0_464), .A2(n_0_81), .ZN(n_0_261));
   AND2_X1 i_0_0_763 (.A1(n_0_0_464), .A2(n_0_82), .ZN(n_0_262));
   AND2_X1 i_0_0_764 (.A1(n_0_0_464), .A2(n_0_83), .ZN(n_0_263));
   AND2_X1 i_0_0_765 (.A1(n_0_0_464), .A2(n_0_84), .ZN(n_0_264));
   AND2_X1 i_0_0_766 (.A1(n_0_0_464), .A2(n_0_85), .ZN(n_0_265));
   AND2_X1 i_0_0_767 (.A1(n_0_0_464), .A2(n_0_86), .ZN(n_0_266));
   AND2_X1 i_0_0_768 (.A1(n_0_0_464), .A2(n_0_87), .ZN(n_0_267));
   AND2_X1 i_0_0_769 (.A1(n_0_0_464), .A2(n_0_88), .ZN(n_0_268));
   AND2_X1 i_0_0_770 (.A1(n_0_0_464), .A2(n_0_89), .ZN(n_0_269));
   AND2_X1 i_0_0_771 (.A1(n_0_0_464), .A2(n_0_90), .ZN(n_0_270));
   AND2_X1 i_0_0_772 (.A1(n_0_0_464), .A2(n_0_91), .ZN(n_0_271));
   AND2_X1 i_0_0_773 (.A1(n_0_0_464), .A2(n_0_92), .ZN(n_0_272));
   AND2_X1 i_0_0_774 (.A1(n_0_0_464), .A2(n_0_93), .ZN(n_0_273));
   AND2_X1 i_0_0_775 (.A1(n_0_0_464), .A2(n_0_94), .ZN(n_0_274));
   AND2_X1 i_0_0_776 (.A1(n_0_0_464), .A2(n_0_95), .ZN(n_0_275));
   AND2_X1 i_0_0_777 (.A1(n_0_0_464), .A2(n_0_96), .ZN(n_0_276));
   AND2_X1 i_0_0_778 (.A1(n_0_0_464), .A2(n_0_97), .ZN(n_0_277));
   AND2_X1 i_0_0_779 (.A1(n_0_0_464), .A2(n_0_98), .ZN(n_0_278));
   OAI21_X1 i_0_0_780 (.A(n_0_0_495), .B1(n_0_0_466), .B2(n_0_0_465), .ZN(
      n_0_0_464));
   OAI22_X1 i_0_0_781 (.A1(n_0_254), .A2(n_0_0_831), .B1(n_0_0_758), .B2(n_0_255), 
      .ZN(n_0_0_465));
   AOI221_X1 i_0_0_782 (.A(n_0_0_467), .B1(n_0_0_829), .B2(n_0_253), .C1(n_0_254), 
      .C2(n_0_0_831), .ZN(n_0_0_466));
   AOI21_X1 i_0_0_783 (.A(n_0_0_468), .B1(n_0_0_470), .B2(n_0_0_469), .ZN(
      n_0_0_467));
   OAI22_X1 i_0_0_784 (.A1(n_0_253), .A2(n_0_0_829), .B1(n_0_0_827), .B2(n_0_252), 
      .ZN(n_0_0_468));
   AOI22_X1 i_0_0_785 (.A1(n_0_252), .A2(n_0_0_827), .B1(n_0_0_825), .B2(n_0_251), 
      .ZN(n_0_0_469));
   OAI221_X1 i_0_0_786 (.A(n_0_0_471), .B1(n_0_0_823), .B2(n_0_250), .C1(n_0_251), 
      .C2(n_0_0_825), .ZN(n_0_0_470));
   OAI21_X1 i_0_0_787 (.A(n_0_0_472), .B1(n_0_0_474), .B2(n_0_0_473), .ZN(
      n_0_0_471));
   AOI22_X1 i_0_0_788 (.A1(n_0_250), .A2(n_0_0_823), .B1(n_0_0_821), .B2(n_0_249), 
      .ZN(n_0_0_472));
   OAI22_X1 i_0_0_789 (.A1(n_0_249), .A2(n_0_0_821), .B1(n_0_0_819), .B2(n_0_248), 
      .ZN(n_0_0_473));
   AOI221_X1 i_0_0_790 (.A(n_0_0_475), .B1(n_0_0_817), .B2(n_0_247), .C1(n_0_248), 
      .C2(n_0_0_819), .ZN(n_0_0_474));
   AOI21_X1 i_0_0_791 (.A(n_0_0_476), .B1(n_0_0_478), .B2(n_0_0_477), .ZN(
      n_0_0_475));
   OAI22_X1 i_0_0_792 (.A1(n_0_247), .A2(n_0_0_817), .B1(n_0_0_815), .B2(n_0_246), 
      .ZN(n_0_0_476));
   AOI22_X1 i_0_0_793 (.A1(n_0_246), .A2(n_0_0_815), .B1(n_0_0_813), .B2(n_0_245), 
      .ZN(n_0_0_477));
   OAI221_X1 i_0_0_794 (.A(n_0_0_479), .B1(n_0_0_811), .B2(n_0_244), .C1(n_0_245), 
      .C2(n_0_0_813), .ZN(n_0_0_478));
   OAI21_X1 i_0_0_795 (.A(n_0_0_480), .B1(n_0_0_482), .B2(n_0_0_481), .ZN(
      n_0_0_479));
   AOI22_X1 i_0_0_796 (.A1(n_0_244), .A2(n_0_0_811), .B1(n_0_0_809), .B2(n_0_243), 
      .ZN(n_0_0_480));
   OAI22_X1 i_0_0_797 (.A1(n_0_243), .A2(n_0_0_809), .B1(n_0_0_807), .B2(n_0_242), 
      .ZN(n_0_0_481));
   AOI221_X1 i_0_0_798 (.A(n_0_0_483), .B1(n_0_0_805), .B2(n_0_241), .C1(n_0_242), 
      .C2(n_0_0_807), .ZN(n_0_0_482));
   AOI21_X1 i_0_0_799 (.A(n_0_0_484), .B1(n_0_0_486), .B2(n_0_0_485), .ZN(
      n_0_0_483));
   OAI22_X1 i_0_0_800 (.A1(n_0_241), .A2(n_0_0_805), .B1(n_0_0_803), .B2(n_0_240), 
      .ZN(n_0_0_484));
   AOI22_X1 i_0_0_801 (.A1(n_0_240), .A2(n_0_0_803), .B1(n_0_0_801), .B2(n_0_239), 
      .ZN(n_0_0_485));
   OAI221_X1 i_0_0_802 (.A(n_0_0_487), .B1(n_0_0_799), .B2(n_0_238), .C1(n_0_239), 
      .C2(n_0_0_801), .ZN(n_0_0_486));
   OAI21_X1 i_0_0_803 (.A(n_0_0_488), .B1(n_0_0_489), .B2(n_0_0_490), .ZN(
      n_0_0_487));
   AOI22_X1 i_0_0_804 (.A1(n_0_238), .A2(n_0_0_799), .B1(n_0_0_797), .B2(n_0_237), 
      .ZN(n_0_0_488));
   NOR2_X1 i_0_0_805 (.A1(n_0_237), .A2(n_0_0_797), .ZN(n_0_0_489));
   AOI21_X1 i_0_0_806 (.A(n_0_0_491), .B1(n_0_0_795), .B2(n_0_236), .ZN(
      n_0_0_490));
   AOI21_X1 i_0_0_807 (.A(n_0_0_492), .B1(n_0_0_494), .B2(n_0_0_493), .ZN(
      n_0_0_491));
   OAI22_X1 i_0_0_808 (.A1(n_0_236), .A2(n_0_0_795), .B1(n_0_0_793), .B2(n_0_235), 
      .ZN(n_0_0_492));
   AOI22_X1 i_0_0_809 (.A1(n_0_235), .A2(n_0_0_793), .B1(n_0_0_791), .B2(n_0_234), 
      .ZN(n_0_0_493));
   OAI22_X1 i_0_0_810 (.A1(n_0_166), .A2(n_0_0_861), .B1(n_0_234), .B2(n_0_0_791), 
      .ZN(n_0_0_494));
   NAND2_X1 i_0_0_811 (.A1(n_0_255), .A2(n_0_0_758), .ZN(n_0_0_495));
   AND2_X1 i_0_0_812 (.A1(n_0_0_496), .A2(in_b[0]), .ZN(n_0_212));
   AND2_X1 i_0_0_813 (.A1(n_0_0_496), .A2(n_0_78), .ZN(n_0_213));
   AND2_X1 i_0_0_814 (.A1(n_0_0_496), .A2(n_0_79), .ZN(n_0_214));
   AND2_X1 i_0_0_815 (.A1(n_0_0_496), .A2(n_0_80), .ZN(n_0_215));
   AND2_X1 i_0_0_816 (.A1(n_0_0_496), .A2(n_0_81), .ZN(n_0_216));
   AND2_X1 i_0_0_817 (.A1(n_0_0_496), .A2(n_0_82), .ZN(n_0_217));
   AND2_X1 i_0_0_818 (.A1(n_0_0_496), .A2(n_0_83), .ZN(n_0_218));
   AND2_X1 i_0_0_819 (.A1(n_0_0_496), .A2(n_0_84), .ZN(n_0_219));
   AND2_X1 i_0_0_820 (.A1(n_0_0_496), .A2(n_0_85), .ZN(n_0_220));
   AND2_X1 i_0_0_821 (.A1(n_0_0_496), .A2(n_0_86), .ZN(n_0_221));
   AND2_X1 i_0_0_822 (.A1(n_0_0_496), .A2(n_0_87), .ZN(n_0_222));
   AND2_X1 i_0_0_823 (.A1(n_0_0_496), .A2(n_0_88), .ZN(n_0_223));
   AND2_X1 i_0_0_824 (.A1(n_0_0_496), .A2(n_0_89), .ZN(n_0_224));
   AND2_X1 i_0_0_825 (.A1(n_0_0_496), .A2(n_0_90), .ZN(n_0_225));
   AND2_X1 i_0_0_826 (.A1(n_0_0_496), .A2(n_0_91), .ZN(n_0_226));
   AND2_X1 i_0_0_827 (.A1(n_0_0_496), .A2(n_0_92), .ZN(n_0_227));
   AND2_X1 i_0_0_828 (.A1(n_0_0_496), .A2(n_0_93), .ZN(n_0_228));
   AND2_X1 i_0_0_829 (.A1(n_0_0_496), .A2(n_0_94), .ZN(n_0_229));
   AND2_X1 i_0_0_830 (.A1(n_0_0_496), .A2(n_0_95), .ZN(n_0_230));
   AND2_X1 i_0_0_831 (.A1(n_0_0_496), .A2(n_0_96), .ZN(n_0_231));
   AND2_X1 i_0_0_832 (.A1(n_0_0_496), .A2(n_0_97), .ZN(n_0_232));
   AND2_X1 i_0_0_833 (.A1(n_0_0_496), .A2(n_0_98), .ZN(n_0_233));
   NAND2_X1 i_0_0_834 (.A1(n_0_0_527), .A2(n_0_0_497), .ZN(n_0_0_496));
   OAI221_X1 i_0_0_835 (.A(n_0_0_498), .B1(n_0_0_831), .B2(n_0_209), .C1(n_0_210), 
      .C2(n_0_0_758), .ZN(n_0_0_497));
   NAND2_X1 i_0_0_836 (.A1(n_0_0_500), .A2(n_0_0_499), .ZN(n_0_0_498));
   AOI22_X1 i_0_0_837 (.A1(n_0_209), .A2(n_0_0_831), .B1(n_0_0_829), .B2(n_0_208), 
      .ZN(n_0_0_499));
   OAI221_X1 i_0_0_838 (.A(n_0_0_501), .B1(n_0_0_827), .B2(n_0_207), .C1(n_0_208), 
      .C2(n_0_0_829), .ZN(n_0_0_500));
   OAI21_X1 i_0_0_839 (.A(n_0_0_502), .B1(n_0_0_504), .B2(n_0_0_503), .ZN(
      n_0_0_501));
   AOI22_X1 i_0_0_840 (.A1(n_0_207), .A2(n_0_0_827), .B1(n_0_0_825), .B2(n_0_206), 
      .ZN(n_0_0_502));
   OAI22_X1 i_0_0_841 (.A1(n_0_206), .A2(n_0_0_825), .B1(n_0_0_823), .B2(n_0_205), 
      .ZN(n_0_0_503));
   AOI221_X1 i_0_0_842 (.A(n_0_0_505), .B1(n_0_0_821), .B2(n_0_204), .C1(n_0_205), 
      .C2(n_0_0_823), .ZN(n_0_0_504));
   AOI21_X1 i_0_0_843 (.A(n_0_0_506), .B1(n_0_0_508), .B2(n_0_0_507), .ZN(
      n_0_0_505));
   OAI22_X1 i_0_0_844 (.A1(n_0_204), .A2(n_0_0_821), .B1(n_0_0_819), .B2(n_0_203), 
      .ZN(n_0_0_506));
   AOI22_X1 i_0_0_845 (.A1(n_0_202), .A2(n_0_0_817), .B1(n_0_0_819), .B2(n_0_203), 
      .ZN(n_0_0_507));
   OAI221_X1 i_0_0_846 (.A(n_0_0_509), .B1(n_0_0_815), .B2(n_0_201), .C1(n_0_202), 
      .C2(n_0_0_817), .ZN(n_0_0_508));
   OAI21_X1 i_0_0_847 (.A(n_0_0_510), .B1(n_0_0_512), .B2(n_0_0_511), .ZN(
      n_0_0_509));
   AOI22_X1 i_0_0_848 (.A1(n_0_201), .A2(n_0_0_815), .B1(n_0_0_813), .B2(n_0_200), 
      .ZN(n_0_0_510));
   OAI22_X1 i_0_0_849 (.A1(n_0_200), .A2(n_0_0_813), .B1(n_0_0_811), .B2(n_0_199), 
      .ZN(n_0_0_511));
   AOI221_X1 i_0_0_850 (.A(n_0_0_513), .B1(n_0_0_809), .B2(n_0_198), .C1(n_0_199), 
      .C2(n_0_0_811), .ZN(n_0_0_512));
   AOI21_X1 i_0_0_851 (.A(n_0_0_514), .B1(n_0_0_516), .B2(n_0_0_515), .ZN(
      n_0_0_513));
   OAI22_X1 i_0_0_852 (.A1(n_0_198), .A2(n_0_0_809), .B1(n_0_0_807), .B2(n_0_197), 
      .ZN(n_0_0_514));
   AOI22_X1 i_0_0_853 (.A1(n_0_197), .A2(n_0_0_807), .B1(n_0_0_805), .B2(n_0_196), 
      .ZN(n_0_0_515));
   OAI221_X1 i_0_0_854 (.A(n_0_0_517), .B1(n_0_0_803), .B2(n_0_195), .C1(n_0_196), 
      .C2(n_0_0_805), .ZN(n_0_0_516));
   OAI21_X1 i_0_0_855 (.A(n_0_0_518), .B1(n_0_0_520), .B2(n_0_0_519), .ZN(
      n_0_0_517));
   AOI22_X1 i_0_0_856 (.A1(n_0_195), .A2(n_0_0_803), .B1(n_0_0_801), .B2(n_0_194), 
      .ZN(n_0_0_518));
   OAI22_X1 i_0_0_857 (.A1(n_0_194), .A2(n_0_0_801), .B1(n_0_0_799), .B2(n_0_193), 
      .ZN(n_0_0_519));
   AOI221_X1 i_0_0_858 (.A(n_0_0_521), .B1(n_0_0_797), .B2(n_0_192), .C1(n_0_193), 
      .C2(n_0_0_799), .ZN(n_0_0_520));
   AOI21_X1 i_0_0_859 (.A(n_0_0_522), .B1(n_0_526), .B2(n_0_0_860), .ZN(
      n_0_0_521));
   AOI21_X1 i_0_0_860 (.A(n_0_0_523), .B1(n_0_0_795), .B2(n_0_191), .ZN(
      n_0_0_522));
   AOI21_X1 i_0_0_861 (.A(n_0_0_524), .B1(n_0_0_526), .B2(n_0_0_525), .ZN(
      n_0_0_523));
   OAI22_X1 i_0_0_862 (.A1(n_0_191), .A2(n_0_0_795), .B1(n_0_0_793), .B2(n_0_190), 
      .ZN(n_0_0_524));
   AOI22_X1 i_0_0_863 (.A1(n_0_190), .A2(n_0_0_793), .B1(n_0_0_791), .B2(n_0_189), 
      .ZN(n_0_0_525));
   OAI22_X1 i_0_0_864 (.A1(n_0_211), .A2(n_0_0_861), .B1(n_0_189), .B2(n_0_0_791), 
      .ZN(n_0_0_526));
   NAND2_X1 i_0_0_865 (.A1(n_0_210), .A2(n_0_0_758), .ZN(n_0_0_527));
   AND2_X1 i_0_0_866 (.A1(n_0_0_528), .A2(in_b[0]), .ZN(n_0_167));
   AND2_X1 i_0_0_867 (.A1(n_0_0_528), .A2(n_0_78), .ZN(n_0_168));
   AND2_X1 i_0_0_868 (.A1(n_0_0_528), .A2(n_0_79), .ZN(n_0_169));
   AND2_X1 i_0_0_869 (.A1(n_0_0_528), .A2(n_0_80), .ZN(n_0_170));
   AND2_X1 i_0_0_870 (.A1(n_0_0_528), .A2(n_0_81), .ZN(n_0_171));
   AND2_X1 i_0_0_871 (.A1(n_0_0_528), .A2(n_0_82), .ZN(n_0_172));
   AND2_X1 i_0_0_872 (.A1(n_0_0_528), .A2(n_0_83), .ZN(n_0_173));
   AND2_X1 i_0_0_873 (.A1(n_0_0_528), .A2(n_0_84), .ZN(n_0_174));
   AND2_X1 i_0_0_874 (.A1(n_0_0_528), .A2(n_0_85), .ZN(n_0_175));
   AND2_X1 i_0_0_875 (.A1(n_0_0_528), .A2(n_0_86), .ZN(n_0_176));
   AND2_X1 i_0_0_876 (.A1(n_0_0_528), .A2(n_0_87), .ZN(n_0_177));
   AND2_X1 i_0_0_877 (.A1(n_0_0_528), .A2(n_0_88), .ZN(n_0_178));
   AND2_X1 i_0_0_878 (.A1(n_0_0_528), .A2(n_0_89), .ZN(n_0_179));
   AND2_X1 i_0_0_879 (.A1(n_0_0_528), .A2(n_0_90), .ZN(n_0_180));
   AND2_X1 i_0_0_880 (.A1(n_0_0_528), .A2(n_0_91), .ZN(n_0_181));
   AND2_X1 i_0_0_881 (.A1(n_0_0_528), .A2(n_0_92), .ZN(n_0_182));
   AND2_X1 i_0_0_882 (.A1(n_0_0_528), .A2(n_0_93), .ZN(n_0_183));
   AND2_X1 i_0_0_883 (.A1(n_0_0_528), .A2(n_0_94), .ZN(n_0_184));
   AND2_X1 i_0_0_884 (.A1(n_0_0_528), .A2(n_0_95), .ZN(n_0_185));
   AND2_X1 i_0_0_885 (.A1(n_0_0_528), .A2(n_0_96), .ZN(n_0_186));
   AND2_X1 i_0_0_886 (.A1(n_0_0_528), .A2(n_0_97), .ZN(n_0_187));
   AND2_X1 i_0_0_887 (.A1(n_0_0_528), .A2(n_0_98), .ZN(n_0_188));
   OAI21_X1 i_0_0_888 (.A(n_0_0_560), .B1(n_0_0_530), .B2(n_0_0_529), .ZN(
      n_0_0_528));
   OAI22_X1 i_0_0_889 (.A1(n_0_164), .A2(n_0_0_831), .B1(n_0_0_758), .B2(n_0_165), 
      .ZN(n_0_0_529));
   AOI221_X1 i_0_0_890 (.A(n_0_0_531), .B1(n_0_0_829), .B2(n_0_163), .C1(n_0_164), 
      .C2(n_0_0_831), .ZN(n_0_0_530));
   AOI21_X1 i_0_0_891 (.A(n_0_0_532), .B1(n_0_0_534), .B2(n_0_0_533), .ZN(
      n_0_0_531));
   OAI22_X1 i_0_0_892 (.A1(n_0_163), .A2(n_0_0_829), .B1(n_0_0_827), .B2(n_0_162), 
      .ZN(n_0_0_532));
   AOI22_X1 i_0_0_893 (.A1(n_0_162), .A2(n_0_0_827), .B1(n_0_0_825), .B2(n_0_161), 
      .ZN(n_0_0_533));
   OAI221_X1 i_0_0_894 (.A(n_0_0_535), .B1(n_0_0_823), .B2(n_0_160), .C1(n_0_161), 
      .C2(n_0_0_825), .ZN(n_0_0_534));
   OAI21_X1 i_0_0_895 (.A(n_0_0_536), .B1(n_0_0_538), .B2(n_0_0_537), .ZN(
      n_0_0_535));
   AOI22_X1 i_0_0_896 (.A1(n_0_160), .A2(n_0_0_823), .B1(n_0_0_821), .B2(n_0_159), 
      .ZN(n_0_0_536));
   OAI22_X1 i_0_0_897 (.A1(n_0_159), .A2(n_0_0_821), .B1(n_0_0_819), .B2(n_0_158), 
      .ZN(n_0_0_537));
   AOI221_X1 i_0_0_898 (.A(n_0_0_539), .B1(n_0_0_817), .B2(n_0_157), .C1(n_0_158), 
      .C2(n_0_0_819), .ZN(n_0_0_538));
   AOI21_X1 i_0_0_899 (.A(n_0_0_540), .B1(n_0_0_542), .B2(n_0_0_541), .ZN(
      n_0_0_539));
   OAI22_X1 i_0_0_900 (.A1(n_0_157), .A2(n_0_0_817), .B1(n_0_0_815), .B2(n_0_156), 
      .ZN(n_0_0_540));
   AOI22_X1 i_0_0_901 (.A1(n_0_156), .A2(n_0_0_815), .B1(n_0_0_813), .B2(n_0_155), 
      .ZN(n_0_0_541));
   OAI221_X1 i_0_0_902 (.A(n_0_0_543), .B1(n_0_0_811), .B2(n_0_154), .C1(n_0_155), 
      .C2(n_0_0_813), .ZN(n_0_0_542));
   NAND2_X1 i_0_0_903 (.A1(n_0_0_545), .A2(n_0_0_544), .ZN(n_0_0_543));
   AOI22_X1 i_0_0_904 (.A1(n_0_154), .A2(n_0_0_811), .B1(n_0_0_809), .B2(n_0_153), 
      .ZN(n_0_0_544));
   OAI221_X1 i_0_0_905 (.A(n_0_0_546), .B1(n_0_0_807), .B2(n_0_152), .C1(n_0_153), 
      .C2(n_0_0_809), .ZN(n_0_0_545));
   OAI21_X1 i_0_0_906 (.A(n_0_0_547), .B1(n_0_0_549), .B2(n_0_0_548), .ZN(
      n_0_0_546));
   AOI22_X1 i_0_0_907 (.A1(n_0_152), .A2(n_0_0_807), .B1(n_0_0_805), .B2(n_0_151), 
      .ZN(n_0_0_547));
   OAI22_X1 i_0_0_908 (.A1(n_0_151), .A2(n_0_0_805), .B1(n_0_0_803), .B2(n_0_150), 
      .ZN(n_0_0_548));
   AOI221_X1 i_0_0_909 (.A(n_0_0_550), .B1(n_0_0_801), .B2(n_0_149), .C1(n_0_150), 
      .C2(n_0_0_803), .ZN(n_0_0_549));
   AOI21_X1 i_0_0_910 (.A(n_0_0_551), .B1(n_0_0_553), .B2(n_0_0_552), .ZN(
      n_0_0_550));
   OAI22_X1 i_0_0_911 (.A1(n_0_149), .A2(n_0_0_801), .B1(n_0_0_799), .B2(n_0_148), 
      .ZN(n_0_0_551));
   AOI22_X1 i_0_0_912 (.A1(n_0_148), .A2(n_0_0_799), .B1(n_0_0_797), .B2(n_0_147), 
      .ZN(n_0_0_552));
   OAI21_X1 i_0_0_913 (.A(n_0_0_554), .B1(n_0_0_797), .B2(n_0_147), .ZN(
      n_0_0_553));
   OAI21_X1 i_0_0_914 (.A(n_0_0_559), .B1(n_0_0_556), .B2(n_0_0_555), .ZN(
      n_0_0_554));
   OAI22_X1 i_0_0_915 (.A1(n_0_146), .A2(n_0_0_795), .B1(n_0_0_793), .B2(n_0_145), 
      .ZN(n_0_0_555));
   AOI221_X1 i_0_0_916 (.A(n_0_0_557), .B1(n_0_0_791), .B2(n_0_144), .C1(n_0_145), 
      .C2(n_0_0_793), .ZN(n_0_0_556));
   AOI21_X1 i_0_0_917 (.A(n_0_0_558), .B1(n_0_0_764), .B2(in_b[0]), .ZN(
      n_0_0_557));
   NOR2_X1 i_0_0_918 (.A1(n_0_144), .A2(n_0_0_791), .ZN(n_0_0_558));
   NAND2_X1 i_0_0_919 (.A1(n_0_146), .A2(n_0_0_795), .ZN(n_0_0_559));
   NAND2_X1 i_0_0_920 (.A1(n_0_165), .A2(n_0_0_758), .ZN(n_0_0_560));
   AND2_X1 i_0_0_921 (.A1(n_0_0_561), .A2(in_b[0]), .ZN(n_0_122));
   AND2_X1 i_0_0_922 (.A1(n_0_0_561), .A2(n_0_78), .ZN(n_0_123));
   AND2_X1 i_0_0_923 (.A1(n_0_0_561), .A2(n_0_79), .ZN(n_0_124));
   AND2_X1 i_0_0_924 (.A1(n_0_0_561), .A2(n_0_80), .ZN(n_0_125));
   AND2_X1 i_0_0_925 (.A1(n_0_0_561), .A2(n_0_81), .ZN(n_0_126));
   AND2_X1 i_0_0_926 (.A1(n_0_0_561), .A2(n_0_82), .ZN(n_0_127));
   AND2_X1 i_0_0_927 (.A1(n_0_0_561), .A2(n_0_83), .ZN(n_0_128));
   AND2_X1 i_0_0_928 (.A1(n_0_0_561), .A2(n_0_84), .ZN(n_0_129));
   AND2_X1 i_0_0_929 (.A1(n_0_0_561), .A2(n_0_85), .ZN(n_0_130));
   AND2_X1 i_0_0_930 (.A1(n_0_0_561), .A2(n_0_86), .ZN(n_0_131));
   AND2_X1 i_0_0_931 (.A1(n_0_0_561), .A2(n_0_87), .ZN(n_0_132));
   AND2_X1 i_0_0_932 (.A1(n_0_0_561), .A2(n_0_88), .ZN(n_0_133));
   AND2_X1 i_0_0_933 (.A1(n_0_0_561), .A2(n_0_89), .ZN(n_0_134));
   AND2_X1 i_0_0_934 (.A1(n_0_0_561), .A2(n_0_90), .ZN(n_0_135));
   AND2_X1 i_0_0_935 (.A1(n_0_0_561), .A2(n_0_91), .ZN(n_0_136));
   AND2_X1 i_0_0_936 (.A1(n_0_0_561), .A2(n_0_92), .ZN(n_0_137));
   AND2_X1 i_0_0_937 (.A1(n_0_0_561), .A2(n_0_93), .ZN(n_0_138));
   AND2_X1 i_0_0_938 (.A1(n_0_0_561), .A2(n_0_94), .ZN(n_0_139));
   AND2_X1 i_0_0_939 (.A1(n_0_0_561), .A2(n_0_95), .ZN(n_0_140));
   AND2_X1 i_0_0_940 (.A1(n_0_0_561), .A2(n_0_96), .ZN(n_0_141));
   AND2_X1 i_0_0_941 (.A1(n_0_0_561), .A2(n_0_97), .ZN(n_0_142));
   AND2_X1 i_0_0_942 (.A1(n_0_0_561), .A2(n_0_98), .ZN(n_0_143));
   NAND2_X1 i_0_0_943 (.A1(n_0_0_594), .A2(n_0_0_562), .ZN(n_0_0_561));
   OAI221_X1 i_0_0_944 (.A(n_0_0_563), .B1(n_0_0_831), .B2(divider[20]), 
      .C1(divider[21]), .C2(n_0_0_758), .ZN(n_0_0_562));
   NAND2_X1 i_0_0_945 (.A1(n_0_0_565), .A2(n_0_0_564), .ZN(n_0_0_563));
   AOI22_X1 i_0_0_946 (.A1(divider[20]), .A2(n_0_0_831), .B1(n_0_0_829), 
      .B2(divider[19]), .ZN(n_0_0_564));
   OAI221_X1 i_0_0_947 (.A(n_0_0_566), .B1(n_0_0_827), .B2(divider[18]), 
      .C1(divider[19]), .C2(n_0_0_829), .ZN(n_0_0_565));
   OAI21_X1 i_0_0_948 (.A(n_0_0_567), .B1(n_0_0_569), .B2(n_0_0_568), .ZN(
      n_0_0_566));
   AOI22_X1 i_0_0_949 (.A1(divider[18]), .A2(n_0_0_827), .B1(n_0_0_825), 
      .B2(divider[17]), .ZN(n_0_0_567));
   OAI22_X1 i_0_0_950 (.A1(divider[17]), .A2(n_0_0_825), .B1(n_0_0_823), 
      .B2(divider[16]), .ZN(n_0_0_568));
   AOI221_X1 i_0_0_951 (.A(n_0_0_570), .B1(n_0_0_821), .B2(divider[15]), 
      .C1(divider[16]), .C2(n_0_0_823), .ZN(n_0_0_569));
   AOI21_X1 i_0_0_952 (.A(n_0_0_571), .B1(n_0_0_573), .B2(n_0_0_572), .ZN(
      n_0_0_570));
   OAI22_X1 i_0_0_953 (.A1(divider[15]), .A2(n_0_0_821), .B1(n_0_0_819), 
      .B2(divider[14]), .ZN(n_0_0_571));
   AOI22_X1 i_0_0_954 (.A1(divider[13]), .A2(n_0_0_817), .B1(n_0_0_819), 
      .B2(divider[14]), .ZN(n_0_0_572));
   OAI221_X1 i_0_0_955 (.A(n_0_0_574), .B1(n_0_0_815), .B2(divider[12]), 
      .C1(divider[13]), .C2(n_0_0_817), .ZN(n_0_0_573));
   NAND2_X1 i_0_0_956 (.A1(n_0_0_576), .A2(n_0_0_575), .ZN(n_0_0_574));
   AOI22_X1 i_0_0_957 (.A1(divider[12]), .A2(n_0_0_815), .B1(n_0_0_813), 
      .B2(divider[11]), .ZN(n_0_0_575));
   OAI221_X1 i_0_0_958 (.A(n_0_0_577), .B1(n_0_0_811), .B2(divider[10]), 
      .C1(divider[11]), .C2(n_0_0_813), .ZN(n_0_0_576));
   NAND2_X1 i_0_0_959 (.A1(n_0_0_579), .A2(n_0_0_578), .ZN(n_0_0_577));
   AOI22_X1 i_0_0_960 (.A1(divider[10]), .A2(n_0_0_811), .B1(n_0_0_809), 
      .B2(divider[9]), .ZN(n_0_0_578));
   OAI221_X1 i_0_0_961 (.A(n_0_0_580), .B1(n_0_0_807), .B2(divider[8]), .C1(
      divider[9]), .C2(n_0_0_809), .ZN(n_0_0_579));
   OAI21_X1 i_0_0_962 (.A(n_0_0_581), .B1(n_0_0_583), .B2(n_0_0_582), .ZN(
      n_0_0_580));
   AOI22_X1 i_0_0_963 (.A1(divider[8]), .A2(n_0_0_807), .B1(n_0_0_805), .B2(
      divider[7]), .ZN(n_0_0_581));
   OAI22_X1 i_0_0_964 (.A1(divider[7]), .A2(n_0_0_805), .B1(n_0_0_803), .B2(
      divider[6]), .ZN(n_0_0_582));
   AOI221_X1 i_0_0_965 (.A(n_0_0_584), .B1(n_0_0_801), .B2(divider[5]), .C1(
      divider[6]), .C2(n_0_0_803), .ZN(n_0_0_583));
   AOI21_X1 i_0_0_966 (.A(n_0_0_585), .B1(n_0_0_587), .B2(n_0_0_586), .ZN(
      n_0_0_584));
   OAI22_X1 i_0_0_967 (.A1(divider[5]), .A2(n_0_0_801), .B1(n_0_0_799), .B2(
      divider[4]), .ZN(n_0_0_585));
   AOI22_X1 i_0_0_968 (.A1(divider[4]), .A2(n_0_0_799), .B1(n_0_0_797), .B2(
      divider[3]), .ZN(n_0_0_586));
   OAI21_X1 i_0_0_969 (.A(n_0_0_588), .B1(n_0_0_797), .B2(divider[3]), .ZN(
      n_0_0_587));
   OAI21_X1 i_0_0_970 (.A(n_0_0_593), .B1(n_0_0_590), .B2(n_0_0_589), .ZN(
      n_0_0_588));
   OAI22_X1 i_0_0_971 (.A1(divider[2]), .A2(n_0_0_795), .B1(n_0_0_793), .B2(
      divider[1]), .ZN(n_0_0_589));
   AOI221_X1 i_0_0_972 (.A(n_0_0_591), .B1(n_0_0_791), .B2(divider[0]), .C1(
      divider[1]), .C2(n_0_0_793), .ZN(n_0_0_590));
   AOI21_X1 i_0_0_973 (.A(n_0_0_592), .B1(n_0_0_765), .B2(in_b[0]), .ZN(
      n_0_0_591));
   NOR2_X1 i_0_0_974 (.A1(divider[0]), .A2(n_0_0_791), .ZN(n_0_0_592));
   NAND2_X1 i_0_0_975 (.A1(divider[2]), .A2(n_0_0_795), .ZN(n_0_0_593));
   NAND2_X1 i_0_0_976 (.A1(divider[21]), .A2(n_0_0_758), .ZN(n_0_0_594));
   NOR3_X1 i_0_0_977 (.A1(n_0_0_861), .A2(n_0_0_766), .A3(n_0_0_596), .ZN(n_0_99));
   AND2_X1 i_0_0_978 (.A1(n_0_78), .A2(n_0_0_595), .ZN(n_0_100));
   AND2_X1 i_0_0_979 (.A1(n_0_79), .A2(n_0_0_595), .ZN(n_0_101));
   AND2_X1 i_0_0_980 (.A1(n_0_80), .A2(n_0_0_595), .ZN(n_0_102));
   AND2_X1 i_0_0_981 (.A1(n_0_81), .A2(n_0_0_595), .ZN(n_0_103));
   AND2_X1 i_0_0_982 (.A1(n_0_82), .A2(n_0_0_595), .ZN(n_0_104));
   AND2_X1 i_0_0_983 (.A1(n_0_83), .A2(n_0_0_595), .ZN(n_0_105));
   AND2_X1 i_0_0_984 (.A1(n_0_84), .A2(n_0_0_595), .ZN(n_0_106));
   AND2_X1 i_0_0_985 (.A1(n_0_85), .A2(n_0_0_595), .ZN(n_0_107));
   AND2_X1 i_0_0_986 (.A1(n_0_86), .A2(n_0_0_595), .ZN(n_0_108));
   AND2_X1 i_0_0_987 (.A1(n_0_87), .A2(n_0_0_595), .ZN(n_0_109));
   AND2_X1 i_0_0_988 (.A1(n_0_88), .A2(n_0_0_595), .ZN(n_0_110));
   AND2_X1 i_0_0_989 (.A1(n_0_89), .A2(n_0_0_595), .ZN(n_0_111));
   AND2_X1 i_0_0_990 (.A1(n_0_90), .A2(n_0_0_595), .ZN(n_0_112));
   AND2_X1 i_0_0_991 (.A1(n_0_91), .A2(n_0_0_595), .ZN(n_0_113));
   AND2_X1 i_0_0_992 (.A1(n_0_92), .A2(n_0_0_595), .ZN(n_0_114));
   AND2_X1 i_0_0_993 (.A1(n_0_93), .A2(n_0_0_595), .ZN(n_0_115));
   AND2_X1 i_0_0_994 (.A1(n_0_94), .A2(n_0_0_595), .ZN(n_0_116));
   AND2_X1 i_0_0_995 (.A1(n_0_95), .A2(n_0_0_595), .ZN(n_0_117));
   AND2_X1 i_0_0_996 (.A1(n_0_96), .A2(n_0_0_595), .ZN(n_0_118));
   AND2_X1 i_0_0_997 (.A1(n_0_97), .A2(n_0_0_595), .ZN(n_0_119));
   AND2_X1 i_0_0_998 (.A1(n_0_98), .A2(n_0_0_595), .ZN(n_0_120));
   AOI21_X1 i_0_0_999 (.A(n_0_0_596), .B1(n_0_0_766), .B2(in_b[0]), .ZN(
      n_0_0_595));
   INV_X1 i_0_0_1000 (.A(n_0_0_597), .ZN(n_0_0_596));
   NOR3_X1 i_0_0_1001 (.A1(n_0_0_603), .A2(n_0_0_602), .A3(n_0_0_598), .ZN(
      n_0_0_597));
   NAND4_X1 i_0_0_1002 (.A1(n_0_0_825), .A2(n_0_0_823), .A3(n_0_0_604), .A4(
      n_0_0_599), .ZN(n_0_0_598));
   NOR3_X1 i_0_0_1003 (.A1(n_0_661), .A2(n_0_0_601), .A3(n_0_0_600), .ZN(
      n_0_0_599));
   NAND3_X1 i_0_0_1004 (.A1(n_0_0_801), .A2(n_0_0_799), .A3(n_0_0_797), .ZN(
      n_0_0_600));
   NAND4_X1 i_0_0_1005 (.A1(n_0_0_795), .A2(n_0_0_793), .A3(n_0_0_791), .A4(
      n_0_0_758), .ZN(n_0_0_601));
   NAND4_X1 i_0_0_1006 (.A1(n_0_0_817), .A2(n_0_0_815), .A3(n_0_0_813), .A4(
      n_0_0_819), .ZN(n_0_0_602));
   NAND4_X1 i_0_0_1007 (.A1(n_0_0_811), .A2(n_0_0_809), .A3(n_0_0_807), .A4(
      n_0_0_805), .ZN(n_0_0_603));
   NOR4_X1 i_0_0_1008 (.A1(n_0_1064), .A2(n_0_1063), .A3(n_0_1062), .A4(n_0_1017), 
      .ZN(n_0_0_604));
   OR2_X1 i_0_0_1009 (.A1(ovfl_flag), .A2(divide_by_zero_error), .ZN(err));
   AND2_X1 i_0_0_1010 (.A1(in_b[0]), .A2(n_0_1068), .ZN(n_0_973));
   AND2_X1 i_0_0_1011 (.A1(n_0_78), .A2(n_0_1068), .ZN(n_0_974));
   AND2_X1 i_0_0_1012 (.A1(n_0_79), .A2(n_0_1068), .ZN(n_0_975));
   AND2_X1 i_0_0_1013 (.A1(n_0_80), .A2(n_0_1068), .ZN(n_0_976));
   AND2_X1 i_0_0_1014 (.A1(n_0_81), .A2(n_0_1068), .ZN(n_0_977));
   AND2_X1 i_0_0_1015 (.A1(n_0_82), .A2(n_0_1068), .ZN(n_0_978));
   AND2_X1 i_0_0_1016 (.A1(n_0_83), .A2(n_0_1068), .ZN(n_0_979));
   AND2_X1 i_0_0_1017 (.A1(n_0_84), .A2(n_0_1068), .ZN(n_0_980));
   AND2_X1 i_0_0_1018 (.A1(n_0_85), .A2(n_0_1068), .ZN(n_0_981));
   AND2_X1 i_0_0_1019 (.A1(n_0_86), .A2(n_0_1068), .ZN(n_0_982));
   AND2_X1 i_0_0_1020 (.A1(n_0_87), .A2(n_0_1068), .ZN(n_0_983));
   AND2_X1 i_0_0_1021 (.A1(n_0_88), .A2(n_0_1068), .ZN(n_0_984));
   AND2_X1 i_0_0_1022 (.A1(n_0_89), .A2(n_0_1068), .ZN(n_0_985));
   AND2_X1 i_0_0_1023 (.A1(n_0_90), .A2(n_0_1068), .ZN(n_0_986));
   AND2_X1 i_0_0_1024 (.A1(n_0_91), .A2(n_0_1068), .ZN(n_0_987));
   AND2_X1 i_0_0_1025 (.A1(n_0_92), .A2(n_0_1068), .ZN(n_0_988));
   AND2_X1 i_0_0_1026 (.A1(n_0_93), .A2(n_0_1068), .ZN(n_0_989));
   AND2_X1 i_0_0_1027 (.A1(n_0_94), .A2(n_0_1068), .ZN(n_0_990));
   AND2_X1 i_0_0_1028 (.A1(n_0_95), .A2(n_0_1068), .ZN(n_0_991));
   AND2_X1 i_0_0_1029 (.A1(n_0_96), .A2(n_0_1068), .ZN(n_0_992));
   AND2_X1 i_0_0_1030 (.A1(n_0_97), .A2(n_0_1068), .ZN(n_0_993));
   AND2_X1 i_0_0_1031 (.A1(n_0_98), .A2(n_0_1068), .ZN(n_0_994));
   AOI21_X1 i_0_0_1032 (.A(n_0_0_636), .B1(n_0_0_606), .B2(n_0_0_605), .ZN(
      n_0_1068));
   AOI22_X1 i_0_0_1033 (.A1(n_0_970), .A2(n_0_0_831), .B1(n_0_0_758), .B2(
      n_0_971), .ZN(n_0_0_605));
   OAI221_X1 i_0_0_1034 (.A(n_0_0_607), .B1(n_0_0_829), .B2(n_0_969), .C1(
      n_0_970), .C2(n_0_0_831), .ZN(n_0_0_606));
   NAND2_X1 i_0_0_1035 (.A1(n_0_0_609), .A2(n_0_0_608), .ZN(n_0_0_607));
   AOI22_X1 i_0_0_1036 (.A1(n_0_969), .A2(n_0_0_829), .B1(n_0_0_827), .B2(
      n_0_968), .ZN(n_0_0_608));
   OAI221_X1 i_0_0_1037 (.A(n_0_0_610), .B1(n_0_0_825), .B2(n_0_967), .C1(
      n_0_968), .C2(n_0_0_827), .ZN(n_0_0_609));
   OAI21_X1 i_0_0_1038 (.A(n_0_0_611), .B1(n_0_0_613), .B2(n_0_0_612), .ZN(
      n_0_0_610));
   AOI22_X1 i_0_0_1039 (.A1(n_0_967), .A2(n_0_0_825), .B1(n_0_0_823), .B2(
      n_0_966), .ZN(n_0_0_611));
   OAI22_X1 i_0_0_1040 (.A1(n_0_966), .A2(n_0_0_823), .B1(n_0_0_821), .B2(
      n_0_965), .ZN(n_0_0_612));
   AOI221_X1 i_0_0_1041 (.A(n_0_0_614), .B1(n_0_0_819), .B2(n_0_964), .C1(
      n_0_965), .C2(n_0_0_821), .ZN(n_0_0_613));
   INV_X1 i_0_0_1042 (.A(n_0_0_615), .ZN(n_0_0_614));
   OAI21_X1 i_0_0_1043 (.A(n_0_0_616), .B1(n_0_0_819), .B2(n_0_964), .ZN(
      n_0_0_615));
   OAI21_X1 i_0_0_1044 (.A(n_0_0_635), .B1(n_0_0_618), .B2(n_0_0_617), .ZN(
      n_0_0_616));
   OAI22_X1 i_0_0_1045 (.A1(n_0_963), .A2(n_0_0_817), .B1(n_0_0_815), .B2(
      n_0_962), .ZN(n_0_0_617));
   AOI221_X1 i_0_0_1046 (.A(n_0_0_619), .B1(n_0_0_813), .B2(n_0_961), .C1(
      n_0_962), .C2(n_0_0_815), .ZN(n_0_0_618));
   AOI21_X1 i_0_0_1047 (.A(n_0_0_620), .B1(n_0_0_622), .B2(n_0_0_621), .ZN(
      n_0_0_619));
   OAI22_X1 i_0_0_1048 (.A1(n_0_961), .A2(n_0_0_813), .B1(n_0_0_811), .B2(
      n_0_960), .ZN(n_0_0_620));
   AOI22_X1 i_0_0_1049 (.A1(n_0_960), .A2(n_0_0_811), .B1(n_0_0_809), .B2(
      n_0_959), .ZN(n_0_0_621));
   OAI221_X1 i_0_0_1050 (.A(n_0_0_623), .B1(n_0_0_807), .B2(n_0_958), .C1(
      n_0_959), .C2(n_0_0_809), .ZN(n_0_0_622));
   OAI21_X1 i_0_0_1051 (.A(n_0_0_624), .B1(n_0_0_626), .B2(n_0_0_625), .ZN(
      n_0_0_623));
   AOI22_X1 i_0_0_1052 (.A1(n_0_958), .A2(n_0_0_807), .B1(n_0_0_805), .B2(
      n_0_957), .ZN(n_0_0_624));
   OAI22_X1 i_0_0_1053 (.A1(n_0_957), .A2(n_0_0_805), .B1(n_0_0_803), .B2(
      n_0_956), .ZN(n_0_0_625));
   AOI221_X1 i_0_0_1054 (.A(n_0_0_627), .B1(n_0_0_801), .B2(n_0_955), .C1(
      n_0_956), .C2(n_0_0_803), .ZN(n_0_0_626));
   AOI21_X1 i_0_0_1055 (.A(n_0_0_628), .B1(n_0_0_630), .B2(n_0_0_629), .ZN(
      n_0_0_627));
   OAI22_X1 i_0_0_1056 (.A1(n_0_955), .A2(n_0_0_801), .B1(n_0_0_799), .B2(
      n_0_954), .ZN(n_0_0_628));
   AOI22_X1 i_0_0_1057 (.A1(n_0_954), .A2(n_0_0_799), .B1(n_0_0_797), .B2(
      n_0_953), .ZN(n_0_0_629));
   OAI21_X1 i_0_0_1058 (.A(n_0_0_631), .B1(n_0_0_797), .B2(n_0_953), .ZN(
      n_0_0_630));
   OAI21_X1 i_0_0_1059 (.A(n_0_0_634), .B1(n_0_0_633), .B2(n_0_0_632), .ZN(
      n_0_0_631));
   OAI22_X1 i_0_0_1060 (.A1(n_0_952), .A2(n_0_0_795), .B1(n_0_0_793), .B2(
      n_0_951), .ZN(n_0_0_632));
   AOI221_X1 i_0_0_1061 (.A(n_0_0_754), .B1(n_0_0_793), .B2(n_0_951), .C1(
      n_0_1069), .C2(n_0_0_791), .ZN(n_0_0_633));
   NAND2_X1 i_0_0_1062 (.A1(n_0_952), .A2(n_0_0_795), .ZN(n_0_0_634));
   NAND2_X1 i_0_0_1063 (.A1(n_0_963), .A2(n_0_0_817), .ZN(n_0_0_635));
   NOR2_X1 i_0_0_1064 (.A1(n_0_971), .A2(n_0_0_758), .ZN(n_0_0_636));
   AND2_X1 i_0_0_1065 (.A1(n_0_1069), .A2(in_b[0]), .ZN(n_0_929));
   AND2_X1 i_0_0_1066 (.A1(n_0_1069), .A2(n_0_78), .ZN(n_0_930));
   AND2_X1 i_0_0_1067 (.A1(n_0_1069), .A2(n_0_79), .ZN(n_0_931));
   AND2_X1 i_0_0_1068 (.A1(n_0_1069), .A2(n_0_80), .ZN(n_0_932));
   AND2_X1 i_0_0_1069 (.A1(n_0_1069), .A2(n_0_81), .ZN(n_0_933));
   AND2_X1 i_0_0_1070 (.A1(n_0_1069), .A2(n_0_82), .ZN(n_0_934));
   AND2_X1 i_0_0_1071 (.A1(n_0_1069), .A2(n_0_83), .ZN(n_0_935));
   AND2_X1 i_0_0_1072 (.A1(n_0_1069), .A2(n_0_84), .ZN(n_0_936));
   AND2_X1 i_0_0_1073 (.A1(n_0_1069), .A2(n_0_85), .ZN(n_0_937));
   AND2_X1 i_0_0_1074 (.A1(n_0_1069), .A2(n_0_86), .ZN(n_0_938));
   AND2_X1 i_0_0_1075 (.A1(n_0_1069), .A2(n_0_87), .ZN(n_0_939));
   AND2_X1 i_0_0_1076 (.A1(n_0_1069), .A2(n_0_88), .ZN(n_0_940));
   AND2_X1 i_0_0_1077 (.A1(n_0_1069), .A2(n_0_89), .ZN(n_0_941));
   AND2_X1 i_0_0_1078 (.A1(n_0_1069), .A2(n_0_90), .ZN(n_0_942));
   AND2_X1 i_0_0_1079 (.A1(n_0_1069), .A2(n_0_91), .ZN(n_0_943));
   AND2_X1 i_0_0_1080 (.A1(n_0_1069), .A2(n_0_92), .ZN(n_0_944));
   AND2_X1 i_0_0_1081 (.A1(n_0_1069), .A2(n_0_93), .ZN(n_0_945));
   AND2_X1 i_0_0_1082 (.A1(n_0_1069), .A2(n_0_94), .ZN(n_0_946));
   AND2_X1 i_0_0_1083 (.A1(n_0_1069), .A2(n_0_95), .ZN(n_0_947));
   AND2_X1 i_0_0_1084 (.A1(n_0_1069), .A2(n_0_96), .ZN(n_0_948));
   AND2_X1 i_0_0_1085 (.A1(n_0_1069), .A2(n_0_97), .ZN(n_0_949));
   AND2_X1 i_0_0_1086 (.A1(n_0_1069), .A2(n_0_98), .ZN(n_0_950));
   OAI21_X1 i_0_0_1087 (.A(n_0_0_665), .B1(n_0_0_638), .B2(n_0_0_637), .ZN(
      n_0_1069));
   OAI22_X1 i_0_0_1088 (.A1(n_0_926), .A2(n_0_0_831), .B1(n_0_0_758), .B2(
      n_0_927), .ZN(n_0_0_637));
   AOI221_X1 i_0_0_1089 (.A(n_0_0_639), .B1(n_0_0_829), .B2(n_0_925), .C1(
      n_0_926), .C2(n_0_0_831), .ZN(n_0_0_638));
   AOI21_X1 i_0_0_1090 (.A(n_0_0_640), .B1(n_0_0_642), .B2(n_0_0_641), .ZN(
      n_0_0_639));
   OAI22_X1 i_0_0_1091 (.A1(n_0_925), .A2(n_0_0_829), .B1(n_0_0_827), .B2(
      n_0_924), .ZN(n_0_0_640));
   AOI22_X1 i_0_0_1092 (.A1(n_0_924), .A2(n_0_0_827), .B1(n_0_0_825), .B2(
      n_0_923), .ZN(n_0_0_641));
   OAI221_X1 i_0_0_1093 (.A(n_0_0_643), .B1(n_0_0_823), .B2(n_0_922), .C1(
      n_0_923), .C2(n_0_0_825), .ZN(n_0_0_642));
   OAI21_X1 i_0_0_1094 (.A(n_0_0_644), .B1(n_0_0_646), .B2(n_0_0_645), .ZN(
      n_0_0_643));
   AOI22_X1 i_0_0_1095 (.A1(n_0_922), .A2(n_0_0_823), .B1(n_0_0_821), .B2(
      n_0_921), .ZN(n_0_0_644));
   OAI22_X1 i_0_0_1096 (.A1(n_0_921), .A2(n_0_0_821), .B1(n_0_0_819), .B2(
      n_0_920), .ZN(n_0_0_645));
   AOI221_X1 i_0_0_1097 (.A(n_0_0_647), .B1(n_0_0_817), .B2(n_0_919), .C1(
      n_0_920), .C2(n_0_0_819), .ZN(n_0_0_646));
   AOI21_X1 i_0_0_1098 (.A(n_0_0_648), .B1(n_0_0_650), .B2(n_0_0_649), .ZN(
      n_0_0_647));
   OAI22_X1 i_0_0_1099 (.A1(n_0_919), .A2(n_0_0_817), .B1(n_0_0_815), .B2(
      n_0_918), .ZN(n_0_0_648));
   AOI22_X1 i_0_0_1100 (.A1(n_0_918), .A2(n_0_0_815), .B1(n_0_0_813), .B2(
      n_0_917), .ZN(n_0_0_649));
   OAI221_X1 i_0_0_1101 (.A(n_0_0_651), .B1(n_0_0_811), .B2(n_0_916), .C1(
      n_0_917), .C2(n_0_0_813), .ZN(n_0_0_650));
   OAI21_X1 i_0_0_1102 (.A(n_0_0_652), .B1(n_0_0_654), .B2(n_0_0_653), .ZN(
      n_0_0_651));
   AOI22_X1 i_0_0_1103 (.A1(n_0_916), .A2(n_0_0_811), .B1(n_0_0_809), .B2(
      n_0_915), .ZN(n_0_0_652));
   OAI22_X1 i_0_0_1104 (.A1(n_0_915), .A2(n_0_0_809), .B1(n_0_0_807), .B2(
      n_0_914), .ZN(n_0_0_653));
   AOI221_X1 i_0_0_1105 (.A(n_0_0_655), .B1(n_0_0_805), .B2(n_0_913), .C1(
      n_0_914), .C2(n_0_0_807), .ZN(n_0_0_654));
   AOI21_X1 i_0_0_1106 (.A(n_0_0_656), .B1(n_0_0_658), .B2(n_0_0_657), .ZN(
      n_0_0_655));
   OAI22_X1 i_0_0_1107 (.A1(n_0_913), .A2(n_0_0_805), .B1(n_0_0_803), .B2(
      n_0_912), .ZN(n_0_0_656));
   AOI22_X1 i_0_0_1108 (.A1(n_0_912), .A2(n_0_0_803), .B1(n_0_0_801), .B2(
      n_0_911), .ZN(n_0_0_657));
   OAI221_X1 i_0_0_1109 (.A(n_0_0_659), .B1(n_0_0_799), .B2(n_0_910), .C1(
      n_0_911), .C2(n_0_0_801), .ZN(n_0_0_658));
   OAI21_X1 i_0_0_1110 (.A(n_0_0_660), .B1(n_0_0_662), .B2(n_0_0_661), .ZN(
      n_0_0_659));
   AOI22_X1 i_0_0_1111 (.A1(n_0_910), .A2(n_0_0_799), .B1(n_0_0_797), .B2(
      n_0_909), .ZN(n_0_0_660));
   OAI22_X1 i_0_0_1112 (.A1(n_0_909), .A2(n_0_0_797), .B1(n_0_0_795), .B2(
      n_0_908), .ZN(n_0_0_661));
   AOI221_X1 i_0_0_1113 (.A(n_0_0_663), .B1(n_0_0_793), .B2(n_0_907), .C1(
      n_0_908), .C2(n_0_0_795), .ZN(n_0_0_662));
   AOI21_X1 i_0_0_1114 (.A(n_0_0_664), .B1(n_0_0_666), .B2(in_b[0]), .ZN(
      n_0_0_663));
   OAI21_X1 i_0_0_1115 (.A(n_0_0_791), .B1(n_0_0_793), .B2(n_0_907), .ZN(
      n_0_0_664));
   NAND2_X1 i_0_0_1116 (.A1(n_0_927), .A2(n_0_0_758), .ZN(n_0_0_665));
   NOR2_X1 i_0_0_1117 (.A1(n_0_0_666), .A2(n_0_0_861), .ZN(n_0_885));
   NOR2_X1 i_0_0_1118 (.A1(n_0_0_666), .A2(n_0_0_834), .ZN(n_0_886));
   NOR2_X1 i_0_0_1119 (.A1(n_0_0_666), .A2(n_0_0_835), .ZN(n_0_887));
   NOR2_X1 i_0_0_1120 (.A1(n_0_0_666), .A2(n_0_0_836), .ZN(n_0_888));
   NOR2_X1 i_0_0_1121 (.A1(n_0_0_666), .A2(n_0_0_837), .ZN(n_0_889));
   NOR2_X1 i_0_0_1122 (.A1(n_0_0_666), .A2(n_0_0_838), .ZN(n_0_890));
   NOR2_X1 i_0_0_1123 (.A1(n_0_0_666), .A2(n_0_0_839), .ZN(n_0_891));
   NOR2_X1 i_0_0_1124 (.A1(n_0_0_666), .A2(n_0_0_840), .ZN(n_0_892));
   NOR2_X1 i_0_0_1125 (.A1(n_0_0_666), .A2(n_0_0_841), .ZN(n_0_893));
   NOR2_X1 i_0_0_1126 (.A1(n_0_0_666), .A2(n_0_0_842), .ZN(n_0_894));
   NOR2_X1 i_0_0_1127 (.A1(n_0_0_666), .A2(n_0_0_843), .ZN(n_0_895));
   NOR2_X1 i_0_0_1128 (.A1(n_0_0_666), .A2(n_0_0_844), .ZN(n_0_896));
   NOR2_X1 i_0_0_1129 (.A1(n_0_0_666), .A2(n_0_0_845), .ZN(n_0_897));
   NOR2_X1 i_0_0_1130 (.A1(n_0_0_666), .A2(n_0_0_846), .ZN(n_0_898));
   NOR2_X1 i_0_0_1131 (.A1(n_0_0_666), .A2(n_0_0_847), .ZN(n_0_899));
   NOR2_X1 i_0_0_1132 (.A1(n_0_0_666), .A2(n_0_0_848), .ZN(n_0_900));
   NOR2_X1 i_0_0_1133 (.A1(n_0_0_666), .A2(n_0_0_849), .ZN(n_0_901));
   NOR2_X1 i_0_0_1134 (.A1(n_0_0_666), .A2(n_0_0_850), .ZN(n_0_902));
   NOR2_X1 i_0_0_1135 (.A1(n_0_0_666), .A2(n_0_0_851), .ZN(n_0_903));
   NOR2_X1 i_0_0_1136 (.A1(n_0_0_666), .A2(n_0_0_852), .ZN(n_0_904));
   NOR2_X1 i_0_0_1137 (.A1(n_0_0_666), .A2(n_0_0_853), .ZN(n_0_905));
   NOR2_X1 i_0_0_1138 (.A1(n_0_0_666), .A2(n_0_0_854), .ZN(n_0_906));
   INV_X1 i_0_0_1139 (.A(n_0_1070), .ZN(n_0_0_666));
   OAI21_X1 i_0_0_1140 (.A(n_0_0_667), .B1(n_0_0_669), .B2(n_0_0_668), .ZN(
      n_0_1070));
   NAND2_X1 i_0_0_1141 (.A1(n_0_883), .A2(n_0_0_758), .ZN(n_0_0_667));
   OAI22_X1 i_0_0_1142 (.A1(n_0_882), .A2(n_0_0_831), .B1(n_0_0_758), .B2(
      n_0_883), .ZN(n_0_0_668));
   AOI221_X1 i_0_0_1143 (.A(n_0_0_670), .B1(n_0_0_829), .B2(n_0_881), .C1(
      n_0_882), .C2(n_0_0_831), .ZN(n_0_0_669));
   AOI21_X1 i_0_0_1144 (.A(n_0_0_671), .B1(n_0_0_673), .B2(n_0_0_672), .ZN(
      n_0_0_670));
   OAI22_X1 i_0_0_1145 (.A1(n_0_881), .A2(n_0_0_829), .B1(n_0_0_827), .B2(
      n_0_880), .ZN(n_0_0_671));
   AOI22_X1 i_0_0_1146 (.A1(n_0_880), .A2(n_0_0_827), .B1(n_0_0_825), .B2(
      n_0_879), .ZN(n_0_0_672));
   OAI221_X1 i_0_0_1147 (.A(n_0_0_674), .B1(n_0_0_823), .B2(n_0_878), .C1(
      n_0_879), .C2(n_0_0_825), .ZN(n_0_0_673));
   OAI21_X1 i_0_0_1148 (.A(n_0_0_675), .B1(n_0_0_677), .B2(n_0_0_676), .ZN(
      n_0_0_674));
   AOI22_X1 i_0_0_1149 (.A1(n_0_878), .A2(n_0_0_823), .B1(n_0_0_821), .B2(
      n_0_877), .ZN(n_0_0_675));
   OAI22_X1 i_0_0_1150 (.A1(n_0_877), .A2(n_0_0_821), .B1(n_0_0_819), .B2(
      n_0_876), .ZN(n_0_0_676));
   AOI221_X1 i_0_0_1151 (.A(n_0_0_678), .B1(n_0_0_817), .B2(n_0_875), .C1(
      n_0_876), .C2(n_0_0_819), .ZN(n_0_0_677));
   AOI21_X1 i_0_0_1152 (.A(n_0_0_679), .B1(n_0_0_681), .B2(n_0_0_680), .ZN(
      n_0_0_678));
   OAI22_X1 i_0_0_1153 (.A1(n_0_875), .A2(n_0_0_817), .B1(n_0_0_815), .B2(
      n_0_874), .ZN(n_0_0_679));
   AOI22_X1 i_0_0_1154 (.A1(n_0_874), .A2(n_0_0_815), .B1(n_0_0_813), .B2(
      n_0_873), .ZN(n_0_0_680));
   OAI221_X1 i_0_0_1155 (.A(n_0_0_682), .B1(n_0_0_811), .B2(n_0_872), .C1(
      n_0_873), .C2(n_0_0_813), .ZN(n_0_0_681));
   OAI21_X1 i_0_0_1156 (.A(n_0_0_683), .B1(n_0_0_685), .B2(n_0_0_684), .ZN(
      n_0_0_682));
   AOI22_X1 i_0_0_1157 (.A1(n_0_872), .A2(n_0_0_811), .B1(n_0_0_809), .B2(
      n_0_871), .ZN(n_0_0_683));
   OAI22_X1 i_0_0_1158 (.A1(n_0_871), .A2(n_0_0_809), .B1(n_0_0_807), .B2(
      n_0_870), .ZN(n_0_0_684));
   AOI221_X1 i_0_0_1159 (.A(n_0_0_686), .B1(n_0_0_805), .B2(n_0_869), .C1(
      n_0_870), .C2(n_0_0_807), .ZN(n_0_0_685));
   AOI21_X1 i_0_0_1160 (.A(n_0_0_687), .B1(n_0_0_689), .B2(n_0_0_688), .ZN(
      n_0_0_686));
   OAI22_X1 i_0_0_1161 (.A1(n_0_869), .A2(n_0_0_805), .B1(n_0_0_803), .B2(
      n_0_868), .ZN(n_0_0_687));
   AOI22_X1 i_0_0_1162 (.A1(n_0_868), .A2(n_0_0_803), .B1(n_0_0_801), .B2(
      n_0_867), .ZN(n_0_0_688));
   OAI221_X1 i_0_0_1163 (.A(n_0_0_690), .B1(n_0_0_799), .B2(n_0_866), .C1(
      n_0_867), .C2(n_0_0_801), .ZN(n_0_0_689));
   OAI21_X1 i_0_0_1164 (.A(n_0_0_691), .B1(n_0_0_693), .B2(n_0_0_692), .ZN(
      n_0_0_690));
   AOI22_X1 i_0_0_1165 (.A1(n_0_866), .A2(n_0_0_799), .B1(n_0_0_797), .B2(
      n_0_865), .ZN(n_0_0_691));
   OAI22_X1 i_0_0_1166 (.A1(n_0_865), .A2(n_0_0_797), .B1(n_0_0_795), .B2(
      n_0_864), .ZN(n_0_0_692));
   AOI221_X1 i_0_0_1167 (.A(n_0_0_694), .B1(n_0_0_793), .B2(n_0_863), .C1(
      n_0_864), .C2(n_0_0_795), .ZN(n_0_0_693));
   AOI21_X1 i_0_0_1168 (.A(n_0_0_695), .B1(n_0_0_696), .B2(in_b[0]), .ZN(
      n_0_0_694));
   OAI21_X1 i_0_0_1169 (.A(n_0_0_791), .B1(n_0_0_793), .B2(n_0_863), .ZN(
      n_0_0_695));
   NOR2_X1 i_0_0_1170 (.A1(n_0_0_696), .A2(n_0_0_861), .ZN(n_0_841));
   NOR2_X1 i_0_0_1171 (.A1(n_0_0_696), .A2(n_0_0_834), .ZN(n_0_842));
   NOR2_X1 i_0_0_1172 (.A1(n_0_0_696), .A2(n_0_0_835), .ZN(n_0_843));
   NOR2_X1 i_0_0_1173 (.A1(n_0_0_696), .A2(n_0_0_836), .ZN(n_0_844));
   NOR2_X1 i_0_0_1174 (.A1(n_0_0_696), .A2(n_0_0_837), .ZN(n_0_845));
   NOR2_X1 i_0_0_1175 (.A1(n_0_0_696), .A2(n_0_0_838), .ZN(n_0_846));
   NOR2_X1 i_0_0_1176 (.A1(n_0_0_696), .A2(n_0_0_839), .ZN(n_0_847));
   NOR2_X1 i_0_0_1177 (.A1(n_0_0_696), .A2(n_0_0_840), .ZN(n_0_848));
   NOR2_X1 i_0_0_1178 (.A1(n_0_0_696), .A2(n_0_0_841), .ZN(n_0_849));
   NOR2_X1 i_0_0_1179 (.A1(n_0_0_696), .A2(n_0_0_842), .ZN(n_0_850));
   NOR2_X1 i_0_0_1180 (.A1(n_0_0_696), .A2(n_0_0_843), .ZN(n_0_851));
   NOR2_X1 i_0_0_1181 (.A1(n_0_0_696), .A2(n_0_0_844), .ZN(n_0_852));
   NOR2_X1 i_0_0_1182 (.A1(n_0_0_696), .A2(n_0_0_845), .ZN(n_0_853));
   NOR2_X1 i_0_0_1183 (.A1(n_0_0_696), .A2(n_0_0_846), .ZN(n_0_854));
   NOR2_X1 i_0_0_1184 (.A1(n_0_0_696), .A2(n_0_0_847), .ZN(n_0_855));
   NOR2_X1 i_0_0_1185 (.A1(n_0_0_696), .A2(n_0_0_848), .ZN(n_0_856));
   NOR2_X1 i_0_0_1186 (.A1(n_0_0_696), .A2(n_0_0_849), .ZN(n_0_857));
   NOR2_X1 i_0_0_1187 (.A1(n_0_0_696), .A2(n_0_0_850), .ZN(n_0_858));
   NOR2_X1 i_0_0_1188 (.A1(n_0_0_696), .A2(n_0_0_851), .ZN(n_0_859));
   NOR2_X1 i_0_0_1189 (.A1(n_0_0_696), .A2(n_0_0_852), .ZN(n_0_860));
   NOR2_X1 i_0_0_1190 (.A1(n_0_0_696), .A2(n_0_0_853), .ZN(n_0_861));
   NOR2_X1 i_0_0_1191 (.A1(n_0_0_696), .A2(n_0_0_854), .ZN(n_0_862));
   INV_X1 i_0_0_1192 (.A(n_0_1071), .ZN(n_0_0_696));
   NAND2_X1 i_0_0_1193 (.A1(n_0_0_725), .A2(n_0_0_697), .ZN(n_0_1071));
   OAI221_X1 i_0_0_1194 (.A(n_0_0_698), .B1(n_0_0_831), .B2(n_0_838), .C1(
      n_0_839), .C2(n_0_0_758), .ZN(n_0_0_697));
   NAND2_X1 i_0_0_1195 (.A1(n_0_0_700), .A2(n_0_0_699), .ZN(n_0_0_698));
   AOI22_X1 i_0_0_1196 (.A1(n_0_838), .A2(n_0_0_831), .B1(n_0_0_829), .B2(
      n_0_837), .ZN(n_0_0_699));
   OAI221_X1 i_0_0_1197 (.A(n_0_0_701), .B1(n_0_0_827), .B2(n_0_836), .C1(
      n_0_837), .C2(n_0_0_829), .ZN(n_0_0_700));
   OAI21_X1 i_0_0_1198 (.A(n_0_0_702), .B1(n_0_0_704), .B2(n_0_0_703), .ZN(
      n_0_0_701));
   AOI22_X1 i_0_0_1199 (.A1(n_0_836), .A2(n_0_0_827), .B1(n_0_0_825), .B2(
      n_0_835), .ZN(n_0_0_702));
   OAI22_X1 i_0_0_1200 (.A1(n_0_835), .A2(n_0_0_825), .B1(n_0_0_823), .B2(
      n_0_834), .ZN(n_0_0_703));
   AOI221_X1 i_0_0_1201 (.A(n_0_0_705), .B1(n_0_0_821), .B2(n_0_833), .C1(
      n_0_834), .C2(n_0_0_823), .ZN(n_0_0_704));
   AOI21_X1 i_0_0_1202 (.A(n_0_0_706), .B1(n_0_0_708), .B2(n_0_0_707), .ZN(
      n_0_0_705));
   OAI22_X1 i_0_0_1203 (.A1(n_0_833), .A2(n_0_0_821), .B1(n_0_0_819), .B2(
      n_0_832), .ZN(n_0_0_706));
   AOI22_X1 i_0_0_1204 (.A1(n_0_831), .A2(n_0_0_817), .B1(n_0_0_819), .B2(
      n_0_832), .ZN(n_0_0_707));
   OAI221_X1 i_0_0_1205 (.A(n_0_0_709), .B1(n_0_0_815), .B2(n_0_830), .C1(
      n_0_831), .C2(n_0_0_817), .ZN(n_0_0_708));
   OAI21_X1 i_0_0_1206 (.A(n_0_0_710), .B1(n_0_0_712), .B2(n_0_0_711), .ZN(
      n_0_0_709));
   AOI22_X1 i_0_0_1207 (.A1(n_0_830), .A2(n_0_0_815), .B1(n_0_0_813), .B2(
      n_0_829), .ZN(n_0_0_710));
   OAI22_X1 i_0_0_1208 (.A1(n_0_829), .A2(n_0_0_813), .B1(n_0_0_811), .B2(
      n_0_828), .ZN(n_0_0_711));
   AOI221_X1 i_0_0_1209 (.A(n_0_0_713), .B1(n_0_0_809), .B2(n_0_827), .C1(
      n_0_828), .C2(n_0_0_811), .ZN(n_0_0_712));
   AOI21_X1 i_0_0_1210 (.A(n_0_0_714), .B1(n_0_0_716), .B2(n_0_0_715), .ZN(
      n_0_0_713));
   OAI22_X1 i_0_0_1211 (.A1(n_0_827), .A2(n_0_0_809), .B1(n_0_0_807), .B2(
      n_0_826), .ZN(n_0_0_714));
   AOI22_X1 i_0_0_1212 (.A1(n_0_826), .A2(n_0_0_807), .B1(n_0_0_805), .B2(
      n_0_825), .ZN(n_0_0_715));
   OAI221_X1 i_0_0_1213 (.A(n_0_0_717), .B1(n_0_0_803), .B2(n_0_824), .C1(
      n_0_825), .C2(n_0_0_805), .ZN(n_0_0_716));
   OAI21_X1 i_0_0_1214 (.A(n_0_0_718), .B1(n_0_0_720), .B2(n_0_0_719), .ZN(
      n_0_0_717));
   AOI22_X1 i_0_0_1215 (.A1(n_0_824), .A2(n_0_0_803), .B1(n_0_0_801), .B2(
      n_0_823), .ZN(n_0_0_718));
   OAI22_X1 i_0_0_1216 (.A1(n_0_823), .A2(n_0_0_801), .B1(n_0_0_799), .B2(
      n_0_822), .ZN(n_0_0_719));
   AOI221_X1 i_0_0_1217 (.A(n_0_0_721), .B1(n_0_0_797), .B2(n_0_821), .C1(
      n_0_822), .C2(n_0_0_799), .ZN(n_0_0_720));
   AOI21_X1 i_0_0_1218 (.A(n_0_0_722), .B1(n_0_0_724), .B2(n_0_0_723), .ZN(
      n_0_0_721));
   OAI22_X1 i_0_0_1219 (.A1(n_0_821), .A2(n_0_0_797), .B1(n_0_0_795), .B2(
      n_0_820), .ZN(n_0_0_722));
   AOI22_X1 i_0_0_1220 (.A1(n_0_820), .A2(n_0_0_795), .B1(n_0_0_793), .B2(
      n_0_819), .ZN(n_0_0_723));
   OAI221_X1 i_0_0_1221 (.A(n_0_0_791), .B1(n_0_0_793), .B2(n_0_819), .C1(
      n_0_0_861), .C2(n_0_1072), .ZN(n_0_0_724));
   NAND2_X1 i_0_0_1222 (.A1(n_0_839), .A2(n_0_0_758), .ZN(n_0_0_725));
   AND2_X1 i_0_0_1223 (.A1(n_0_1072), .A2(in_b[0]), .ZN(n_0_797));
   AND2_X1 i_0_0_1224 (.A1(n_0_1072), .A2(n_0_78), .ZN(n_0_798));
   AND2_X1 i_0_0_1225 (.A1(n_0_1072), .A2(n_0_79), .ZN(n_0_799));
   AND2_X1 i_0_0_1226 (.A1(n_0_1072), .A2(n_0_80), .ZN(n_0_800));
   AND2_X1 i_0_0_1227 (.A1(n_0_1072), .A2(n_0_81), .ZN(n_0_801));
   AND2_X1 i_0_0_1228 (.A1(n_0_1072), .A2(n_0_82), .ZN(n_0_802));
   AND2_X1 i_0_0_1229 (.A1(n_0_1072), .A2(n_0_83), .ZN(n_0_803));
   AND2_X1 i_0_0_1230 (.A1(n_0_1072), .A2(n_0_84), .ZN(n_0_804));
   AND2_X1 i_0_0_1231 (.A1(n_0_1072), .A2(n_0_85), .ZN(n_0_805));
   AND2_X1 i_0_0_1232 (.A1(n_0_1072), .A2(n_0_86), .ZN(n_0_806));
   AND2_X1 i_0_0_1233 (.A1(n_0_1072), .A2(n_0_87), .ZN(n_0_807));
   AND2_X1 i_0_0_1234 (.A1(n_0_1072), .A2(n_0_88), .ZN(n_0_808));
   AND2_X1 i_0_0_1235 (.A1(n_0_1072), .A2(n_0_89), .ZN(n_0_809));
   AND2_X1 i_0_0_1236 (.A1(n_0_1072), .A2(n_0_90), .ZN(n_0_810));
   AND2_X1 i_0_0_1237 (.A1(n_0_1072), .A2(n_0_91), .ZN(n_0_811));
   AND2_X1 i_0_0_1238 (.A1(n_0_1072), .A2(n_0_92), .ZN(n_0_812));
   AND2_X1 i_0_0_1239 (.A1(n_0_1072), .A2(n_0_93), .ZN(n_0_813));
   AND2_X1 i_0_0_1240 (.A1(n_0_1072), .A2(n_0_94), .ZN(n_0_814));
   AND2_X1 i_0_0_1241 (.A1(n_0_1072), .A2(n_0_95), .ZN(n_0_815));
   AND2_X1 i_0_0_1242 (.A1(n_0_1072), .A2(n_0_96), .ZN(n_0_816));
   AND2_X1 i_0_0_1243 (.A1(n_0_1072), .A2(n_0_97), .ZN(n_0_817));
   AND2_X1 i_0_0_1244 (.A1(n_0_1072), .A2(n_0_98), .ZN(n_0_818));
   NAND2_X1 i_0_0_1245 (.A1(n_0_0_757), .A2(n_0_0_726), .ZN(n_0_1072));
   OAI221_X1 i_0_0_1246 (.A(n_0_0_727), .B1(n_0_0_831), .B2(n_0_794), .C1(
      n_0_795), .C2(n_0_0_758), .ZN(n_0_0_726));
   OAI21_X1 i_0_0_1247 (.A(n_0_0_728), .B1(n_0_0_730), .B2(n_0_0_729), .ZN(
      n_0_0_727));
   AOI22_X1 i_0_0_1248 (.A1(n_0_794), .A2(n_0_0_831), .B1(n_0_0_829), .B2(
      n_0_793), .ZN(n_0_0_728));
   OAI22_X1 i_0_0_1249 (.A1(n_0_793), .A2(n_0_0_829), .B1(n_0_0_827), .B2(
      n_0_792), .ZN(n_0_0_729));
   AOI221_X1 i_0_0_1250 (.A(n_0_0_731), .B1(n_0_0_825), .B2(n_0_791), .C1(
      n_0_792), .C2(n_0_0_827), .ZN(n_0_0_730));
   AOI21_X1 i_0_0_1251 (.A(n_0_0_732), .B1(n_0_0_734), .B2(n_0_0_733), .ZN(
      n_0_0_731));
   OAI22_X1 i_0_0_1252 (.A1(n_0_791), .A2(n_0_0_825), .B1(n_0_0_823), .B2(
      n_0_790), .ZN(n_0_0_732));
   AOI22_X1 i_0_0_1253 (.A1(n_0_790), .A2(n_0_0_823), .B1(n_0_0_821), .B2(
      n_0_789), .ZN(n_0_0_733));
   OAI221_X1 i_0_0_1254 (.A(n_0_0_735), .B1(n_0_0_819), .B2(n_0_788), .C1(
      n_0_789), .C2(n_0_0_821), .ZN(n_0_0_734));
   OAI21_X1 i_0_0_1255 (.A(n_0_0_736), .B1(n_0_0_738), .B2(n_0_0_737), .ZN(
      n_0_0_735));
   AOI22_X1 i_0_0_1256 (.A1(n_0_787), .A2(n_0_0_817), .B1(n_0_0_819), .B2(
      n_0_788), .ZN(n_0_0_736));
   OAI22_X1 i_0_0_1257 (.A1(n_0_787), .A2(n_0_0_817), .B1(n_0_0_815), .B2(
      n_0_786), .ZN(n_0_0_737));
   AOI221_X1 i_0_0_1258 (.A(n_0_0_739), .B1(n_0_0_813), .B2(n_0_785), .C1(
      n_0_786), .C2(n_0_0_815), .ZN(n_0_0_738));
   AOI21_X1 i_0_0_1259 (.A(n_0_0_740), .B1(n_0_0_742), .B2(n_0_0_741), .ZN(
      n_0_0_739));
   OAI22_X1 i_0_0_1260 (.A1(n_0_785), .A2(n_0_0_813), .B1(n_0_0_811), .B2(
      n_0_784), .ZN(n_0_0_740));
   AOI22_X1 i_0_0_1261 (.A1(n_0_784), .A2(n_0_0_811), .B1(n_0_0_809), .B2(
      n_0_783), .ZN(n_0_0_741));
   OAI221_X1 i_0_0_1262 (.A(n_0_0_743), .B1(n_0_0_807), .B2(n_0_782), .C1(
      n_0_783), .C2(n_0_0_809), .ZN(n_0_0_742));
   OAI21_X1 i_0_0_1263 (.A(n_0_0_744), .B1(n_0_0_746), .B2(n_0_0_745), .ZN(
      n_0_0_743));
   AOI22_X1 i_0_0_1264 (.A1(n_0_782), .A2(n_0_0_807), .B1(n_0_0_805), .B2(
      n_0_781), .ZN(n_0_0_744));
   OAI22_X1 i_0_0_1265 (.A1(n_0_781), .A2(n_0_0_805), .B1(n_0_0_803), .B2(
      n_0_780), .ZN(n_0_0_745));
   AOI221_X1 i_0_0_1266 (.A(n_0_0_747), .B1(n_0_0_801), .B2(n_0_779), .C1(
      n_0_780), .C2(n_0_0_803), .ZN(n_0_0_746));
   AOI21_X1 i_0_0_1267 (.A(n_0_0_748), .B1(n_0_0_750), .B2(n_0_0_749), .ZN(
      n_0_0_747));
   OAI22_X1 i_0_0_1268 (.A1(n_0_779), .A2(n_0_0_801), .B1(n_0_0_799), .B2(
      n_0_778), .ZN(n_0_0_748));
   AOI22_X1 i_0_0_1269 (.A1(n_0_778), .A2(n_0_0_799), .B1(n_0_0_797), .B2(
      n_0_777), .ZN(n_0_0_749));
   OAI21_X1 i_0_0_1270 (.A(n_0_0_751), .B1(n_0_0_797), .B2(n_0_777), .ZN(
      n_0_0_750));
   OAI21_X1 i_0_0_1271 (.A(n_0_0_756), .B1(n_0_0_753), .B2(n_0_0_752), .ZN(
      n_0_0_751));
   OAI22_X1 i_0_0_1272 (.A1(n_0_776), .A2(n_0_0_795), .B1(n_0_0_793), .B2(
      n_0_775), .ZN(n_0_0_752));
   AOI221_X1 i_0_0_1273 (.A(n_0_0_754), .B1(n_0_0_755), .B2(n_0_774), .C1(
      n_0_775), .C2(n_0_0_793), .ZN(n_0_0_753));
   NOR2_X1 i_0_0_1274 (.A1(n_0_391), .A2(in_b[0]), .ZN(n_0_0_754));
   NAND2_X1 i_0_0_1275 (.A1(n_0_391), .A2(in_b[0]), .ZN(n_0_0_755));
   NAND2_X1 i_0_0_1276 (.A1(n_0_776), .A2(n_0_0_795), .ZN(n_0_0_756));
   NAND2_X1 i_0_0_1277 (.A1(n_0_795), .A2(n_0_0_758), .ZN(n_0_0_757));
   OAI21_X1 i_0_0_1278 (.A(n_0_0_759), .B1(n_0_22), .B2(n_0_0_862), .ZN(
      n_0_0_758));
   OR2_X1 i_0_0_1279 (.A1(in_b[63]), .A2(in_b[22]), .ZN(n_0_0_759));
   XNOR2_X1 i_0_0_1280 (.A(in_a[1]), .B(n_0_0_789), .ZN(n_0_69));
   XNOR2_X1 i_0_0_1281 (.A(in_a[2]), .B(n_0_0_788), .ZN(n_0_70));
   XNOR2_X1 i_0_0_1282 (.A(in_a[3]), .B(n_0_0_786), .ZN(n_0_71));
   XOR2_X1 i_0_0_1283 (.A(in_a[4]), .B(n_0_0_784), .Z(n_0_72));
   INV_X1 i_0_0_1284 (.A(n_0_0_760), .ZN(n_0_73));
   XOR2_X1 i_0_0_1285 (.A(in_a[5]), .B(n_0_0_783), .Z(n_0_0_760));
   INV_X1 i_0_0_1286 (.A(n_0_0_761), .ZN(n_0_74));
   NAND2_X1 i_0_0_1287 (.A1(n_0_0_781), .A2(n_0_0_762), .ZN(n_0_0_761));
   NAND2_X1 i_0_0_1288 (.A1(n_0_0_782), .A2(in_a[6]), .ZN(n_0_0_762));
   XNOR2_X1 i_0_0_1289 (.A(in_a[7]), .B(n_0_0_780), .ZN(n_0_75));
   INV_X1 i_0_0_1290 (.A(n_0_0_763), .ZN(n_0_76));
   XOR2_X1 i_0_0_1291 (.A(in_a[8]), .B(n_0_0_779), .Z(n_0_0_763));
   XOR2_X1 i_0_0_1292 (.A(in_a[9]), .B(n_0_0_777), .Z(n_0_77));
   XNOR2_X1 i_0_0_1293 (.A(in_a[10]), .B(n_0_0_773), .ZN(n_0_121));
   XNOR2_X1 i_0_0_1294 (.A(in_a[11]), .B(n_0_0_772), .ZN(n_0_166));
   XNOR2_X1 i_0_0_1295 (.A(in_a[12]), .B(n_0_0_771), .ZN(n_0_211));
   INV_X1 i_0_0_1296 (.A(n_0_0_764), .ZN(n_0_256));
   XNOR2_X1 i_0_0_1297 (.A(in_a[13]), .B(n_0_0_770), .ZN(n_0_0_764));
   INV_X1 i_0_0_1298 (.A(n_0_0_765), .ZN(n_0_301));
   XNOR2_X1 i_0_0_1299 (.A(in_a[14]), .B(n_0_0_768), .ZN(n_0_0_765));
   INV_X1 i_0_0_1300 (.A(n_0_346), .ZN(n_0_0_766));
   XNOR2_X1 i_0_0_1301 (.A(in_a[15]), .B(n_0_0_767), .ZN(n_0_346));
   OAI21_X1 i_0_0_1302 (.A(in_a[63]), .B1(n_0_0_769), .B2(in_a[14]), .ZN(
      n_0_0_767));
   AND2_X1 i_0_0_1303 (.A1(n_0_0_769), .A2(in_a[63]), .ZN(n_0_0_768));
   OR2_X1 i_0_0_1304 (.A1(in_a[13]), .A2(n_0_0_770), .ZN(n_0_0_769));
   NAND2_X1 i_0_0_1305 (.A1(n_0_0_771), .A2(n_0_0_775), .ZN(n_0_0_770));
   AND2_X1 i_0_0_1306 (.A1(n_0_0_772), .A2(n_0_0_774), .ZN(n_0_0_771));
   OAI21_X1 i_0_0_1307 (.A(in_a[63]), .B1(n_0_0_776), .B2(in_a[10]), .ZN(
      n_0_0_772));
   NAND2_X1 i_0_0_1308 (.A1(n_0_0_776), .A2(in_a[63]), .ZN(n_0_0_773));
   NAND2_X1 i_0_0_1309 (.A1(in_a[63]), .A2(in_a[11]), .ZN(n_0_0_774));
   NAND2_X1 i_0_0_1310 (.A1(in_a[63]), .A2(in_a[12]), .ZN(n_0_0_775));
   OR2_X1 i_0_0_1311 (.A1(in_a[9]), .A2(n_0_0_777), .ZN(n_0_0_776));
   NAND2_X1 i_0_0_1312 (.A1(n_0_0_779), .A2(n_0_0_778), .ZN(n_0_0_777));
   NAND2_X1 i_0_0_1313 (.A1(in_a[63]), .A2(in_a[8]), .ZN(n_0_0_778));
   OAI21_X1 i_0_0_1314 (.A(in_a[63]), .B1(n_0_0_781), .B2(in_a[7]), .ZN(
      n_0_0_779));
   NAND2_X1 i_0_0_1315 (.A1(n_0_0_781), .A2(in_a[63]), .ZN(n_0_0_780));
   OR2_X1 i_0_0_1316 (.A1(n_0_0_782), .A2(in_a[6]), .ZN(n_0_0_781));
   NAND2_X1 i_0_0_1317 (.A1(n_0_0_790), .A2(n_0_0_783), .ZN(n_0_0_782));
   OAI21_X1 i_0_0_1318 (.A(in_a[63]), .B1(in_a[4]), .B2(n_0_0_784), .ZN(
      n_0_0_783));
   NAND2_X1 i_0_0_1319 (.A1(n_0_0_786), .A2(n_0_0_785), .ZN(n_0_0_784));
   NAND2_X1 i_0_0_1320 (.A1(in_a[63]), .A2(in_a[3]), .ZN(n_0_0_785));
   AOI21_X1 i_0_0_1321 (.A(n_0_0_787), .B1(in_a[2]), .B2(in_a[63]), .ZN(
      n_0_0_786));
   INV_X1 i_0_0_1322 (.A(n_0_0_788), .ZN(n_0_0_787));
   OAI21_X1 i_0_0_1323 (.A(in_a[63]), .B1(in_a[1]), .B2(in_a[0]), .ZN(n_0_0_788));
   NAND2_X1 i_0_0_1324 (.A1(in_a[63]), .A2(in_a[0]), .ZN(n_0_0_789));
   NAND2_X1 i_0_0_1325 (.A1(in_a[63]), .A2(in_a[5]), .ZN(n_0_0_790));
   INV_X1 i_0_0_1326 (.A(n_0_0_791), .ZN(n_0_391));
   OAI21_X1 i_0_0_1327 (.A(n_0_0_792), .B1(in_b[1]), .B2(in_b[63]), .ZN(
      n_0_0_791));
   NAND2_X1 i_0_0_1328 (.A1(n_0_0_855), .A2(in_b[63]), .ZN(n_0_0_792));
   INV_X1 i_0_0_1329 (.A(n_0_0_793), .ZN(n_0_436));
   OAI21_X1 i_0_0_1330 (.A(n_0_0_794), .B1(n_0_2), .B2(n_0_0_862), .ZN(n_0_0_793));
   OR2_X1 i_0_0_1331 (.A1(in_b[63]), .A2(in_b[2]), .ZN(n_0_0_794));
   INV_X1 i_0_0_1332 (.A(n_0_0_795), .ZN(n_0_481));
   OAI21_X1 i_0_0_1333 (.A(n_0_0_796), .B1(n_0_3), .B2(n_0_0_862), .ZN(n_0_0_795));
   OR2_X1 i_0_0_1334 (.A1(in_b[63]), .A2(in_b[3]), .ZN(n_0_0_796));
   INV_X1 i_0_0_1335 (.A(n_0_0_797), .ZN(n_0_526));
   OAI21_X1 i_0_0_1336 (.A(n_0_0_798), .B1(n_0_4), .B2(n_0_0_862), .ZN(n_0_0_797));
   OR2_X1 i_0_0_1337 (.A1(in_b[63]), .A2(in_b[4]), .ZN(n_0_0_798));
   INV_X1 i_0_0_1338 (.A(n_0_0_799), .ZN(n_0_571));
   OAI21_X1 i_0_0_1339 (.A(n_0_0_800), .B1(n_0_5), .B2(n_0_0_862), .ZN(n_0_0_799));
   OR2_X1 i_0_0_1340 (.A1(in_b[63]), .A2(in_b[5]), .ZN(n_0_0_800));
   INV_X1 i_0_0_1341 (.A(n_0_0_801), .ZN(n_0_616));
   OAI21_X1 i_0_0_1342 (.A(n_0_0_802), .B1(n_0_6), .B2(n_0_0_862), .ZN(n_0_0_801));
   OR2_X1 i_0_0_1343 (.A1(in_b[63]), .A2(in_b[6]), .ZN(n_0_0_802));
   INV_X1 i_0_0_1344 (.A(n_0_0_803), .ZN(n_0_661));
   OAI21_X1 i_0_0_1345 (.A(n_0_0_804), .B1(n_0_7), .B2(n_0_0_862), .ZN(n_0_0_803));
   OR2_X1 i_0_0_1346 (.A1(in_b[63]), .A2(in_b[7]), .ZN(n_0_0_804));
   INV_X1 i_0_0_1347 (.A(n_0_0_805), .ZN(n_0_706));
   OAI21_X1 i_0_0_1348 (.A(n_0_0_806), .B1(n_0_8), .B2(n_0_0_862), .ZN(n_0_0_805));
   OR2_X1 i_0_0_1349 (.A1(in_b[63]), .A2(in_b[8]), .ZN(n_0_0_806));
   INV_X1 i_0_0_1350 (.A(n_0_0_807), .ZN(n_0_751));
   OAI21_X1 i_0_0_1351 (.A(n_0_0_808), .B1(n_0_9), .B2(n_0_0_862), .ZN(n_0_0_807));
   OR2_X1 i_0_0_1352 (.A1(in_b[63]), .A2(in_b[9]), .ZN(n_0_0_808));
   INV_X1 i_0_0_1353 (.A(n_0_0_809), .ZN(n_0_796));
   OAI21_X1 i_0_0_1354 (.A(n_0_0_810), .B1(n_0_10), .B2(n_0_0_862), .ZN(
      n_0_0_809));
   OR2_X1 i_0_0_1355 (.A1(in_b[63]), .A2(in_b[10]), .ZN(n_0_0_810));
   INV_X1 i_0_0_1356 (.A(n_0_0_811), .ZN(n_0_840));
   OAI21_X1 i_0_0_1357 (.A(n_0_0_812), .B1(n_0_11), .B2(n_0_0_862), .ZN(
      n_0_0_811));
   OR2_X1 i_0_0_1358 (.A1(in_b[63]), .A2(in_b[11]), .ZN(n_0_0_812));
   INV_X1 i_0_0_1359 (.A(n_0_0_813), .ZN(n_0_884));
   OAI21_X1 i_0_0_1360 (.A(n_0_0_814), .B1(n_0_12), .B2(n_0_0_862), .ZN(
      n_0_0_813));
   OR2_X1 i_0_0_1361 (.A1(in_b[63]), .A2(in_b[12]), .ZN(n_0_0_814));
   INV_X1 i_0_0_1362 (.A(n_0_0_815), .ZN(n_0_928));
   OAI21_X1 i_0_0_1363 (.A(n_0_0_816), .B1(n_0_13), .B2(n_0_0_862), .ZN(
      n_0_0_815));
   OR2_X1 i_0_0_1364 (.A1(in_b[63]), .A2(in_b[13]), .ZN(n_0_0_816));
   INV_X1 i_0_0_1365 (.A(n_0_0_817), .ZN(n_0_972));
   OAI21_X1 i_0_0_1366 (.A(n_0_0_818), .B1(n_0_14), .B2(n_0_0_862), .ZN(
      n_0_0_817));
   OR2_X1 i_0_0_1367 (.A1(in_b[63]), .A2(in_b[14]), .ZN(n_0_0_818));
   INV_X1 i_0_0_1368 (.A(n_0_0_819), .ZN(n_0_1016));
   OAI21_X1 i_0_0_1369 (.A(n_0_0_820), .B1(n_0_15), .B2(n_0_0_862), .ZN(
      n_0_0_819));
   OR2_X1 i_0_0_1370 (.A1(in_b[63]), .A2(in_b[15]), .ZN(n_0_0_820));
   INV_X1 i_0_0_1371 (.A(n_0_0_821), .ZN(n_0_1017));
   OAI21_X1 i_0_0_1372 (.A(n_0_0_822), .B1(n_0_16), .B2(n_0_0_862), .ZN(
      n_0_0_821));
   OR2_X1 i_0_0_1373 (.A1(in_b[63]), .A2(in_b[16]), .ZN(n_0_0_822));
   INV_X1 i_0_0_1374 (.A(n_0_0_823), .ZN(n_0_1060));
   OAI21_X1 i_0_0_1375 (.A(n_0_0_824), .B1(n_0_17), .B2(n_0_0_862), .ZN(
      n_0_0_823));
   OR2_X1 i_0_0_1376 (.A1(in_b[63]), .A2(in_b[17]), .ZN(n_0_0_824));
   INV_X1 i_0_0_1377 (.A(n_0_0_825), .ZN(n_0_1061));
   OAI21_X1 i_0_0_1378 (.A(n_0_0_826), .B1(n_0_18), .B2(n_0_0_862), .ZN(
      n_0_0_825));
   OR2_X1 i_0_0_1379 (.A1(in_b[63]), .A2(in_b[18]), .ZN(n_0_0_826));
   INV_X1 i_0_0_1380 (.A(n_0_0_827), .ZN(n_0_1062));
   OAI21_X1 i_0_0_1381 (.A(n_0_0_828), .B1(n_0_19), .B2(n_0_0_862), .ZN(
      n_0_0_827));
   OR2_X1 i_0_0_1382 (.A1(in_b[63]), .A2(in_b[19]), .ZN(n_0_0_828));
   INV_X1 i_0_0_1383 (.A(n_0_0_829), .ZN(n_0_1063));
   OAI21_X1 i_0_0_1384 (.A(n_0_0_830), .B1(n_0_20), .B2(n_0_0_862), .ZN(
      n_0_0_829));
   OR2_X1 i_0_0_1385 (.A1(in_b[63]), .A2(in_b[20]), .ZN(n_0_0_830));
   INV_X1 i_0_0_1386 (.A(n_0_0_831), .ZN(n_0_1064));
   OAI21_X1 i_0_0_1387 (.A(n_0_0_832), .B1(n_0_21), .B2(n_0_0_862), .ZN(
      n_0_0_831));
   OR2_X1 i_0_0_1388 (.A1(in_b[63]), .A2(in_b[21]), .ZN(n_0_0_832));
   INV_X1 i_0_0_1389 (.A(rst), .ZN(n_0_39));
   INV_X1 i_0_0_1390 (.A(n_0_36), .ZN(n_0_0_833));
   INV_X1 i_0_0_1391 (.A(n_0_78), .ZN(n_0_0_834));
   INV_X1 i_0_0_1392 (.A(n_0_79), .ZN(n_0_0_835));
   INV_X1 i_0_0_1393 (.A(n_0_80), .ZN(n_0_0_836));
   INV_X1 i_0_0_1394 (.A(n_0_81), .ZN(n_0_0_837));
   INV_X1 i_0_0_1395 (.A(n_0_82), .ZN(n_0_0_838));
   INV_X1 i_0_0_1396 (.A(n_0_83), .ZN(n_0_0_839));
   INV_X1 i_0_0_1397 (.A(n_0_84), .ZN(n_0_0_840));
   INV_X1 i_0_0_1398 (.A(n_0_85), .ZN(n_0_0_841));
   INV_X1 i_0_0_1399 (.A(n_0_86), .ZN(n_0_0_842));
   INV_X1 i_0_0_1400 (.A(n_0_87), .ZN(n_0_0_843));
   INV_X1 i_0_0_1401 (.A(n_0_88), .ZN(n_0_0_844));
   INV_X1 i_0_0_1402 (.A(n_0_89), .ZN(n_0_0_845));
   INV_X1 i_0_0_1403 (.A(n_0_90), .ZN(n_0_0_846));
   INV_X1 i_0_0_1404 (.A(n_0_91), .ZN(n_0_0_847));
   INV_X1 i_0_0_1405 (.A(n_0_92), .ZN(n_0_0_848));
   INV_X1 i_0_0_1406 (.A(n_0_93), .ZN(n_0_0_849));
   INV_X1 i_0_0_1407 (.A(n_0_94), .ZN(n_0_0_850));
   INV_X1 i_0_0_1408 (.A(n_0_95), .ZN(n_0_0_851));
   INV_X1 i_0_0_1409 (.A(n_0_96), .ZN(n_0_0_852));
   INV_X1 i_0_0_1410 (.A(n_0_97), .ZN(n_0_0_853));
   INV_X1 i_0_0_1411 (.A(n_0_98), .ZN(n_0_0_854));
   INV_X1 i_0_0_1412 (.A(n_0_1), .ZN(n_0_0_855));
   INV_X1 i_0_0_1413 (.A(n_0_1042), .ZN(n_0_0_856));
   INV_X1 i_0_0_1414 (.A(n_0_998), .ZN(n_0_0_857));
   INV_X1 i_0_0_1415 (.A(n_0_327), .ZN(n_0_0_858));
   INV_X1 i_0_0_1416 (.A(n_0_282), .ZN(n_0_0_859));
   INV_X1 i_0_0_1417 (.A(n_0_192), .ZN(n_0_0_860));
   INV_X1 i_0_0_1418 (.A(in_b[0]), .ZN(n_0_0_861));
   INV_X1 i_0_0_1419 (.A(in_b[63]), .ZN(n_0_0_862));
endmodule
