/*
 * Created by 
   ../bin/Linux-x86_64-O/oasysGui 19.2-p002 on Sat Apr 25 22:31:16 2020
 * (C) Mentor Graphics Corporation
 */
/* CheckSum: 2796667101 */

module datapath__0_57(R, L, plus);
   input [15:0]R;
   input [15:0]L;
   output [15:0]plus;

   HA_X1 i_1 (.A(R[0]), .B(L[0]), .CO(n_1), .S(plus[0]));
   FA_X1 i_2 (.A(R[1]), .B(L[1]), .CI(n_1), .CO(n_2), .S(plus[1]));
   FA_X1 i_3 (.A(R[2]), .B(L[2]), .CI(n_2), .CO(n_3), .S(plus[2]));
   FA_X1 i_4 (.A(R[3]), .B(L[3]), .CI(n_3), .CO(n_4), .S(plus[3]));
   FA_X1 i_5 (.A(R[4]), .B(L[4]), .CI(n_4), .CO(n_5), .S(plus[4]));
   FA_X1 i_6 (.A(R[5]), .B(L[5]), .CI(n_5), .CO(n_6), .S(plus[5]));
   FA_X1 i_7 (.A(R[6]), .B(L[6]), .CI(n_6), .CO(n_7), .S(plus[6]));
   FA_X1 i_8 (.A(R[7]), .B(L[7]), .CI(n_7), .CO(n_8), .S(plus[7]));
   FA_X1 i_9 (.A(R[8]), .B(L[8]), .CI(n_8), .CO(n_9), .S(plus[8]));
   FA_X1 i_10 (.A(R[9]), .B(L[9]), .CI(n_9), .CO(n_10), .S(plus[9]));
   FA_X1 i_11 (.A(R[10]), .B(L[10]), .CI(n_10), .CO(n_11), .S(plus[10]));
   FA_X1 i_12 (.A(R[11]), .B(L[11]), .CI(n_11), .CO(n_12), .S(plus[11]));
   FA_X1 i_13 (.A(R[12]), .B(L[12]), .CI(n_12), .CO(n_13), .S(plus[12]));
   FA_X1 i_14 (.A(R[13]), .B(L[13]), .CI(n_13), .CO(n_14), .S(plus[13]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(plus[14]));
   OAI22_X1 i_15 (.A1(n_18), .A2(L[14]), .B1(R[14]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(R[15]), .B(n_15), .Z(plus[15]));
   OAI33_X1 i_17 (.A1(n_18), .A2(L[14]), .A3(n_16), .B1(R[14]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(L[14]), .ZN(n_17));
   INV_X1 i_20 (.A(R[14]), .ZN(n_18));
endmodule

module datapath__0_60(minus, L, p_0);
   input [15:0]minus;
   input [15:0]L;
   output [15:0]p_0;

   HA_X1 i_1 (.A(minus[0]), .B(L[0]), .CO(n_1), .S(p_0[0]));
   FA_X1 i_2 (.A(minus[1]), .B(L[1]), .CI(n_1), .CO(n_2), .S(p_0[1]));
   FA_X1 i_3 (.A(minus[2]), .B(L[2]), .CI(n_2), .CO(n_3), .S(p_0[2]));
   FA_X1 i_4 (.A(minus[3]), .B(L[3]), .CI(n_3), .CO(n_4), .S(p_0[3]));
   FA_X1 i_5 (.A(minus[4]), .B(L[4]), .CI(n_4), .CO(n_5), .S(p_0[4]));
   FA_X1 i_6 (.A(minus[5]), .B(L[5]), .CI(n_5), .CO(n_6), .S(p_0[5]));
   FA_X1 i_7 (.A(minus[6]), .B(L[6]), .CI(n_6), .CO(n_7), .S(p_0[6]));
   FA_X1 i_8 (.A(minus[7]), .B(L[7]), .CI(n_7), .CO(n_8), .S(p_0[7]));
   FA_X1 i_9 (.A(minus[8]), .B(L[8]), .CI(n_8), .CO(n_9), .S(p_0[8]));
   FA_X1 i_10 (.A(minus[9]), .B(L[9]), .CI(n_9), .CO(n_10), .S(p_0[9]));
   FA_X1 i_11 (.A(minus[10]), .B(L[10]), .CI(n_10), .CO(n_11), .S(p_0[10]));
   FA_X1 i_12 (.A(minus[11]), .B(L[11]), .CI(n_11), .CO(n_12), .S(p_0[11]));
   FA_X1 i_13 (.A(minus[12]), .B(L[12]), .CI(n_12), .CO(n_13), .S(p_0[12]));
   FA_X1 i_14 (.A(minus[13]), .B(L[13]), .CI(n_13), .CO(n_14), .S(p_0[13]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_0[14]));
   OAI22_X1 i_15 (.A1(n_18), .A2(L[14]), .B1(minus[14]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(minus[15]), .B(n_15), .Z(p_0[15]));
   OAI33_X1 i_17 (.A1(n_18), .A2(L[14]), .A3(n_16), .B1(minus[14]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(L[14]), .ZN(n_17));
   INV_X1 i_20 (.A(minus[14]), .ZN(n_18));
endmodule

module datapath__0_65(R, L, plus);
   input [15:0]R;
   input [15:0]L;
   output [15:0]plus;

   HA_X1 i_1 (.A(R[0]), .B(L[0]), .CO(n_1), .S(plus[0]));
   FA_X1 i_2 (.A(R[1]), .B(L[1]), .CI(n_1), .CO(n_2), .S(plus[1]));
   FA_X1 i_3 (.A(R[2]), .B(L[2]), .CI(n_2), .CO(n_3), .S(plus[2]));
   FA_X1 i_4 (.A(R[3]), .B(L[3]), .CI(n_3), .CO(n_4), .S(plus[3]));
   FA_X1 i_5 (.A(R[4]), .B(L[4]), .CI(n_4), .CO(n_5), .S(plus[4]));
   FA_X1 i_6 (.A(R[5]), .B(L[5]), .CI(n_5), .CO(n_6), .S(plus[5]));
   FA_X1 i_7 (.A(R[6]), .B(L[6]), .CI(n_6), .CO(n_7), .S(plus[6]));
   FA_X1 i_8 (.A(R[7]), .B(L[7]), .CI(n_7), .CO(n_8), .S(plus[7]));
   FA_X1 i_9 (.A(R[8]), .B(L[8]), .CI(n_8), .CO(n_9), .S(plus[8]));
   FA_X1 i_10 (.A(R[9]), .B(L[9]), .CI(n_9), .CO(n_10), .S(plus[9]));
   FA_X1 i_11 (.A(R[10]), .B(L[10]), .CI(n_10), .CO(n_11), .S(plus[10]));
   FA_X1 i_12 (.A(R[11]), .B(L[11]), .CI(n_11), .CO(n_12), .S(plus[11]));
   FA_X1 i_13 (.A(R[12]), .B(L[12]), .CI(n_12), .CO(n_13), .S(plus[12]));
   FA_X1 i_14 (.A(R[13]), .B(L[13]), .CI(n_13), .CO(n_14), .S(plus[13]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(plus[14]));
   OAI22_X1 i_15 (.A1(n_18), .A2(L[14]), .B1(R[14]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(R[15]), .B(n_15), .Z(plus[15]));
   OAI33_X1 i_17 (.A1(n_18), .A2(L[14]), .A3(n_16), .B1(R[14]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(L[14]), .ZN(n_17));
   INV_X1 i_20 (.A(R[14]), .ZN(n_18));
endmodule

module datapath__0_68(minus, L, p_0);
   input [15:0]minus;
   input [15:0]L;
   output [15:0]p_0;

   HA_X1 i_1 (.A(minus[0]), .B(L[0]), .CO(n_1), .S(p_0[0]));
   FA_X1 i_2 (.A(minus[1]), .B(L[1]), .CI(n_1), .CO(n_2), .S(p_0[1]));
   FA_X1 i_3 (.A(minus[2]), .B(L[2]), .CI(n_2), .CO(n_3), .S(p_0[2]));
   FA_X1 i_4 (.A(minus[3]), .B(L[3]), .CI(n_3), .CO(n_4), .S(p_0[3]));
   FA_X1 i_5 (.A(minus[4]), .B(L[4]), .CI(n_4), .CO(n_5), .S(p_0[4]));
   FA_X1 i_6 (.A(minus[5]), .B(L[5]), .CI(n_5), .CO(n_6), .S(p_0[5]));
   FA_X1 i_7 (.A(minus[6]), .B(L[6]), .CI(n_6), .CO(n_7), .S(p_0[6]));
   FA_X1 i_8 (.A(minus[7]), .B(L[7]), .CI(n_7), .CO(n_8), .S(p_0[7]));
   FA_X1 i_9 (.A(minus[8]), .B(L[8]), .CI(n_8), .CO(n_9), .S(p_0[8]));
   FA_X1 i_10 (.A(minus[9]), .B(L[9]), .CI(n_9), .CO(n_10), .S(p_0[9]));
   FA_X1 i_11 (.A(minus[10]), .B(L[10]), .CI(n_10), .CO(n_11), .S(p_0[10]));
   FA_X1 i_12 (.A(minus[11]), .B(L[11]), .CI(n_11), .CO(n_12), .S(p_0[11]));
   FA_X1 i_13 (.A(minus[12]), .B(L[12]), .CI(n_12), .CO(n_13), .S(p_0[12]));
   FA_X1 i_14 (.A(minus[13]), .B(L[13]), .CI(n_13), .CO(n_14), .S(p_0[13]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_0[14]));
   OAI22_X1 i_15 (.A1(n_18), .A2(L[14]), .B1(minus[14]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(minus[15]), .B(n_15), .Z(p_0[15]));
   OAI33_X1 i_17 (.A1(n_18), .A2(L[14]), .A3(n_16), .B1(minus[14]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(L[14]), .ZN(n_17));
   INV_X1 i_20 (.A(minus[14]), .ZN(n_18));
endmodule

module datapath__0_73(R, L, plus);
   input [15:0]R;
   input [15:0]L;
   output [15:0]plus;

   HA_X1 i_1 (.A(R[0]), .B(L[0]), .CO(n_1), .S(plus[0]));
   FA_X1 i_2 (.A(R[1]), .B(L[1]), .CI(n_1), .CO(n_2), .S(plus[1]));
   FA_X1 i_3 (.A(R[2]), .B(L[2]), .CI(n_2), .CO(n_3), .S(plus[2]));
   FA_X1 i_4 (.A(R[3]), .B(L[3]), .CI(n_3), .CO(n_4), .S(plus[3]));
   FA_X1 i_5 (.A(R[4]), .B(L[4]), .CI(n_4), .CO(n_5), .S(plus[4]));
   FA_X1 i_6 (.A(R[5]), .B(L[5]), .CI(n_5), .CO(n_6), .S(plus[5]));
   FA_X1 i_7 (.A(R[6]), .B(L[6]), .CI(n_6), .CO(n_7), .S(plus[6]));
   FA_X1 i_8 (.A(R[7]), .B(L[7]), .CI(n_7), .CO(n_8), .S(plus[7]));
   FA_X1 i_9 (.A(R[8]), .B(L[8]), .CI(n_8), .CO(n_9), .S(plus[8]));
   FA_X1 i_10 (.A(R[9]), .B(L[9]), .CI(n_9), .CO(n_10), .S(plus[9]));
   FA_X1 i_11 (.A(R[10]), .B(L[10]), .CI(n_10), .CO(n_11), .S(plus[10]));
   FA_X1 i_12 (.A(R[11]), .B(L[11]), .CI(n_11), .CO(n_12), .S(plus[11]));
   FA_X1 i_13 (.A(R[12]), .B(L[12]), .CI(n_12), .CO(n_13), .S(plus[12]));
   FA_X1 i_14 (.A(R[13]), .B(L[13]), .CI(n_13), .CO(n_14), .S(plus[13]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(plus[14]));
   OAI22_X1 i_15 (.A1(n_18), .A2(L[14]), .B1(R[14]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(R[15]), .B(n_15), .Z(plus[15]));
   OAI33_X1 i_17 (.A1(n_18), .A2(L[14]), .A3(n_16), .B1(R[14]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(L[14]), .ZN(n_17));
   INV_X1 i_20 (.A(R[14]), .ZN(n_18));
endmodule

module datapath__0_76(minus, L, p_0);
   input [15:0]minus;
   input [15:0]L;
   output [15:0]p_0;

   HA_X1 i_1 (.A(minus[0]), .B(L[0]), .CO(n_1), .S(p_0[0]));
   FA_X1 i_2 (.A(minus[1]), .B(L[1]), .CI(n_1), .CO(n_2), .S(p_0[1]));
   FA_X1 i_3 (.A(minus[2]), .B(L[2]), .CI(n_2), .CO(n_3), .S(p_0[2]));
   FA_X1 i_4 (.A(minus[3]), .B(L[3]), .CI(n_3), .CO(n_4), .S(p_0[3]));
   FA_X1 i_5 (.A(minus[4]), .B(L[4]), .CI(n_4), .CO(n_5), .S(p_0[4]));
   FA_X1 i_6 (.A(minus[5]), .B(L[5]), .CI(n_5), .CO(n_6), .S(p_0[5]));
   FA_X1 i_7 (.A(minus[6]), .B(L[6]), .CI(n_6), .CO(n_7), .S(p_0[6]));
   FA_X1 i_8 (.A(minus[7]), .B(L[7]), .CI(n_7), .CO(n_8), .S(p_0[7]));
   FA_X1 i_9 (.A(minus[8]), .B(L[8]), .CI(n_8), .CO(n_9), .S(p_0[8]));
   FA_X1 i_10 (.A(minus[9]), .B(L[9]), .CI(n_9), .CO(n_10), .S(p_0[9]));
   FA_X1 i_11 (.A(minus[10]), .B(L[10]), .CI(n_10), .CO(n_11), .S(p_0[10]));
   FA_X1 i_12 (.A(minus[11]), .B(L[11]), .CI(n_11), .CO(n_12), .S(p_0[11]));
   FA_X1 i_13 (.A(minus[12]), .B(L[12]), .CI(n_12), .CO(n_13), .S(p_0[12]));
   FA_X1 i_14 (.A(minus[13]), .B(L[13]), .CI(n_13), .CO(n_14), .S(p_0[13]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_0[14]));
   OAI22_X1 i_15 (.A1(n_18), .A2(L[14]), .B1(minus[14]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(minus[15]), .B(n_15), .Z(p_0[15]));
   OAI33_X1 i_17 (.A1(n_18), .A2(L[14]), .A3(n_16), .B1(minus[14]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(L[14]), .ZN(n_17));
   INV_X1 i_20 (.A(minus[14]), .ZN(n_18));
endmodule

module datapath__0_81(R, L, plus);
   input [15:0]R;
   input [15:0]L;
   output [15:0]plus;

   HA_X1 i_1 (.A(R[0]), .B(L[0]), .CO(n_1), .S(plus[0]));
   FA_X1 i_2 (.A(R[1]), .B(L[1]), .CI(n_1), .CO(n_2), .S(plus[1]));
   FA_X1 i_3 (.A(R[2]), .B(L[2]), .CI(n_2), .CO(n_3), .S(plus[2]));
   FA_X1 i_4 (.A(R[3]), .B(L[3]), .CI(n_3), .CO(n_4), .S(plus[3]));
   FA_X1 i_5 (.A(R[4]), .B(L[4]), .CI(n_4), .CO(n_5), .S(plus[4]));
   FA_X1 i_6 (.A(R[5]), .B(L[5]), .CI(n_5), .CO(n_6), .S(plus[5]));
   FA_X1 i_7 (.A(R[6]), .B(L[6]), .CI(n_6), .CO(n_7), .S(plus[6]));
   FA_X1 i_8 (.A(R[7]), .B(L[7]), .CI(n_7), .CO(n_8), .S(plus[7]));
   FA_X1 i_9 (.A(R[8]), .B(L[8]), .CI(n_8), .CO(n_9), .S(plus[8]));
   FA_X1 i_10 (.A(R[9]), .B(L[9]), .CI(n_9), .CO(n_10), .S(plus[9]));
   FA_X1 i_11 (.A(R[10]), .B(L[10]), .CI(n_10), .CO(n_11), .S(plus[10]));
   FA_X1 i_12 (.A(R[11]), .B(L[11]), .CI(n_11), .CO(n_12), .S(plus[11]));
   FA_X1 i_13 (.A(R[12]), .B(L[12]), .CI(n_12), .CO(n_13), .S(plus[12]));
   FA_X1 i_14 (.A(R[13]), .B(L[13]), .CI(n_13), .CO(n_14), .S(plus[13]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(plus[14]));
   OAI22_X1 i_15 (.A1(n_18), .A2(L[14]), .B1(R[14]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(R[15]), .B(n_15), .Z(plus[15]));
   OAI33_X1 i_17 (.A1(n_18), .A2(L[14]), .A3(n_16), .B1(R[14]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(L[14]), .ZN(n_17));
   INV_X1 i_20 (.A(R[14]), .ZN(n_18));
endmodule

module datapath__0_84(minus, L, p_0);
   input [15:0]minus;
   input [15:0]L;
   output [15:0]p_0;

   HA_X1 i_1 (.A(minus[0]), .B(L[0]), .CO(n_1), .S(p_0[0]));
   FA_X1 i_2 (.A(minus[1]), .B(L[1]), .CI(n_1), .CO(n_2), .S(p_0[1]));
   FA_X1 i_3 (.A(minus[2]), .B(L[2]), .CI(n_2), .CO(n_3), .S(p_0[2]));
   FA_X1 i_4 (.A(minus[3]), .B(L[3]), .CI(n_3), .CO(n_4), .S(p_0[3]));
   FA_X1 i_5 (.A(minus[4]), .B(L[4]), .CI(n_4), .CO(n_5), .S(p_0[4]));
   FA_X1 i_6 (.A(minus[5]), .B(L[5]), .CI(n_5), .CO(n_6), .S(p_0[5]));
   FA_X1 i_7 (.A(minus[6]), .B(L[6]), .CI(n_6), .CO(n_7), .S(p_0[6]));
   FA_X1 i_8 (.A(minus[7]), .B(L[7]), .CI(n_7), .CO(n_8), .S(p_0[7]));
   FA_X1 i_9 (.A(minus[8]), .B(L[8]), .CI(n_8), .CO(n_9), .S(p_0[8]));
   FA_X1 i_10 (.A(minus[9]), .B(L[9]), .CI(n_9), .CO(n_10), .S(p_0[9]));
   FA_X1 i_11 (.A(minus[10]), .B(L[10]), .CI(n_10), .CO(n_11), .S(p_0[10]));
   FA_X1 i_12 (.A(minus[11]), .B(L[11]), .CI(n_11), .CO(n_12), .S(p_0[11]));
   FA_X1 i_13 (.A(minus[12]), .B(L[12]), .CI(n_12), .CO(n_13), .S(p_0[12]));
   FA_X1 i_14 (.A(minus[13]), .B(L[13]), .CI(n_13), .CO(n_14), .S(p_0[13]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_0[14]));
   OAI22_X1 i_15 (.A1(n_18), .A2(L[14]), .B1(minus[14]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(minus[15]), .B(n_15), .Z(p_0[15]));
   OAI33_X1 i_17 (.A1(n_18), .A2(L[14]), .A3(n_16), .B1(minus[14]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(L[14]), .ZN(n_17));
   INV_X1 i_20 (.A(minus[14]), .ZN(n_18));
endmodule

module datapath__0_89(R, L, plus);
   input [15:0]R;
   input [15:0]L;
   output [15:0]plus;

   HA_X1 i_1 (.A(R[0]), .B(L[0]), .CO(n_1), .S(plus[0]));
   FA_X1 i_2 (.A(R[1]), .B(L[1]), .CI(n_1), .CO(n_2), .S(plus[1]));
   FA_X1 i_3 (.A(R[2]), .B(L[2]), .CI(n_2), .CO(n_3), .S(plus[2]));
   FA_X1 i_4 (.A(R[3]), .B(L[3]), .CI(n_3), .CO(n_4), .S(plus[3]));
   FA_X1 i_5 (.A(R[4]), .B(L[4]), .CI(n_4), .CO(n_5), .S(plus[4]));
   FA_X1 i_6 (.A(R[5]), .B(L[5]), .CI(n_5), .CO(n_6), .S(plus[5]));
   FA_X1 i_7 (.A(R[6]), .B(L[6]), .CI(n_6), .CO(n_7), .S(plus[6]));
   FA_X1 i_8 (.A(R[7]), .B(L[7]), .CI(n_7), .CO(n_8), .S(plus[7]));
   FA_X1 i_9 (.A(R[8]), .B(L[8]), .CI(n_8), .CO(n_9), .S(plus[8]));
   FA_X1 i_10 (.A(R[9]), .B(L[9]), .CI(n_9), .CO(n_10), .S(plus[9]));
   FA_X1 i_11 (.A(R[10]), .B(L[10]), .CI(n_10), .CO(n_11), .S(plus[10]));
   FA_X1 i_12 (.A(R[11]), .B(L[11]), .CI(n_11), .CO(n_12), .S(plus[11]));
   FA_X1 i_13 (.A(R[12]), .B(L[12]), .CI(n_12), .CO(n_13), .S(plus[12]));
   FA_X1 i_14 (.A(R[13]), .B(L[13]), .CI(n_13), .CO(n_14), .S(plus[13]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(plus[14]));
   OAI22_X1 i_15 (.A1(n_18), .A2(L[14]), .B1(R[14]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(R[15]), .B(n_15), .Z(plus[15]));
   OAI33_X1 i_17 (.A1(n_18), .A2(L[14]), .A3(n_16), .B1(R[14]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(L[14]), .ZN(n_17));
   INV_X1 i_20 (.A(R[14]), .ZN(n_18));
endmodule

module datapath__0_92(minus, L, p_0);
   input [15:0]minus;
   input [15:0]L;
   output [15:0]p_0;

   HA_X1 i_1 (.A(minus[0]), .B(L[0]), .CO(n_1), .S(p_0[0]));
   FA_X1 i_2 (.A(minus[1]), .B(L[1]), .CI(n_1), .CO(n_2), .S(p_0[1]));
   FA_X1 i_3 (.A(minus[2]), .B(L[2]), .CI(n_2), .CO(n_3), .S(p_0[2]));
   FA_X1 i_4 (.A(minus[3]), .B(L[3]), .CI(n_3), .CO(n_4), .S(p_0[3]));
   FA_X1 i_5 (.A(minus[4]), .B(L[4]), .CI(n_4), .CO(n_5), .S(p_0[4]));
   FA_X1 i_6 (.A(minus[5]), .B(L[5]), .CI(n_5), .CO(n_6), .S(p_0[5]));
   FA_X1 i_7 (.A(minus[6]), .B(L[6]), .CI(n_6), .CO(n_7), .S(p_0[6]));
   FA_X1 i_8 (.A(minus[7]), .B(L[7]), .CI(n_7), .CO(n_8), .S(p_0[7]));
   FA_X1 i_9 (.A(minus[8]), .B(L[8]), .CI(n_8), .CO(n_9), .S(p_0[8]));
   FA_X1 i_10 (.A(minus[9]), .B(L[9]), .CI(n_9), .CO(n_10), .S(p_0[9]));
   FA_X1 i_11 (.A(minus[10]), .B(L[10]), .CI(n_10), .CO(n_11), .S(p_0[10]));
   FA_X1 i_12 (.A(minus[11]), .B(L[11]), .CI(n_11), .CO(n_12), .S(p_0[11]));
   FA_X1 i_13 (.A(minus[12]), .B(L[12]), .CI(n_12), .CO(n_13), .S(p_0[12]));
   FA_X1 i_14 (.A(minus[13]), .B(L[13]), .CI(n_13), .CO(n_14), .S(p_0[13]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_0[14]));
   OAI22_X1 i_15 (.A1(n_18), .A2(L[14]), .B1(minus[14]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(minus[15]), .B(n_15), .Z(p_0[15]));
   OAI33_X1 i_17 (.A1(n_18), .A2(L[14]), .A3(n_16), .B1(minus[14]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(L[14]), .ZN(n_17));
   INV_X1 i_20 (.A(minus[14]), .ZN(n_18));
endmodule

module datapath__0_97(R, L, plus);
   input [15:0]R;
   input [15:0]L;
   output [15:0]plus;

   HA_X1 i_1 (.A(R[0]), .B(L[0]), .CO(n_1), .S(plus[0]));
   FA_X1 i_2 (.A(R[1]), .B(L[1]), .CI(n_1), .CO(n_2), .S(plus[1]));
   FA_X1 i_3 (.A(R[2]), .B(L[2]), .CI(n_2), .CO(n_3), .S(plus[2]));
   FA_X1 i_4 (.A(R[3]), .B(L[3]), .CI(n_3), .CO(n_4), .S(plus[3]));
   FA_X1 i_5 (.A(R[4]), .B(L[4]), .CI(n_4), .CO(n_5), .S(plus[4]));
   FA_X1 i_6 (.A(R[5]), .B(L[5]), .CI(n_5), .CO(n_6), .S(plus[5]));
   FA_X1 i_7 (.A(R[6]), .B(L[6]), .CI(n_6), .CO(n_7), .S(plus[6]));
   FA_X1 i_8 (.A(R[7]), .B(L[7]), .CI(n_7), .CO(n_8), .S(plus[7]));
   FA_X1 i_9 (.A(R[8]), .B(L[8]), .CI(n_8), .CO(n_9), .S(plus[8]));
   FA_X1 i_10 (.A(R[9]), .B(L[9]), .CI(n_9), .CO(n_10), .S(plus[9]));
   FA_X1 i_11 (.A(R[10]), .B(L[10]), .CI(n_10), .CO(n_11), .S(plus[10]));
   FA_X1 i_12 (.A(R[11]), .B(L[11]), .CI(n_11), .CO(n_12), .S(plus[11]));
   FA_X1 i_13 (.A(R[12]), .B(L[12]), .CI(n_12), .CO(n_13), .S(plus[12]));
   FA_X1 i_14 (.A(R[13]), .B(L[13]), .CI(n_13), .CO(n_14), .S(plus[13]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(plus[14]));
   OAI22_X1 i_15 (.A1(n_18), .A2(L[14]), .B1(R[14]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(R[15]), .B(n_15), .Z(plus[15]));
   OAI33_X1 i_17 (.A1(n_18), .A2(L[14]), .A3(n_16), .B1(R[14]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(L[14]), .ZN(n_17));
   INV_X1 i_20 (.A(R[14]), .ZN(n_18));
endmodule

module datapath__0_100(minus, L, p_0);
   input [15:0]minus;
   input [15:0]L;
   output [15:0]p_0;

   HA_X1 i_1 (.A(minus[0]), .B(L[0]), .CO(n_1), .S(p_0[0]));
   FA_X1 i_2 (.A(minus[1]), .B(L[1]), .CI(n_1), .CO(n_2), .S(p_0[1]));
   FA_X1 i_3 (.A(minus[2]), .B(L[2]), .CI(n_2), .CO(n_3), .S(p_0[2]));
   FA_X1 i_4 (.A(minus[3]), .B(L[3]), .CI(n_3), .CO(n_4), .S(p_0[3]));
   FA_X1 i_5 (.A(minus[4]), .B(L[4]), .CI(n_4), .CO(n_5), .S(p_0[4]));
   FA_X1 i_6 (.A(minus[5]), .B(L[5]), .CI(n_5), .CO(n_6), .S(p_0[5]));
   FA_X1 i_7 (.A(minus[6]), .B(L[6]), .CI(n_6), .CO(n_7), .S(p_0[6]));
   FA_X1 i_8 (.A(minus[7]), .B(L[7]), .CI(n_7), .CO(n_8), .S(p_0[7]));
   FA_X1 i_9 (.A(minus[8]), .B(L[8]), .CI(n_8), .CO(n_9), .S(p_0[8]));
   FA_X1 i_10 (.A(minus[9]), .B(L[9]), .CI(n_9), .CO(n_10), .S(p_0[9]));
   FA_X1 i_11 (.A(minus[10]), .B(L[10]), .CI(n_10), .CO(n_11), .S(p_0[10]));
   FA_X1 i_12 (.A(minus[11]), .B(L[11]), .CI(n_11), .CO(n_12), .S(p_0[11]));
   FA_X1 i_13 (.A(minus[12]), .B(L[12]), .CI(n_12), .CO(n_13), .S(p_0[12]));
   FA_X1 i_14 (.A(minus[13]), .B(L[13]), .CI(n_13), .CO(n_14), .S(p_0[13]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_0[14]));
   OAI22_X1 i_15 (.A1(n_18), .A2(L[14]), .B1(minus[14]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(minus[15]), .B(n_15), .Z(p_0[15]));
   OAI33_X1 i_17 (.A1(n_18), .A2(L[14]), .A3(n_16), .B1(minus[14]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(L[14]), .ZN(n_17));
   INV_X1 i_20 (.A(minus[14]), .ZN(n_18));
endmodule

module datapath__0_105(R, L, plus);
   input [15:0]R;
   input [15:0]L;
   output [15:0]plus;

   HA_X1 i_1 (.A(R[0]), .B(L[0]), .CO(n_1), .S(plus[0]));
   FA_X1 i_2 (.A(R[1]), .B(L[1]), .CI(n_1), .CO(n_2), .S(plus[1]));
   FA_X1 i_3 (.A(R[2]), .B(L[2]), .CI(n_2), .CO(n_3), .S(plus[2]));
   FA_X1 i_4 (.A(R[3]), .B(L[3]), .CI(n_3), .CO(n_4), .S(plus[3]));
   FA_X1 i_5 (.A(R[4]), .B(L[4]), .CI(n_4), .CO(n_5), .S(plus[4]));
   FA_X1 i_6 (.A(R[5]), .B(L[5]), .CI(n_5), .CO(n_6), .S(plus[5]));
   FA_X1 i_7 (.A(R[6]), .B(L[6]), .CI(n_6), .CO(n_7), .S(plus[6]));
   FA_X1 i_8 (.A(R[7]), .B(L[7]), .CI(n_7), .CO(n_8), .S(plus[7]));
   FA_X1 i_9 (.A(R[8]), .B(L[8]), .CI(n_8), .CO(n_9), .S(plus[8]));
   FA_X1 i_10 (.A(R[9]), .B(L[9]), .CI(n_9), .CO(n_10), .S(plus[9]));
   FA_X1 i_11 (.A(R[10]), .B(L[10]), .CI(n_10), .CO(n_11), .S(plus[10]));
   FA_X1 i_12 (.A(R[11]), .B(L[11]), .CI(n_11), .CO(n_12), .S(plus[11]));
   FA_X1 i_13 (.A(R[12]), .B(L[12]), .CI(n_12), .CO(n_13), .S(plus[12]));
   FA_X1 i_14 (.A(R[13]), .B(L[13]), .CI(n_13), .CO(n_14), .S(plus[13]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(plus[14]));
   OAI22_X1 i_15 (.A1(n_18), .A2(L[14]), .B1(R[14]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(R[15]), .B(n_15), .Z(plus[15]));
   OAI33_X1 i_17 (.A1(n_18), .A2(L[14]), .A3(n_16), .B1(R[14]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(L[14]), .ZN(n_17));
   INV_X1 i_20 (.A(R[14]), .ZN(n_18));
endmodule

module datapath__0_108(minus, L, p_0);
   input [15:0]minus;
   input [15:0]L;
   output [15:0]p_0;

   HA_X1 i_1 (.A(minus[0]), .B(L[0]), .CO(n_1), .S(p_0[0]));
   FA_X1 i_2 (.A(minus[1]), .B(L[1]), .CI(n_1), .CO(n_2), .S(p_0[1]));
   FA_X1 i_3 (.A(minus[2]), .B(L[2]), .CI(n_2), .CO(n_3), .S(p_0[2]));
   FA_X1 i_4 (.A(minus[3]), .B(L[3]), .CI(n_3), .CO(n_4), .S(p_0[3]));
   FA_X1 i_5 (.A(minus[4]), .B(L[4]), .CI(n_4), .CO(n_5), .S(p_0[4]));
   FA_X1 i_6 (.A(minus[5]), .B(L[5]), .CI(n_5), .CO(n_6), .S(p_0[5]));
   FA_X1 i_7 (.A(minus[6]), .B(L[6]), .CI(n_6), .CO(n_7), .S(p_0[6]));
   FA_X1 i_8 (.A(minus[7]), .B(L[7]), .CI(n_7), .CO(n_8), .S(p_0[7]));
   FA_X1 i_9 (.A(minus[8]), .B(L[8]), .CI(n_8), .CO(n_9), .S(p_0[8]));
   FA_X1 i_10 (.A(minus[9]), .B(L[9]), .CI(n_9), .CO(n_10), .S(p_0[9]));
   FA_X1 i_11 (.A(minus[10]), .B(L[10]), .CI(n_10), .CO(n_11), .S(p_0[10]));
   FA_X1 i_12 (.A(minus[11]), .B(L[11]), .CI(n_11), .CO(n_12), .S(p_0[11]));
   FA_X1 i_13 (.A(minus[12]), .B(L[12]), .CI(n_12), .CO(n_13), .S(p_0[12]));
   FA_X1 i_14 (.A(minus[13]), .B(L[13]), .CI(n_13), .CO(n_14), .S(p_0[13]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_0[14]));
   OAI22_X1 i_15 (.A1(n_18), .A2(L[14]), .B1(minus[14]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(minus[15]), .B(n_15), .Z(p_0[15]));
   OAI33_X1 i_17 (.A1(n_18), .A2(L[14]), .A3(n_16), .B1(minus[14]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(L[14]), .ZN(n_17));
   INV_X1 i_20 (.A(minus[14]), .ZN(n_18));
endmodule

module datapath__0_113(R, L, plus);
   input [15:0]R;
   input [15:0]L;
   output [15:0]plus;

   HA_X1 i_1 (.A(R[0]), .B(L[0]), .CO(n_1), .S(plus[0]));
   FA_X1 i_2 (.A(R[1]), .B(L[1]), .CI(n_1), .CO(n_2), .S(plus[1]));
   FA_X1 i_3 (.A(R[2]), .B(L[2]), .CI(n_2), .CO(n_3), .S(plus[2]));
   FA_X1 i_4 (.A(R[3]), .B(L[3]), .CI(n_3), .CO(n_4), .S(plus[3]));
   FA_X1 i_5 (.A(R[4]), .B(L[4]), .CI(n_4), .CO(n_5), .S(plus[4]));
   FA_X1 i_6 (.A(R[5]), .B(L[5]), .CI(n_5), .CO(n_6), .S(plus[5]));
   FA_X1 i_7 (.A(R[6]), .B(L[6]), .CI(n_6), .CO(n_7), .S(plus[6]));
   FA_X1 i_8 (.A(R[7]), .B(L[7]), .CI(n_7), .CO(n_8), .S(plus[7]));
   FA_X1 i_9 (.A(R[8]), .B(L[8]), .CI(n_8), .CO(n_9), .S(plus[8]));
   FA_X1 i_10 (.A(R[9]), .B(L[9]), .CI(n_9), .CO(n_10), .S(plus[9]));
   FA_X1 i_11 (.A(R[10]), .B(L[10]), .CI(n_10), .CO(n_11), .S(plus[10]));
   FA_X1 i_12 (.A(R[11]), .B(L[11]), .CI(n_11), .CO(n_12), .S(plus[11]));
   FA_X1 i_13 (.A(R[12]), .B(L[12]), .CI(n_12), .CO(n_13), .S(plus[12]));
   FA_X1 i_14 (.A(R[13]), .B(L[13]), .CI(n_13), .CO(n_14), .S(plus[13]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(plus[14]));
   OAI22_X1 i_15 (.A1(n_18), .A2(L[14]), .B1(R[14]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(R[15]), .B(n_15), .Z(plus[15]));
   OAI33_X1 i_17 (.A1(n_18), .A2(L[14]), .A3(n_16), .B1(R[14]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(L[14]), .ZN(n_17));
   INV_X1 i_20 (.A(R[14]), .ZN(n_18));
endmodule

module datapath__0_116(minus, L, p_0);
   input [15:0]minus;
   input [15:0]L;
   output [15:0]p_0;

   HA_X1 i_1 (.A(minus[0]), .B(L[0]), .CO(n_1), .S(p_0[0]));
   FA_X1 i_2 (.A(minus[1]), .B(L[1]), .CI(n_1), .CO(n_2), .S(p_0[1]));
   FA_X1 i_3 (.A(minus[2]), .B(L[2]), .CI(n_2), .CO(n_3), .S(p_0[2]));
   FA_X1 i_4 (.A(minus[3]), .B(L[3]), .CI(n_3), .CO(n_4), .S(p_0[3]));
   FA_X1 i_5 (.A(minus[4]), .B(L[4]), .CI(n_4), .CO(n_5), .S(p_0[4]));
   FA_X1 i_6 (.A(minus[5]), .B(L[5]), .CI(n_5), .CO(n_6), .S(p_0[5]));
   FA_X1 i_7 (.A(minus[6]), .B(L[6]), .CI(n_6), .CO(n_7), .S(p_0[6]));
   FA_X1 i_8 (.A(minus[7]), .B(L[7]), .CI(n_7), .CO(n_8), .S(p_0[7]));
   FA_X1 i_9 (.A(minus[8]), .B(L[8]), .CI(n_8), .CO(n_9), .S(p_0[8]));
   FA_X1 i_10 (.A(minus[9]), .B(L[9]), .CI(n_9), .CO(n_10), .S(p_0[9]));
   FA_X1 i_11 (.A(minus[10]), .B(L[10]), .CI(n_10), .CO(n_11), .S(p_0[10]));
   FA_X1 i_12 (.A(minus[11]), .B(L[11]), .CI(n_11), .CO(n_12), .S(p_0[11]));
   FA_X1 i_13 (.A(minus[12]), .B(L[12]), .CI(n_12), .CO(n_13), .S(p_0[12]));
   FA_X1 i_14 (.A(minus[13]), .B(L[13]), .CI(n_13), .CO(n_14), .S(p_0[13]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_0[14]));
   OAI22_X1 i_15 (.A1(n_18), .A2(L[14]), .B1(minus[14]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(minus[15]), .B(n_15), .Z(p_0[15]));
   OAI33_X1 i_17 (.A1(n_18), .A2(L[14]), .A3(n_16), .B1(minus[14]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(L[14]), .ZN(n_17));
   INV_X1 i_20 (.A(minus[14]), .ZN(n_18));
endmodule

module datapath__0_121(R, L, plus);
   input [15:0]R;
   input [15:0]L;
   output [15:0]plus;

   HA_X1 i_1 (.A(R[0]), .B(L[0]), .CO(n_1), .S(plus[0]));
   FA_X1 i_2 (.A(R[1]), .B(L[1]), .CI(n_1), .CO(n_2), .S(plus[1]));
   FA_X1 i_3 (.A(R[2]), .B(L[2]), .CI(n_2), .CO(n_3), .S(plus[2]));
   FA_X1 i_4 (.A(R[3]), .B(L[3]), .CI(n_3), .CO(n_4), .S(plus[3]));
   FA_X1 i_5 (.A(R[4]), .B(L[4]), .CI(n_4), .CO(n_5), .S(plus[4]));
   FA_X1 i_6 (.A(R[5]), .B(L[5]), .CI(n_5), .CO(n_6), .S(plus[5]));
   FA_X1 i_7 (.A(R[6]), .B(L[6]), .CI(n_6), .CO(n_7), .S(plus[6]));
   FA_X1 i_8 (.A(R[7]), .B(L[7]), .CI(n_7), .CO(n_8), .S(plus[7]));
   FA_X1 i_9 (.A(R[8]), .B(L[8]), .CI(n_8), .CO(n_9), .S(plus[8]));
   FA_X1 i_10 (.A(R[9]), .B(L[9]), .CI(n_9), .CO(n_10), .S(plus[9]));
   FA_X1 i_11 (.A(R[10]), .B(L[10]), .CI(n_10), .CO(n_11), .S(plus[10]));
   FA_X1 i_12 (.A(R[11]), .B(L[11]), .CI(n_11), .CO(n_12), .S(plus[11]));
   FA_X1 i_13 (.A(R[12]), .B(L[12]), .CI(n_12), .CO(n_13), .S(plus[12]));
   FA_X1 i_14 (.A(R[13]), .B(L[13]), .CI(n_13), .CO(n_14), .S(plus[13]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(plus[14]));
   OAI22_X1 i_15 (.A1(n_18), .A2(L[14]), .B1(R[14]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(R[15]), .B(n_15), .Z(plus[15]));
   OAI33_X1 i_17 (.A1(n_18), .A2(L[14]), .A3(n_16), .B1(R[14]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(L[14]), .ZN(n_17));
   INV_X1 i_20 (.A(R[14]), .ZN(n_18));
endmodule

module datapath__0_124(minus, L, p_0);
   input [15:0]minus;
   input [15:0]L;
   output [15:0]p_0;

   HA_X1 i_1 (.A(minus[0]), .B(L[0]), .CO(n_1), .S(p_0[0]));
   FA_X1 i_2 (.A(minus[1]), .B(L[1]), .CI(n_1), .CO(n_2), .S(p_0[1]));
   FA_X1 i_3 (.A(minus[2]), .B(L[2]), .CI(n_2), .CO(n_3), .S(p_0[2]));
   FA_X1 i_4 (.A(minus[3]), .B(L[3]), .CI(n_3), .CO(n_4), .S(p_0[3]));
   FA_X1 i_5 (.A(minus[4]), .B(L[4]), .CI(n_4), .CO(n_5), .S(p_0[4]));
   FA_X1 i_6 (.A(minus[5]), .B(L[5]), .CI(n_5), .CO(n_6), .S(p_0[5]));
   FA_X1 i_7 (.A(minus[6]), .B(L[6]), .CI(n_6), .CO(n_7), .S(p_0[6]));
   FA_X1 i_8 (.A(minus[7]), .B(L[7]), .CI(n_7), .CO(n_8), .S(p_0[7]));
   FA_X1 i_9 (.A(minus[8]), .B(L[8]), .CI(n_8), .CO(n_9), .S(p_0[8]));
   FA_X1 i_10 (.A(minus[9]), .B(L[9]), .CI(n_9), .CO(n_10), .S(p_0[9]));
   FA_X1 i_11 (.A(minus[10]), .B(L[10]), .CI(n_10), .CO(n_11), .S(p_0[10]));
   FA_X1 i_12 (.A(minus[11]), .B(L[11]), .CI(n_11), .CO(n_12), .S(p_0[11]));
   FA_X1 i_13 (.A(minus[12]), .B(L[12]), .CI(n_12), .CO(n_13), .S(p_0[12]));
   FA_X1 i_14 (.A(minus[13]), .B(L[13]), .CI(n_13), .CO(n_14), .S(p_0[13]));
   XNOR2_X1 i_0 (.A(n_16), .B(n_0), .ZN(p_0[14]));
   OAI22_X1 i_15 (.A1(n_18), .A2(L[14]), .B1(minus[14]), .B2(n_17), .ZN(n_0));
   XOR2_X1 i_16 (.A(minus[15]), .B(n_15), .Z(p_0[15]));
   OAI33_X1 i_17 (.A1(n_18), .A2(L[14]), .A3(n_16), .B1(minus[14]), .B2(n_17), 
      .B3(n_14), .ZN(n_15));
   INV_X1 i_18 (.A(n_14), .ZN(n_16));
   INV_X1 i_19 (.A(L[14]), .ZN(n_17));
   INV_X1 i_20 (.A(minus[14]), .ZN(n_18));
endmodule

module fpu_multiplier(mode, clk, rst, enbl, in_a, in_b, out_c, done, err, zero, 
      posv);
   input [1:0]mode;
   input clk;
   input rst;
   input enbl;
   input [63:0]in_a;
   input [63:0]in_b;
   output [63:0]out_c;
   output done;
   output err;
   output zero;
   output posv;

   wire n_0_0;
   wire n_0_1;
   wire n_0_2;
   wire n_0_3;
   wire n_0_5;
   wire n_0_6;
   wire n_0_7;
   wire n_0_8;
   wire n_0_9;
   wire n_0_10;
   wire n_0_11;
   wire n_0_12;
   wire n_0_13;
   wire n_0_14;
   wire n_0_15;
   wire n_0_16;
   wire n_0_17;
   wire n_0_18;
   wire n_0_19;
   wire n_0_20;
   wire n_0_21;
   wire n_0_22;
   wire n_0_23;
   wire n_0_24;
   wire n_0_25;
   wire n_0_26;
   wire n_0_27;
   wire n_0_28;
   wire n_0_29;
   wire n_0_30;
   wire n_0_31;
   wire n_0_32;
   wire n_0_33;
   wire n_0_34;
   wire n_0_35;
   wire n_0_36;
   wire n_0_37;
   wire n_0_38;
   wire n_0_39;
   wire n_0_40;
   wire n_0_41;
   wire n_0_42;
   wire n_0_43;
   wire n_0_44;
   wire n_0_45;
   wire n_0_46;
   wire n_0_47;
   wire n_0_48;
   wire n_0_49;
   wire n_0_50;
   wire n_0_51;
   wire n_0_52;
   wire n_0_53;
   wire n_0_54;
   wire n_0_55;
   wire n_0_56;
   wire n_0_57;
   wire n_0_58;
   wire n_0_59;
   wire n_0_60;
   wire n_0_61;
   wire n_0_62;
   wire n_0_63;
   wire n_0_64;
   wire n_0_65;
   wire n_0_66;
   wire n_0_67;
   wire n_0_68;
   wire n_0_69;
   wire n_0_70;
   wire n_0_71;
   wire n_0_72;
   wire n_0_73;
   wire n_0_74;
   wire n_0_75;
   wire n_0_76;
   wire n_0_77;
   wire n_0_78;
   wire n_0_79;
   wire n_0_80;
   wire n_0_81;
   wire n_0_82;
   wire n_0_83;
   wire n_0_84;
   wire n_0_85;
   wire n_0_86;
   wire n_0_87;
   wire n_0_88;
   wire n_0_89;
   wire n_0_90;
   wire n_0_91;
   wire n_0_92;
   wire n_0_93;
   wire n_0_94;
   wire n_0_95;
   wire n_0_96;
   wire n_0_97;
   wire n_0_98;
   wire n_0_99;
   wire n_0_100;
   wire n_0_101;
   wire n_0_102;
   wire n_0_103;
   wire n_0_104;
   wire n_0_105;
   wire n_0_106;
   wire n_0_107;
   wire n_0_108;
   wire n_0_109;
   wire n_0_110;
   wire n_0_111;
   wire n_0_112;
   wire n_0_113;
   wire n_0_114;
   wire n_0_115;
   wire n_0_116;
   wire n_0_117;
   wire n_0_118;
   wire n_0_119;
   wire n_0_120;
   wire n_0_121;
   wire n_0_122;
   wire n_0_123;
   wire n_0_124;
   wire n_0_125;
   wire n_0_126;
   wire n_0_127;
   wire n_0_128;
   wire n_0_129;
   wire n_0_130;
   wire n_0_131;
   wire n_0_132;
   wire n_0_133;
   wire n_0_134;
   wire n_0_135;
   wire n_0_136;
   wire n_0_137;
   wire n_0_138;
   wire n_0_139;
   wire n_0_140;
   wire n_0_141;
   wire n_0_142;
   wire n_0_143;
   wire n_0_144;
   wire n_0_145;
   wire n_0_146;
   wire n_0_147;
   wire n_0_148;
   wire n_0_149;
   wire n_0_150;
   wire n_0_151;
   wire n_0_152;
   wire n_0_153;
   wire n_0_154;
   wire n_0_155;
   wire n_0_156;
   wire n_0_157;
   wire n_0_158;
   wire n_0_159;
   wire n_0_160;
   wire n_0_161;
   wire n_0_162;
   wire n_0_163;
   wire n_0_164;
   wire n_0_165;
   wire n_0_166;
   wire n_0_167;
   wire n_0_168;
   wire n_0_169;
   wire n_0_170;
   wire n_0_171;
   wire n_0_172;
   wire n_0_173;
   wire n_0_174;
   wire n_0_175;
   wire n_0_176;
   wire n_0_177;
   wire n_0_178;
   wire n_0_179;
   wire n_0_180;
   wire n_0_181;
   wire n_0_182;
   wire n_0_183;
   wire n_0_184;
   wire n_0_185;
   wire n_0_186;
   wire n_0_187;
   wire n_0_188;
   wire n_0_189;
   wire n_0_190;
   wire n_0_191;
   wire n_0_192;
   wire n_0_193;
   wire n_0_194;
   wire n_0_195;
   wire n_0_196;
   wire n_0_197;
   wire n_0_198;
   wire n_0_199;
   wire n_0_200;
   wire n_0_201;
   wire n_0_202;
   wire n_0_203;
   wire n_0_204;
   wire n_0_205;
   wire n_0_206;
   wire n_0_207;
   wire n_0_208;
   wire n_0_209;
   wire n_0_210;
   wire n_0_211;
   wire n_0_212;
   wire n_0_213;
   wire n_0_214;
   wire n_0_215;
   wire n_0_216;
   wire n_0_217;
   wire n_0_218;
   wire n_0_219;
   wire n_0_220;
   wire n_0_221;
   wire n_0_222;
   wire n_0_223;
   wire n_0_224;
   wire n_0_225;
   wire n_0_226;
   wire n_0_227;
   wire n_0_228;
   wire n_0_229;
   wire n_0_230;
   wire n_0_231;
   wire n_0_232;
   wire n_0_233;
   wire n_0_234;
   wire n_0_235;
   wire n_0_236;
   wire n_0_237;
   wire n_0_238;
   wire n_0_239;
   wire n_0_240;
   wire n_0_241;
   wire n_0_242;
   wire n_0_243;
   wire n_0_244;
   wire n_0_245;
   wire n_0_246;
   wire n_0_247;
   wire n_0_248;
   wire n_0_249;
   wire n_0_250;
   wire n_0_251;
   wire n_0_252;
   wire n_0_253;
   wire n_0_254;
   wire n_0_255;
   wire n_0_256;
   wire n_0_257;
   wire n_0_258;
   wire n_0_259;
   wire n_0_260;
   wire n_0_261;
   wire n_0_262;
   wire n_0_263;
   wire n_0_264;
   wire n_0_265;
   wire n_0_266;
   wire n_0_267;
   wire n_0_268;
   wire n_0_269;
   wire n_0_270;
   wire n_0_271;
   wire n_0_272;
   wire n_0_273;
   wire n_0_274;
   wire n_0_275;
   wire n_0_276;
   wire n_0_277;
   wire n_0_278;
   wire n_0_279;
   wire n_0_280;
   wire n_0_281;
   wire n_0_282;
   wire n_0_283;
   wire n_0_284;
   wire n_0_285;
   wire n_0_286;
   wire n_0_287;
   wire n_0_288;
   wire error;
   wire n_0_289;
   wire n_0_290;
   wire n_0_4;
   wire n_0_1_168;
   wire n_0_1_3;
   wire n_0_1_169;
   wire n_0_1_4;
   wire n_0_1_170;
   wire n_0_1_5;
   wire n_0_1_171;
   wire n_0_1_6;
   wire n_0_1_172;
   wire n_0_1_7;
   wire n_0_1_173;
   wire n_0_1_8;
   wire n_0_1_174;
   wire n_0_1_9;
   wire n_0_1_175;
   wire n_0_1_10;
   wire n_0_1_176;
   wire n_0_1_11;
   wire n_0_1_177;
   wire n_0_1_12;
   wire n_0_1_178;
   wire n_0_1_13;
   wire n_0_1_179;
   wire n_0_1_14;
   wire n_0_1_180;
   wire n_0_1_15;
   wire n_0_1_181;
   wire n_0_1_0;
   wire n_0_1_182;
   wire n_0_1_1;
   wire n_0_1_183;
   wire n_0_1_2;
   wire n_0_1_184;
   wire n_0_1_16;
   wire n_0_1_185;
   wire n_0_1_17;
   wire n_0_1_186;
   wire n_0_1_18;
   wire n_0_1_187;
   wire n_0_1_19;
   wire n_0_1_188;
   wire n_0_1_20;
   wire n_0_1_189;
   wire n_0_1_21;
   wire n_0_1_190;
   wire n_0_1_22;
   wire n_0_1_191;
   wire n_0_1_23;
   wire n_0_1_192;
   wire n_0_1_24;
   wire n_0_1_193;
   wire n_0_1_25;
   wire n_0_1_194;
   wire n_0_1_26;
   wire n_0_1_195;
   wire n_0_1_27;
   wire n_0_1_196;
   wire n_0_1_28;
   wire n_0_1_197;
   wire n_0_1_29;
   wire n_0_1_198;
   wire n_0_1_30;
   wire n_0_1_199;
   wire n_0_1_31;
   wire n_0_1_200;
   wire n_0_1_32;
   wire n_0_1_201;
   wire n_0_1_33;
   wire n_0_1_202;
   wire n_0_1_34;
   wire n_0_1_203;
   wire n_0_1_35;
   wire n_0_1_204;
   wire n_0_1_36;
   wire n_0_1_205;
   wire n_0_1_37;
   wire n_0_1_206;
   wire n_0_1_38;
   wire n_0_1_207;
   wire n_0_1_39;
   wire n_0_1_208;
   wire n_0_1_40;
   wire n_0_1_209;
   wire n_0_1_41;
   wire n_0_1_210;
   wire n_0_1_42;
   wire n_0_1_211;
   wire n_0_1_43;
   wire n_0_1_212;
   wire n_0_1_44;
   wire n_0_1_213;
   wire n_0_1_45;
   wire n_0_1_214;
   wire n_0_1_46;
   wire n_0_1_215;
   wire n_0_1_47;
   wire n_0_1_216;
   wire n_0_1_48;
   wire n_0_1_217;
   wire n_0_1_49;
   wire n_0_1_218;
   wire n_0_1_50;
   wire n_0_1_219;
   wire n_0_1_51;
   wire n_0_1_220;
   wire n_0_1_52;
   wire n_0_1_221;
   wire n_0_1_53;
   wire n_0_1_222;
   wire n_0_1_54;
   wire n_0_1_223;
   wire n_0_1_55;
   wire n_0_1_224;
   wire n_0_1_56;
   wire n_0_1_225;
   wire n_0_1_57;
   wire n_0_1_226;
   wire n_0_1_58;
   wire n_0_1_227;
   wire n_0_1_59;
   wire n_0_1_228;
   wire n_0_1_60;
   wire n_0_1_229;
   wire n_0_1_61;
   wire n_0_1_230;
   wire n_0_1_62;
   wire n_0_1_231;
   wire n_0_1_63;
   wire n_0_1_232;
   wire n_0_1_64;
   wire n_0_1_233;
   wire n_0_1_65;
   wire n_0_1_234;
   wire n_0_1_66;
   wire n_0_1_235;
   wire n_0_1_67;
   wire n_0_1_236;
   wire n_0_1_68;
   wire n_0_1_237;
   wire n_0_1_69;
   wire n_0_1_238;
   wire n_0_1_70;
   wire n_0_1_239;
   wire n_0_1_71;
   wire n_0_1_240;
   wire n_0_1_72;
   wire n_0_1_241;
   wire n_0_1_73;
   wire n_0_1_242;
   wire n_0_1_74;
   wire n_0_1_243;
   wire n_0_1_75;
   wire n_0_1_244;
   wire n_0_1_76;
   wire n_0_1_245;
   wire n_0_1_77;
   wire n_0_1_246;
   wire n_0_1_78;
   wire n_0_1_247;
   wire n_0_1_79;
   wire n_0_1_248;
   wire n_0_1_80;
   wire n_0_1_249;
   wire n_0_1_81;
   wire n_0_1_250;
   wire n_0_1_82;
   wire n_0_1_251;
   wire n_0_1_83;
   wire n_0_1_252;
   wire n_0_1_84;
   wire n_0_1_253;
   wire n_0_1_85;
   wire n_0_1_254;
   wire n_0_1_86;
   wire n_0_1_255;
   wire n_0_1_87;
   wire n_0_1_256;
   wire n_0_1_88;
   wire n_0_1_257;
   wire n_0_1_89;
   wire n_0_1_258;
   wire n_0_1_90;
   wire n_0_1_259;
   wire n_0_1_91;
   wire n_0_1_260;
   wire n_0_1_92;
   wire n_0_1_261;
   wire n_0_1_93;
   wire n_0_1_262;
   wire n_0_1_94;
   wire n_0_1_263;
   wire n_0_1_95;
   wire n_0_1_264;
   wire n_0_1_96;
   wire n_0_1_265;
   wire n_0_1_97;
   wire n_0_1_266;
   wire n_0_1_98;
   wire n_0_1_267;
   wire n_0_1_99;
   wire n_0_1_268;
   wire n_0_1_100;
   wire n_0_1_269;
   wire n_0_1_101;
   wire n_0_1_270;
   wire n_0_1_102;
   wire n_0_1_271;
   wire n_0_1_103;
   wire n_0_1_272;
   wire n_0_1_104;
   wire n_0_1_273;
   wire n_0_1_105;
   wire n_0_1_274;
   wire n_0_1_106;
   wire n_0_1_275;
   wire n_0_1_107;
   wire n_0_1_276;
   wire n_0_1_108;
   wire n_0_1_277;
   wire n_0_1_109;
   wire n_0_1_278;
   wire n_0_1_110;
   wire n_0_1_279;
   wire n_0_1_111;
   wire n_0_1_280;
   wire n_0_1_112;
   wire n_0_1_281;
   wire n_0_1_113;
   wire n_0_1_282;
   wire n_0_1_114;
   wire n_0_1_283;
   wire n_0_1_115;
   wire n_0_1_284;
   wire n_0_1_116;
   wire n_0_1_285;
   wire n_0_1_117;
   wire n_0_1_286;
   wire n_0_1_118;
   wire n_0_1_287;
   wire n_0_1_119;
   wire n_0_1_288;
   wire n_0_1_120;
   wire n_0_1_289;
   wire n_0_1_121;
   wire n_0_1_290;
   wire n_0_1_122;
   wire n_0_1_291;
   wire n_0_1_123;
   wire n_0_1_292;
   wire n_0_1_124;
   wire n_0_1_293;
   wire n_0_1_125;
   wire n_0_1_294;
   wire n_0_1_126;
   wire n_0_1_295;
   wire n_0_1_127;
   wire n_0_1_296;
   wire n_0_1_128;
   wire n_0_1_297;
   wire n_0_1_129;
   wire n_0_1_298;
   wire n_0_1_130;
   wire n_0_1_299;
   wire n_0_1_131;
   wire n_0_1_300;
   wire n_0_1_132;
   wire n_0_1_301;
   wire n_0_1_133;
   wire n_0_1_302;
   wire n_0_1_134;
   wire n_0_1_303;
   wire n_0_1_135;
   wire n_0_1_304;
   wire n_0_1_136;
   wire n_0_1_305;
   wire n_0_1_137;
   wire n_0_1_306;
   wire n_0_1_138;
   wire n_0_1_307;
   wire n_0_1_139;
   wire n_0_1_308;
   wire n_0_1_140;
   wire n_0_1_309;
   wire n_0_1_141;
   wire n_0_1_310;
   wire n_0_1_142;
   wire n_0_1_311;
   wire n_0_1_143;
   wire n_0_1_312;
   wire n_0_1_144;
   wire n_0_1_313;
   wire n_0_1_145;
   wire n_0_1_314;
   wire n_0_1_146;
   wire n_0_1_315;
   wire n_0_1_147;
   wire n_0_1_316;
   wire n_0_1_148;
   wire n_0_1_317;
   wire n_0_1_149;
   wire n_0_1_318;
   wire n_0_1_150;
   wire n_0_1_319;
   wire n_0_1_151;
   wire n_0_1_320;
   wire n_0_1_152;
   wire n_0_1_321;
   wire n_0_1_153;
   wire n_0_1_322;
   wire n_0_1_154;
   wire n_0_1_323;
   wire n_0_1_155;
   wire n_0_1_156;
   wire n_0_1_157;
   wire n_0_1_158;
   wire n_0_1_159;
   wire n_0_1_160;
   wire n_0_1_161;
   wire n_0_1_162;
   wire n_0_1_163;
   wire n_0_1_164;
   wire n_0_1_165;
   wire n_0_1_166;
   wire n_0_1_167;
   wire n_0_1_324;
   wire n_0_1_325;
   wire n_0_1_326;
   wire n_0_1_327;
   wire n_0_1_328;
   wire n_0_1_329;
   wire n_0_1_330;
   wire n_0_1_331;
   wire n_0_1_332;
   wire n_0_1_333;
   wire n_0_1_334;
   wire n_0_1_335;
   wire n_0_1_336;
   wire n_0_1_337;
   wire n_0_1_338;
   wire n_0_1_339;
   wire n_0_1_340;
   wire n_0_1_341;
   wire n_0_1_342;
   wire n_0_1_343;
   wire n_0_1_344;
   wire n_0_1_345;
   wire n_0_1_346;
   wire n_0_1_347;
   wire n_0_1_348;
   wire n_0_1_349;
   wire n_0_1_350;
   wire n_0_1_351;
   wire n_0_1_352;
   wire n_0_1_353;
   wire n_0_1_354;
   wire n_0_1_355;
   wire n_0_1_356;
   wire n_0_1_357;
   wire n_0_1_358;
   wire n_0_1_359;
   wire n_0_291;
   wire n_0_1_360;
   wire n_0_1_361;
   wire n_0_1_362;
   wire n_0_1_363;
   wire n_0_1_364;
   wire n_0_1_365;
   wire n_0_1_366;
   wire n_0_1_367;
   wire n_0_1_368;
   wire n_0_1_369;
   wire n_0_1_370;
   wire n_0_1_371;
   wire n_0_1_372;
   wire n_0_292;
   wire n_0_293;
   wire n_0_1_373;
   wire n_0_1_374;
   wire n_0_1_375;
   wire n_0_1_376;
   wire n_0_294;
   wire n_0_1_377;
   wire n_0_295;
   wire n_0_1_378;
   wire n_0_296;
   wire n_0_1_379;
   wire n_0_297;
   wire n_0_1_380;
   wire n_0_298;
   wire n_0_1_381;
   wire n_0_299;
   wire n_0_1_382;
   wire n_0_300;
   wire n_0_1_383;
   wire n_0_301;
   wire n_0_1_384;
   wire n_0_302;
   wire n_0_1_385;
   wire n_0_303;
   wire n_0_1_386;
   wire n_0_304;
   wire n_0_1_387;
   wire n_0_305;
   wire n_0_1_388;
   wire n_0_306;
   wire n_0_1_389;
   wire n_0_307;
   wire n_0_1_390;
   wire n_0_308;
   wire n_0_1_391;
   wire n_0_309;
   wire n_0_1_392;
   wire \output ;
   wire n_0_1_393;
   wire n_0_1_394;
   wire n_0_1_395;
   wire n_0_1_396;
   wire n_0_1_397;
   wire n_0_310;
   wire n_0_1_398;
   wire n_0_311;
   wire n_0_1_399;
   wire n_0_312;
   wire n_0_1_400;
   wire n_0_313;
   wire n_0_1_401;
   wire n_0_314;
   wire n_0_1_402;
   wire n_0_315;
   wire n_0_1_403;
   wire n_0_316;
   wire n_0_1_404;
   wire n_0_317;
   wire n_0_1_405;
   wire n_0_318;
   wire n_0_1_406;
   wire n_0_319;
   wire n_0_1_407;
   wire n_0_320;
   wire n_0_1_408;
   wire n_0_321;
   wire n_0_1_409;
   wire n_0_322;
   wire n_0_1_410;
   wire n_0_323;
   wire n_0_1_411;
   wire n_0_324;
   wire n_0_1_412;
   wire n_0_1_413;
   wire n_0_1_414;
   wire n_0_1_415;
   wire n_0_1_416;
   wire n_0_325;
   wire n_0_1_417;
   wire n_0_326;
   wire n_0_1_418;
   wire n_0_327;
   wire n_0_1_419;
   wire n_0_328;
   wire n_0_1_420;
   wire n_0_329;
   wire n_0_1_421;
   wire n_0_330;
   wire n_0_1_422;
   wire n_0_331;
   wire n_0_1_423;
   wire n_0_332;
   wire n_0_1_424;
   wire n_0_333;
   wire n_0_1_425;
   wire n_0_334;
   wire n_0_1_426;
   wire n_0_335;
   wire n_0_1_427;
   wire n_0_336;
   wire n_0_1_428;
   wire n_0_337;
   wire n_0_1_429;
   wire n_0_338;
   wire n_0_1_430;
   wire n_0_339;
   wire n_0_1_431;
   wire n_0_1_432;
   wire n_0_1_433;
   wire n_0_1_434;
   wire n_0_1_435;
   wire n_0_340;
   wire n_0_1_436;
   wire n_0_341;
   wire n_0_1_437;
   wire n_0_342;
   wire n_0_1_438;
   wire n_0_343;
   wire n_0_1_439;
   wire n_0_344;
   wire n_0_1_440;
   wire n_0_345;
   wire n_0_1_441;
   wire n_0_346;
   wire n_0_1_442;
   wire n_0_347;
   wire n_0_1_443;
   wire n_0_348;
   wire n_0_1_444;
   wire n_0_349;
   wire n_0_1_445;
   wire n_0_350;
   wire n_0_1_446;
   wire n_0_351;
   wire n_0_1_447;
   wire n_0_352;
   wire n_0_1_448;
   wire n_0_353;
   wire n_0_1_449;
   wire n_0_354;
   wire n_0_1_450;
   wire n_0_1_451;
   wire n_0_1_452;
   wire n_0_1_453;
   wire n_0_1_454;
   wire n_0_355;
   wire n_0_1_455;
   wire n_0_356;
   wire n_0_1_456;
   wire n_0_357;
   wire n_0_1_457;
   wire n_0_358;
   wire n_0_1_458;
   wire n_0_359;
   wire n_0_1_459;
   wire n_0_360;
   wire n_0_1_460;
   wire n_0_361;
   wire n_0_1_461;
   wire n_0_362;
   wire n_0_1_462;
   wire n_0_363;
   wire n_0_1_463;
   wire n_0_364;
   wire n_0_1_464;
   wire n_0_365;
   wire n_0_1_465;
   wire n_0_366;
   wire n_0_1_466;
   wire n_0_367;
   wire n_0_1_467;
   wire n_0_368;
   wire n_0_1_468;
   wire n_0_369;
   wire n_0_1_469;
   wire n_0_1_470;
   wire n_0_1_471;
   wire n_0_1_472;
   wire n_0_1_473;
   wire n_0_370;
   wire n_0_1_474;
   wire n_0_371;
   wire n_0_1_475;
   wire n_0_372;
   wire n_0_1_476;
   wire n_0_373;
   wire n_0_1_477;
   wire n_0_374;
   wire n_0_1_478;
   wire n_0_375;
   wire n_0_1_479;
   wire n_0_376;
   wire n_0_1_480;
   wire n_0_377;
   wire n_0_1_481;
   wire n_0_378;
   wire n_0_1_482;
   wire n_0_379;
   wire n_0_1_483;
   wire n_0_380;
   wire n_0_1_484;
   wire n_0_381;
   wire n_0_1_485;
   wire n_0_382;
   wire n_0_1_486;
   wire n_0_383;
   wire n_0_1_487;
   wire n_0_384;
   wire n_0_1_488;
   wire n_0_1_489;
   wire n_0_1_490;
   wire n_0_1_491;
   wire n_0_1_492;
   wire n_0_385;
   wire n_0_1_493;
   wire n_0_386;
   wire n_0_1_494;
   wire n_0_387;
   wire n_0_1_495;
   wire n_0_388;
   wire n_0_1_496;
   wire n_0_389;
   wire n_0_1_497;
   wire n_0_390;
   wire n_0_1_498;
   wire n_0_391;
   wire n_0_1_499;
   wire n_0_392;
   wire n_0_1_500;
   wire n_0_393;
   wire n_0_1_501;
   wire n_0_394;
   wire n_0_1_502;
   wire n_0_395;
   wire n_0_1_503;
   wire n_0_396;
   wire n_0_1_504;
   wire n_0_397;
   wire n_0_1_505;
   wire n_0_398;
   wire n_0_1_506;
   wire n_0_399;
   wire n_0_1_507;
   wire n_0_1_508;
   wire n_0_1_509;
   wire n_0_1_510;
   wire n_0_1_511;
   wire n_0_400;
   wire n_0_1_512;
   wire n_0_401;
   wire n_0_1_513;
   wire n_0_402;
   wire n_0_1_514;
   wire n_0_403;
   wire n_0_1_515;
   wire n_0_404;
   wire n_0_1_516;
   wire n_0_405;
   wire n_0_1_517;
   wire n_0_406;
   wire n_0_1_518;
   wire n_0_407;
   wire n_0_1_519;
   wire n_0_408;
   wire n_0_1_520;
   wire n_0_409;
   wire n_0_1_521;
   wire n_0_410;
   wire n_0_1_522;
   wire n_0_411;
   wire n_0_1_523;
   wire n_0_412;
   wire n_0_1_524;
   wire n_0_413;
   wire n_0_1_525;
   wire n_0_414;
   wire n_0_1_526;
   wire n_0_1_527;
   wire n_0_1_528;
   wire n_0_1_529;
   wire n_0_1_530;
   wire n_0_415;
   wire n_0_1_531;
   wire n_0_416;
   wire n_0_1_532;
   wire n_0_417;
   wire n_0_1_533;
   wire n_0_418;
   wire n_0_1_534;
   wire n_0_419;
   wire n_0_1_535;
   wire n_0_420;
   wire n_0_1_536;
   wire n_0_421;
   wire n_0_1_537;
   wire n_0_422;
   wire n_0_1_538;
   wire n_0_423;
   wire n_0_1_539;
   wire n_0_424;
   wire n_0_1_540;
   wire n_0_425;
   wire n_0_1_541;
   wire n_0_426;
   wire n_0_1_542;
   wire n_0_427;
   wire n_0_1_543;
   wire n_0_428;
   wire n_0_1_544;
   wire n_0_429;
   wire n_0_1_545;
   wire n_0_1_546;
   wire n_0_1_547;
   wire n_0_1_548;
   wire n_0_1_549;
   wire n_0_430;
   wire n_0_1_550;
   wire n_0_1_551;
   wire n_0_1_552;
   wire n_0_1_553;
   wire n_0_1_554;
   wire n_0_1_555;
   wire n_0_1_556;
   wire n_0_1_557;
   wire n_0_1_558;
   wire n_0_1_559;
   wire n_0_1_560;
   wire n_0_1_561;
   wire n_0_431;
   wire n_0_1_562;
   wire n_0_1_563;
   wire n_0_1_564;
   wire n_0_1_565;
   wire n_0_1_566;
   wire n_0_1_567;
   wire n_0_1_568;
   wire n_0_1_569;
   wire n_0_1_570;
   wire n_0_1_571;
   wire n_0_1_572;
   wire n_0_1_573;
   wire n_0_432;
   wire n_0_1_574;
   wire n_0_1_575;
   wire n_0_1_576;
   wire n_0_1_577;
   wire n_0_1_578;
   wire n_0_1_579;
   wire n_0_1_580;
   wire n_0_1_581;
   wire n_0_1_582;
   wire n_0_1_583;
   wire n_0_1_584;
   wire n_0_1_585;
   wire n_0_433;
   wire n_0_1_586;
   wire n_0_1_587;
   wire n_0_1_588;
   wire n_0_1_589;
   wire n_0_1_590;
   wire n_0_1_591;
   wire n_0_1_592;
   wire n_0_1_593;
   wire n_0_1_594;
   wire n_0_1_595;
   wire n_0_1_596;
   wire n_0_1_597;
   wire n_0_434;
   wire n_0_1_598;
   wire n_0_1_599;
   wire n_0_1_600;
   wire n_0_1_601;
   wire n_0_1_602;
   wire n_0_1_603;
   wire n_0_1_604;
   wire n_0_1_605;
   wire n_0_1_606;
   wire n_0_1_607;
   wire n_0_1_608;
   wire n_0_1_609;
   wire n_0_435;
   wire n_0_1_610;
   wire n_0_1_611;
   wire n_0_1_612;
   wire n_0_1_613;
   wire n_0_1_614;
   wire n_0_1_615;
   wire n_0_1_616;
   wire n_0_1_617;
   wire n_0_1_618;
   wire n_0_1_619;
   wire n_0_1_620;
   wire n_0_1_621;
   wire n_0_436;
   wire n_0_1_622;
   wire n_0_1_623;
   wire n_0_1_624;
   wire n_0_1_625;
   wire n_0_1_626;
   wire n_0_1_627;
   wire n_0_1_628;
   wire n_0_1_629;
   wire n_0_1_630;
   wire n_0_1_631;
   wire n_0_1_632;
   wire n_0_1_633;
   wire n_0_437;
   wire n_0_1_634;
   wire n_0_1_635;
   wire n_0_1_636;
   wire n_0_1_637;
   wire n_0_1_638;
   wire n_0_1_639;
   wire n_0_1_640;
   wire n_0_1_641;
   wire n_0_1_642;
   wire n_0_1_643;
   wire n_0_1_644;
   wire n_0_438;
   wire n_0_1_645;
   wire n_0_1_646;
   wire n_0_1_647;
   wire n_0_1_648;
   wire n_0_1_649;
   wire n_0_1_650;
   wire n_0_1_651;
   wire n_0_1_652;
   wire n_0_1_653;
   wire n_0_1_654;
   wire n_0_1_655;
   wire n_0_1_656;
   wire n_0_1_657;
   wire n_0_1_658;
   wire n_0_1_659;
   wire n_0_1_660;
   wire n_0_439;
   wire n_0_1_661;
   wire n_0_1_662;
   wire n_0_1_663;
   wire n_0_1_664;
   wire n_0_1_665;
   wire n_0_1_666;
   wire n_0_1_667;
   wire n_0_1_668;
   wire n_0_1_669;
   wire n_0_1_670;
   wire n_0_1_671;
   wire n_0_1_672;
   wire n_0_1_673;
   wire n_0_440;
   wire n_0_1_674;
   wire n_0_1_675;
   wire n_0_1_676;
   wire n_0_1_677;
   wire n_0_1_678;
   wire n_0_1_679;
   wire n_0_1_680;
   wire n_0_1_681;
   wire n_0_1_682;
   wire n_0_441;
   wire n_0_1_683;
   wire n_0_1_684;
   wire n_0_1_685;
   wire n_0_1_686;
   wire n_0_1_687;
   wire n_0_1_688;
   wire n_0_1_689;
   wire n_0_442;
   wire n_0_1_690;
   wire n_0_1_691;
   wire n_0_1_692;
   wire n_0_1_693;
   wire n_0_1_694;
   wire n_0_1_695;
   wire n_0_1_696;
   wire n_0_443;
   wire n_0_1_697;
   wire n_0_1_698;
   wire n_0_1_699;
   wire n_0_444;
   wire n_0_1_700;
   wire n_0_1_701;
   wire n_0_1_702;
   wire n_0_1_703;
   wire n_0_1_704;
   wire n_0_1_705;
   wire n_0_1_706;
   wire n_0_1_707;
   wire n_0_1_708;
   wire n_0_1_709;
   wire n_0_1_710;
   wire n_0_1_711;
   wire n_0_1_712;
   wire n_0_1_713;
   wire n_0_1_714;
   wire n_0_1_715;
   wire n_0_1_716;
   wire n_0_1_717;
   wire n_0_1_718;
   wire n_0_1_719;
   wire n_0_1_720;
   wire n_0_1_721;
   wire n_0_1_722;
   wire n_0_1_723;
   wire n_0_1_724;
   wire n_0_1_725;
   wire n_0_1_726;
   wire n_0_1_727;
   wire n_0_1_728;
   wire n_0_1_729;
   wire n_0_1_730;
   wire n_0_1_731;
   wire n_0_1_732;
   wire n_0_1_733;
   wire n_0_1_734;
   wire n_0_1_735;
   wire n_0_1_736;
   wire n_0_1_737;
   wire n_0_1_738;
   wire n_0_1_739;
   wire n_0_1_740;
   wire n_0_1_741;
   wire n_0_1_742;
   wire n_0_1_743;
   wire n_0_1_744;
   wire n_0_1_745;
   wire n_0_1_746;
   wire n_0_1_747;
   wire n_0_1_748;
   wire n_0_1_749;
   wire n_0_1_750;
   wire n_0_1_751;
   wire n_0_1_752;
   wire n_0_1_753;
   wire n_0_1_754;
   wire n_0_1_755;
   wire n_0_1_756;
   wire n_0_1_757;
   wire n_0_1_758;
   wire n_0_1_759;
   wire n_0_1_760;
   wire n_0_1_761;
   wire n_0_1_762;
   wire n_0_1_763;
   wire n_0_1_764;
   wire n_0_1_765;
   wire n_0_1_766;
   wire n_0_1_767;
   wire n_0_1_768;
   wire n_0_1_769;
   wire n_0_1_770;
   wire n_0_1_771;
   wire n_0_1_772;
   wire n_0_1_773;
   wire n_0_445;
   wire n_0_446;
   wire n_0_447;
   wire n_0_448;
   wire n_0_449;
   wire n_0_450;
   wire n_0_451;
   wire n_0_452;
   wire n_0_453;
   wire n_0_454;
   wire n_0_455;
   wire n_0_456;
   wire n_0_457;
   wire n_0_458;
   wire n_0_1_774;
   wire n_0_1_775;
   wire n_0_459;
   wire n_0_1_776;
   wire n_0_1_777;
   wire n_0_1_778;
   wire n_0_1_779;
   wire n_0_1_780;
   wire n_0_1_781;
   wire n_0_1_782;
   wire n_0_1_783;
   wire n_0_1_784;
   wire n_0_1_785;
   wire n_0_1_786;
   wire n_0_1_787;
   wire n_0_1_788;
   wire n_0_1_789;
   wire n_0_1_790;
   wire n_0_1_791;
   wire n_0_1_792;
   wire n_0_1_793;
   wire n_0_1_794;
   wire n_0_1_795;
   wire n_0_1_796;
   wire n_0_1_797;
   wire n_0_1_798;
   wire n_0_1_799;
   wire n_0_1_800;
   wire n_0_1_801;
   wire n_0_1_802;
   wire n_0_1_803;
   wire n_0_1_804;
   wire n_0_1_805;
   wire n_0_1_806;
   wire n_0_1_807;
   wire n_0_1_808;
   wire n_0_1_809;
   wire n_0_1_810;
   wire n_0_1_811;
   wire n_0_1_812;
   wire n_0_1_813;
   wire n_0_1_814;
   wire n_0_1_815;
   wire n_0_1_816;
   wire n_0_1_817;
   wire n_0_1_818;
   wire n_0_1_819;
   wire n_0_1_820;
   wire n_0_1_821;
   wire n_0_1_822;
   wire n_0_1_823;
   wire n_0_1_824;
   wire n_0_1_825;
   wire n_0_1_826;
   wire n_0_1_827;
   wire n_0_460;
   wire n_0_463;
   wire n_0_462;
   wire n_0_465;
   wire n_0_461;
   wire n_0_2_0;
   wire n_0_464;

   assign out_c[63] = out_c[16];
   assign out_c[62] = out_c[16];
   assign out_c[61] = out_c[16];
   assign out_c[60] = out_c[16];
   assign out_c[59] = out_c[16];
   assign out_c[58] = out_c[16];
   assign out_c[57] = out_c[16];
   assign out_c[56] = out_c[16];
   assign out_c[55] = out_c[16];
   assign out_c[54] = out_c[16];
   assign out_c[53] = out_c[16];
   assign out_c[52] = out_c[16];
   assign out_c[51] = out_c[16];
   assign out_c[50] = out_c[16];
   assign out_c[49] = out_c[16];
   assign out_c[48] = out_c[16];
   assign out_c[47] = out_c[16];
   assign out_c[46] = out_c[16];
   assign out_c[45] = out_c[16];
   assign out_c[44] = out_c[16];
   assign out_c[43] = out_c[16];
   assign out_c[42] = out_c[16];
   assign out_c[41] = out_c[16];
   assign out_c[40] = out_c[16];
   assign out_c[39] = out_c[16];
   assign out_c[38] = out_c[16];
   assign out_c[37] = out_c[16];
   assign out_c[36] = out_c[16];
   assign out_c[35] = out_c[16];
   assign out_c[34] = out_c[16];
   assign out_c[33] = out_c[16];
   assign out_c[32] = out_c[16];
   assign out_c[31] = out_c[16];
   assign out_c[30] = out_c[16];
   assign out_c[29] = out_c[16];
   assign out_c[28] = out_c[16];
   assign out_c[27] = out_c[16];
   assign out_c[26] = out_c[16];
   assign out_c[25] = out_c[16];
   assign out_c[24] = out_c[16];
   assign out_c[23] = out_c[16];
   assign out_c[22] = out_c[16];
   assign out_c[21] = out_c[16];
   assign out_c[20] = out_c[16];
   assign out_c[19] = out_c[16];
   assign out_c[18] = out_c[16];
   assign out_c[17] = out_c[16];

   DFFR_X1 posv_reg (.D(n_0_292), .RN(n_0_462), .CK(n_0_4), .Q(posv), .QN());
   datapath__0_57 i_0_31 (.R({in_a[15], in_a[14], in_a[13], in_a[12], in_a[11], 
      in_a[10], in_a[9], in_a[8], in_a[7], in_a[6], in_a[5], in_a[4], in_a[3], 
      in_a[2], in_a[1], in_a[0]}), .L({uc_0, n_0_444, n_0_443, n_0_442, n_0_441, 
      n_0_440, n_0_439, n_0_438, n_0_437, n_0_436, n_0_435, n_0_434, n_0_433, 
      n_0_432, n_0_431, n_0_430}), .plus({n_0_16, n_0_15, n_0_14, n_0_13, n_0_12, 
      n_0_11, n_0_10, n_0_9, n_0_8, n_0_7, n_0_6, n_0_5, n_0_3, n_0_2, n_0_1, 
      n_0_0}));
   datapath__0_60 i_0_32 (.minus({n_0_459, n_0_458, n_0_457, n_0_456, n_0_455, 
      n_0_454, n_0_453, n_0_452, n_0_451, n_0_450, n_0_449, n_0_448, n_0_447, 
      n_0_446, n_0_445, in_a[0]}), .L({uc_1, n_0_444, n_0_443, n_0_442, n_0_441, 
      n_0_440, n_0_439, n_0_438, n_0_437, n_0_436, n_0_435, n_0_434, n_0_433, 
      n_0_432, n_0_431, n_0_430}), .p_0({n_0_32, n_0_31, n_0_30, n_0_29, n_0_28, 
      n_0_27, n_0_26, n_0_25, n_0_24, n_0_23, n_0_22, n_0_21, n_0_20, n_0_19, 
      n_0_18, n_0_17}));
   datapath__0_65 i_0_35 (.R({in_a[15], in_a[14], in_a[13], in_a[12], in_a[11], 
      in_a[10], in_a[9], in_a[8], in_a[7], in_a[6], in_a[5], in_a[4], in_a[3], 
      in_a[2], in_a[1], in_a[0]}), .L({uc_2, n_0_429, n_0_428, n_0_427, n_0_426, 
      n_0_425, n_0_424, n_0_423, n_0_422, n_0_421, n_0_420, n_0_419, n_0_418, 
      n_0_417, n_0_416, n_0_415}), .plus({n_0_48, n_0_47, n_0_46, n_0_45, n_0_44, 
      n_0_43, n_0_42, n_0_41, n_0_40, n_0_39, n_0_38, n_0_37, n_0_36, n_0_35, 
      n_0_34, n_0_33}));
   datapath__0_68 i_0_36 (.minus({n_0_459, n_0_458, n_0_457, n_0_456, n_0_455, 
      n_0_454, n_0_453, n_0_452, n_0_451, n_0_450, n_0_449, n_0_448, n_0_447, 
      n_0_446, n_0_445, in_a[0]}), .L({uc_3, n_0_429, n_0_428, n_0_427, n_0_426, 
      n_0_425, n_0_424, n_0_423, n_0_422, n_0_421, n_0_420, n_0_419, n_0_418, 
      n_0_417, n_0_416, n_0_415}), .p_0({n_0_64, n_0_63, n_0_62, n_0_61, n_0_60, 
      n_0_59, n_0_58, n_0_57, n_0_56, n_0_55, n_0_54, n_0_53, n_0_52, n_0_51, 
      n_0_50, n_0_49}));
   datapath__0_73 i_0_39 (.R({in_a[15], in_a[14], in_a[13], in_a[12], in_a[11], 
      in_a[10], in_a[9], in_a[8], in_a[7], in_a[6], in_a[5], in_a[4], in_a[3], 
      in_a[2], in_a[1], in_a[0]}), .L({uc_4, n_0_414, n_0_413, n_0_412, n_0_411, 
      n_0_410, n_0_409, n_0_408, n_0_407, n_0_406, n_0_405, n_0_404, n_0_403, 
      n_0_402, n_0_401, n_0_400}), .plus({n_0_80, n_0_79, n_0_78, n_0_77, n_0_76, 
      n_0_75, n_0_74, n_0_73, n_0_72, n_0_71, n_0_70, n_0_69, n_0_68, n_0_67, 
      n_0_66, n_0_65}));
   datapath__0_76 i_0_40 (.minus({n_0_459, n_0_458, n_0_457, n_0_456, n_0_455, 
      n_0_454, n_0_453, n_0_452, n_0_451, n_0_450, n_0_449, n_0_448, n_0_447, 
      n_0_446, n_0_445, in_a[0]}), .L({uc_5, n_0_414, n_0_413, n_0_412, n_0_411, 
      n_0_410, n_0_409, n_0_408, n_0_407, n_0_406, n_0_405, n_0_404, n_0_403, 
      n_0_402, n_0_401, n_0_400}), .p_0({n_0_96, n_0_95, n_0_94, n_0_93, n_0_92, 
      n_0_91, n_0_90, n_0_89, n_0_88, n_0_87, n_0_86, n_0_85, n_0_84, n_0_83, 
      n_0_82, n_0_81}));
   datapath__0_81 i_0_43 (.R({in_a[15], in_a[14], in_a[13], in_a[12], in_a[11], 
      in_a[10], in_a[9], in_a[8], in_a[7], in_a[6], in_a[5], in_a[4], in_a[3], 
      in_a[2], in_a[1], in_a[0]}), .L({uc_6, n_0_399, n_0_398, n_0_397, n_0_396, 
      n_0_395, n_0_394, n_0_393, n_0_392, n_0_391, n_0_390, n_0_389, n_0_388, 
      n_0_387, n_0_386, n_0_385}), .plus({n_0_112, n_0_111, n_0_110, n_0_109, 
      n_0_108, n_0_107, n_0_106, n_0_105, n_0_104, n_0_103, n_0_102, n_0_101, 
      n_0_100, n_0_99, n_0_98, n_0_97}));
   datapath__0_84 i_0_44 (.minus({n_0_459, n_0_458, n_0_457, n_0_456, n_0_455, 
      n_0_454, n_0_453, n_0_452, n_0_451, n_0_450, n_0_449, n_0_448, n_0_447, 
      n_0_446, n_0_445, in_a[0]}), .L({uc_7, n_0_399, n_0_398, n_0_397, n_0_396, 
      n_0_395, n_0_394, n_0_393, n_0_392, n_0_391, n_0_390, n_0_389, n_0_388, 
      n_0_387, n_0_386, n_0_385}), .p_0({n_0_128, n_0_127, n_0_126, n_0_125, 
      n_0_124, n_0_123, n_0_122, n_0_121, n_0_120, n_0_119, n_0_118, n_0_117, 
      n_0_116, n_0_115, n_0_114, n_0_113}));
   datapath__0_89 i_0_47 (.R({in_a[15], in_a[14], in_a[13], in_a[12], in_a[11], 
      in_a[10], in_a[9], in_a[8], in_a[7], in_a[6], in_a[5], in_a[4], in_a[3], 
      in_a[2], in_a[1], in_a[0]}), .L({uc_8, n_0_384, n_0_383, n_0_382, n_0_381, 
      n_0_380, n_0_379, n_0_378, n_0_377, n_0_376, n_0_375, n_0_374, n_0_373, 
      n_0_372, n_0_371, n_0_370}), .plus({n_0_144, n_0_143, n_0_142, n_0_141, 
      n_0_140, n_0_139, n_0_138, n_0_137, n_0_136, n_0_135, n_0_134, n_0_133, 
      n_0_132, n_0_131, n_0_130, n_0_129}));
   datapath__0_92 i_0_48 (.minus({n_0_459, n_0_458, n_0_457, n_0_456, n_0_455, 
      n_0_454, n_0_453, n_0_452, n_0_451, n_0_450, n_0_449, n_0_448, n_0_447, 
      n_0_446, n_0_445, in_a[0]}), .L({uc_9, n_0_384, n_0_383, n_0_382, n_0_381, 
      n_0_380, n_0_379, n_0_378, n_0_377, n_0_376, n_0_375, n_0_374, n_0_373, 
      n_0_372, n_0_371, n_0_370}), .p_0({n_0_160, n_0_159, n_0_158, n_0_157, 
      n_0_156, n_0_155, n_0_154, n_0_153, n_0_152, n_0_151, n_0_150, n_0_149, 
      n_0_148, n_0_147, n_0_146, n_0_145}));
   datapath__0_97 i_0_51 (.R({in_a[15], in_a[14], in_a[13], in_a[12], in_a[11], 
      in_a[10], in_a[9], in_a[8], in_a[7], in_a[6], in_a[5], in_a[4], in_a[3], 
      in_a[2], in_a[1], in_a[0]}), .L({uc_10, n_0_369, n_0_368, n_0_367, n_0_366, 
      n_0_365, n_0_364, n_0_363, n_0_362, n_0_361, n_0_360, n_0_359, n_0_358, 
      n_0_357, n_0_356, n_0_355}), .plus({n_0_176, n_0_175, n_0_174, n_0_173, 
      n_0_172, n_0_171, n_0_170, n_0_169, n_0_168, n_0_167, n_0_166, n_0_165, 
      n_0_164, n_0_163, n_0_162, n_0_161}));
   datapath__0_100 i_0_52 (.minus({n_0_459, n_0_458, n_0_457, n_0_456, n_0_455, 
      n_0_454, n_0_453, n_0_452, n_0_451, n_0_450, n_0_449, n_0_448, n_0_447, 
      n_0_446, n_0_445, in_a[0]}), .L({uc_11, n_0_369, n_0_368, n_0_367, n_0_366, 
      n_0_365, n_0_364, n_0_363, n_0_362, n_0_361, n_0_360, n_0_359, n_0_358, 
      n_0_357, n_0_356, n_0_355}), .p_0({n_0_192, n_0_191, n_0_190, n_0_189, 
      n_0_188, n_0_187, n_0_186, n_0_185, n_0_184, n_0_183, n_0_182, n_0_181, 
      n_0_180, n_0_179, n_0_178, n_0_177}));
   datapath__0_105 i_0_55 (.R({in_a[15], in_a[14], in_a[13], in_a[12], in_a[11], 
      in_a[10], in_a[9], in_a[8], in_a[7], in_a[6], in_a[5], in_a[4], in_a[3], 
      in_a[2], in_a[1], in_a[0]}), .L({uc_12, n_0_354, n_0_353, n_0_352, n_0_351, 
      n_0_350, n_0_349, n_0_348, n_0_347, n_0_346, n_0_345, n_0_344, n_0_343, 
      n_0_342, n_0_341, n_0_340}), .plus({n_0_208, n_0_207, n_0_206, n_0_205, 
      n_0_204, n_0_203, n_0_202, n_0_201, n_0_200, n_0_199, n_0_198, n_0_197, 
      n_0_196, n_0_195, n_0_194, n_0_193}));
   datapath__0_108 i_0_56 (.minus({n_0_459, n_0_458, n_0_457, n_0_456, n_0_455, 
      n_0_454, n_0_453, n_0_452, n_0_451, n_0_450, n_0_449, n_0_448, n_0_447, 
      n_0_446, n_0_445, in_a[0]}), .L({uc_13, n_0_354, n_0_353, n_0_352, n_0_351, 
      n_0_350, n_0_349, n_0_348, n_0_347, n_0_346, n_0_345, n_0_344, n_0_343, 
      n_0_342, n_0_341, n_0_340}), .p_0({n_0_224, n_0_223, n_0_222, n_0_221, 
      n_0_220, n_0_219, n_0_218, n_0_217, n_0_216, n_0_215, n_0_214, n_0_213, 
      n_0_212, n_0_211, n_0_210, n_0_209}));
   datapath__0_113 i_0_59 (.R({in_a[15], in_a[14], in_a[13], in_a[12], in_a[11], 
      in_a[10], in_a[9], in_a[8], in_a[7], in_a[6], in_a[5], in_a[4], in_a[3], 
      in_a[2], in_a[1], in_a[0]}), .L({uc_14, n_0_339, n_0_338, n_0_337, n_0_336, 
      n_0_335, n_0_334, n_0_333, n_0_332, n_0_331, n_0_330, n_0_329, n_0_328, 
      n_0_327, n_0_326, n_0_325}), .plus({n_0_240, n_0_239, n_0_238, n_0_237, 
      n_0_236, n_0_235, n_0_234, n_0_233, n_0_232, n_0_231, n_0_230, n_0_229, 
      n_0_228, n_0_227, n_0_226, n_0_225}));
   datapath__0_116 i_0_60 (.minus({n_0_459, n_0_458, n_0_457, n_0_456, n_0_455, 
      n_0_454, n_0_453, n_0_452, n_0_451, n_0_450, n_0_449, n_0_448, n_0_447, 
      n_0_446, n_0_445, in_a[0]}), .L({uc_15, n_0_339, n_0_338, n_0_337, n_0_336, 
      n_0_335, n_0_334, n_0_333, n_0_332, n_0_331, n_0_330, n_0_329, n_0_328, 
      n_0_327, n_0_326, n_0_325}), .p_0({n_0_256, n_0_255, n_0_254, n_0_253, 
      n_0_252, n_0_251, n_0_250, n_0_249, n_0_248, n_0_247, n_0_246, n_0_245, 
      n_0_244, n_0_243, n_0_242, n_0_241}));
   datapath__0_121 i_0_63 (.R({in_a[15], in_a[14], in_a[13], in_a[12], in_a[11], 
      in_a[10], in_a[9], in_a[8], in_a[7], in_a[6], in_a[5], in_a[4], in_a[3], 
      in_a[2], in_a[1], in_a[0]}), .L({uc_16, n_0_324, n_0_323, n_0_322, n_0_321, 
      n_0_320, n_0_319, n_0_318, n_0_317, n_0_316, n_0_315, n_0_314, n_0_313, 
      n_0_312, n_0_311, n_0_310}), .plus({n_0_272, n_0_271, n_0_270, n_0_269, 
      n_0_268, n_0_267, n_0_266, n_0_265, n_0_264, n_0_263, n_0_262, n_0_261, 
      n_0_260, n_0_259, n_0_258, n_0_257}));
   datapath__0_124 i_0_64 (.minus({n_0_459, n_0_458, n_0_457, n_0_456, n_0_455, 
      n_0_454, n_0_453, n_0_452, n_0_451, n_0_450, n_0_449, n_0_448, n_0_447, 
      n_0_446, n_0_445, in_a[0]}), .L({uc_17, n_0_324, n_0_323, n_0_322, n_0_321, 
      n_0_320, n_0_319, n_0_318, n_0_317, n_0_316, n_0_315, n_0_314, n_0_313, 
      n_0_312, n_0_311, n_0_310}), .p_0({n_0_288, n_0_287, n_0_286, n_0_285, 
      n_0_284, n_0_283, n_0_282, n_0_281, n_0_280, n_0_279, n_0_278, n_0_277, 
      n_0_276, n_0_275, n_0_274, n_0_273}));
   DFFR_X1 zero_reg (.D(n_0_293), .RN(n_0_462), .CK(n_0_4), .Q(zero), .QN());
   DFFRS_X1 err_reg (.D(n_0_291), .RN(n_0_463), .SN(n_0_465), .CK(n_0_4), 
      .Q(err), .QN());
   DFFRS_X1 done_reg (.D(1'b1), .RN(n_0_461), .SN(n_0_290), .CK(n_0_4), .Q(done), 
      .QN());
   DFFR_X1 \out_c_reg[63]  (.D(\output ), .RN(n_0_462), .CK(n_0_4), .Q(out_c[16]), 
      .QN());
   DFFR_X1 \out_c_reg[15]  (.D(n_0_309), .RN(n_0_462), .CK(n_0_4), .Q(out_c[15]), 
      .QN());
   DFFR_X1 \out_c_reg[14]  (.D(n_0_308), .RN(n_0_462), .CK(n_0_4), .Q(out_c[14]), 
      .QN());
   DFFR_X1 \out_c_reg[13]  (.D(n_0_307), .RN(n_0_462), .CK(n_0_4), .Q(out_c[13]), 
      .QN());
   DFFR_X1 \out_c_reg[12]  (.D(n_0_306), .RN(n_0_462), .CK(n_0_4), .Q(out_c[12]), 
      .QN());
   DFFR_X1 \out_c_reg[11]  (.D(n_0_305), .RN(n_0_462), .CK(n_0_4), .Q(out_c[11]), 
      .QN());
   DFFR_X1 \out_c_reg[10]  (.D(n_0_304), .RN(n_0_462), .CK(n_0_4), .Q(out_c[10]), 
      .QN());
   DFFR_X1 \out_c_reg[9]  (.D(n_0_303), .RN(n_0_462), .CK(n_0_4), .Q(out_c[9]), 
      .QN());
   DFFR_X1 \out_c_reg[8]  (.D(n_0_302), .RN(n_0_462), .CK(n_0_4), .Q(out_c[8]), 
      .QN());
   DFFR_X1 \out_c_reg[7]  (.D(n_0_301), .RN(n_0_462), .CK(n_0_4), .Q(out_c[7]), 
      .QN());
   DFFR_X1 \out_c_reg[6]  (.D(n_0_300), .RN(n_0_462), .CK(n_0_4), .Q(out_c[6]), 
      .QN());
   DFFR_X1 \out_c_reg[5]  (.D(n_0_299), .RN(n_0_462), .CK(n_0_4), .Q(out_c[5]), 
      .QN());
   DFFR_X1 \out_c_reg[4]  (.D(n_0_298), .RN(n_0_462), .CK(n_0_4), .Q(out_c[4]), 
      .QN());
   DFFR_X1 \out_c_reg[3]  (.D(n_0_297), .RN(n_0_462), .CK(n_0_4), .Q(out_c[3]), 
      .QN());
   DFFR_X1 \out_c_reg[2]  (.D(n_0_296), .RN(n_0_462), .CK(n_0_4), .Q(out_c[2]), 
      .QN());
   DFFR_X1 \out_c_reg[1]  (.D(n_0_295), .RN(n_0_462), .CK(n_0_4), .Q(out_c[1]), 
      .QN());
   DFFR_X1 \out_c_reg[0]  (.D(n_0_294), .RN(n_0_462), .CK(n_0_4), .Q(out_c[0]), 
      .QN());
   DFFR_X1 error_reg (.D(n_0_289), .RN(n_0_290), .CK(clk), .Q(error), .QN());
   MUX2_X1 error_reg_enable_mux_0 (.A(error), .B(n_0_291), .S(n_0_460), .Z(
      n_0_289));
   INV_X1 i_0_0_0 (.A(rst), .ZN(n_0_290));
   CLKGATETST_X1 clk_gate_posv_reg (.CK(clk), .E(n_0_464), .SE(1'b0), .GCK(n_0_4));
   FA_X1 i_0_1_0 (.A(in_a[1]), .B(n_0_1_358), .CI(n_0_1_157), .CO(n_0_1_3), 
      .S(n_0_1_168));
   FA_X1 i_0_1_1 (.A(in_a[2]), .B(n_0_1_357), .CI(n_0_1_3), .CO(n_0_1_4), 
      .S(n_0_1_169));
   FA_X1 i_0_1_2 (.A(in_a[3]), .B(n_0_1_356), .CI(n_0_1_4), .CO(n_0_1_5), 
      .S(n_0_1_170));
   FA_X1 i_0_1_3 (.A(in_a[4]), .B(n_0_1_355), .CI(n_0_1_5), .CO(n_0_1_6), 
      .S(n_0_1_171));
   FA_X1 i_0_1_4 (.A(in_a[5]), .B(n_0_1_354), .CI(n_0_1_6), .CO(n_0_1_7), 
      .S(n_0_1_172));
   FA_X1 i_0_1_5 (.A(in_a[6]), .B(n_0_1_561), .CI(n_0_1_7), .CO(n_0_1_8), 
      .S(n_0_1_173));
   FA_X1 i_0_1_6 (.A(in_a[7]), .B(n_0_1_573), .CI(n_0_1_8), .CO(n_0_1_9), 
      .S(n_0_1_174));
   FA_X1 i_0_1_7 (.A(in_a[8]), .B(n_0_1_585), .CI(n_0_1_9), .CO(n_0_1_10), 
      .S(n_0_1_175));
   FA_X1 i_0_1_8 (.A(in_a[9]), .B(n_0_1_597), .CI(n_0_1_10), .CO(n_0_1_11), 
      .S(n_0_1_176));
   FA_X1 i_0_1_9 (.A(in_a[10]), .B(n_0_1_609), .CI(n_0_1_11), .CO(n_0_1_12), 
      .S(n_0_1_177));
   FA_X1 i_0_1_10 (.A(in_a[11]), .B(n_0_1_621), .CI(n_0_1_12), .CO(n_0_1_13), 
      .S(n_0_1_178));
   FA_X1 i_0_1_11 (.A(in_a[12]), .B(n_0_1_633), .CI(n_0_1_13), .CO(n_0_1_14), 
      .S(n_0_1_179));
   FA_X1 i_0_1_12 (.A(in_a[13]), .B(n_0_1_769), .CI(n_0_1_14), .CO(n_0_1_15), 
      .S(n_0_1_180));
   FA_X1 i_0_1_13 (.A(n_0_445), .B(n_0_1_358), .CI(n_0_1_157), .CO(n_0_1_0), 
      .S(n_0_1_181));
   FA_X1 i_0_1_14 (.A(n_0_446), .B(n_0_1_357), .CI(n_0_1_0), .CO(n_0_1_1), 
      .S(n_0_1_182));
   FA_X1 i_0_1_15 (.A(n_0_447), .B(n_0_1_356), .CI(n_0_1_1), .CO(n_0_1_2), 
      .S(n_0_1_183));
   FA_X1 i_0_1_16 (.A(n_0_448), .B(n_0_1_355), .CI(n_0_1_2), .CO(n_0_1_16), 
      .S(n_0_1_184));
   FA_X1 i_0_1_17 (.A(n_0_449), .B(n_0_1_354), .CI(n_0_1_16), .CO(n_0_1_17), 
      .S(n_0_1_185));
   FA_X1 i_0_1_18 (.A(n_0_450), .B(n_0_1_561), .CI(n_0_1_17), .CO(n_0_1_18), 
      .S(n_0_1_186));
   FA_X1 i_0_1_19 (.A(n_0_451), .B(n_0_1_573), .CI(n_0_1_18), .CO(n_0_1_19), 
      .S(n_0_1_187));
   FA_X1 i_0_1_20 (.A(n_0_452), .B(n_0_1_585), .CI(n_0_1_19), .CO(n_0_1_20), 
      .S(n_0_1_188));
   FA_X1 i_0_1_21 (.A(n_0_453), .B(n_0_1_597), .CI(n_0_1_20), .CO(n_0_1_21), 
      .S(n_0_1_189));
   FA_X1 i_0_1_22 (.A(n_0_454), .B(n_0_1_609), .CI(n_0_1_21), .CO(n_0_1_22), 
      .S(n_0_1_190));
   FA_X1 i_0_1_23 (.A(n_0_455), .B(n_0_1_621), .CI(n_0_1_22), .CO(n_0_1_23), 
      .S(n_0_1_191));
   FA_X1 i_0_1_24 (.A(n_0_456), .B(n_0_1_633), .CI(n_0_1_23), .CO(n_0_1_24), 
      .S(n_0_1_192));
   FA_X1 i_0_1_25 (.A(n_0_457), .B(n_0_1_769), .CI(n_0_1_24), .CO(n_0_1_25), 
      .S(n_0_1_193));
   FA_X1 i_0_1_26 (.A(in_a[1]), .B(n_0_1_350), .CI(n_0_1_159), .CO(n_0_1_26), 
      .S(n_0_1_194));
   FA_X1 i_0_1_27 (.A(in_a[2]), .B(n_0_1_348), .CI(n_0_1_26), .CO(n_0_1_27), 
      .S(n_0_1_195));
   FA_X1 i_0_1_28 (.A(in_a[3]), .B(n_0_1_346), .CI(n_0_1_27), .CO(n_0_1_28), 
      .S(n_0_1_196));
   FA_X1 i_0_1_29 (.A(in_a[4]), .B(n_0_1_344), .CI(n_0_1_28), .CO(n_0_1_29), 
      .S(n_0_1_197));
   FA_X1 i_0_1_30 (.A(in_a[5]), .B(n_0_1_559), .CI(n_0_1_29), .CO(n_0_1_30), 
      .S(n_0_1_198));
   FA_X1 i_0_1_31 (.A(in_a[6]), .B(n_0_1_571), .CI(n_0_1_30), .CO(n_0_1_31), 
      .S(n_0_1_199));
   FA_X1 i_0_1_32 (.A(in_a[7]), .B(n_0_1_583), .CI(n_0_1_31), .CO(n_0_1_32), 
      .S(n_0_1_200));
   FA_X1 i_0_1_33 (.A(in_a[8]), .B(n_0_1_595), .CI(n_0_1_32), .CO(n_0_1_33), 
      .S(n_0_1_201));
   FA_X1 i_0_1_34 (.A(in_a[9]), .B(n_0_1_607), .CI(n_0_1_33), .CO(n_0_1_34), 
      .S(n_0_1_202));
   FA_X1 i_0_1_35 (.A(in_a[10]), .B(n_0_1_619), .CI(n_0_1_34), .CO(n_0_1_35), 
      .S(n_0_1_203));
   FA_X1 i_0_1_36 (.A(in_a[11]), .B(n_0_1_631), .CI(n_0_1_35), .CO(n_0_1_36), 
      .S(n_0_1_204));
   FA_X1 i_0_1_37 (.A(in_a[12]), .B(n_0_1_643), .CI(n_0_1_36), .CO(n_0_1_37), 
      .S(n_0_1_205));
   FA_X1 i_0_1_38 (.A(in_a[13]), .B(n_0_1_654), .CI(n_0_1_37), .CO(n_0_1_38), 
      .S(n_0_1_206));
   FA_X1 i_0_1_39 (.A(n_0_445), .B(n_0_1_350), .CI(n_0_1_159), .CO(n_0_1_39), 
      .S(n_0_1_207));
   FA_X1 i_0_1_40 (.A(n_0_446), .B(n_0_1_348), .CI(n_0_1_39), .CO(n_0_1_40), 
      .S(n_0_1_208));
   FA_X1 i_0_1_41 (.A(n_0_447), .B(n_0_1_346), .CI(n_0_1_40), .CO(n_0_1_41), 
      .S(n_0_1_209));
   FA_X1 i_0_1_42 (.A(n_0_448), .B(n_0_1_344), .CI(n_0_1_41), .CO(n_0_1_42), 
      .S(n_0_1_210));
   FA_X1 i_0_1_43 (.A(n_0_449), .B(n_0_1_559), .CI(n_0_1_42), .CO(n_0_1_43), 
      .S(n_0_1_211));
   FA_X1 i_0_1_44 (.A(n_0_450), .B(n_0_1_571), .CI(n_0_1_43), .CO(n_0_1_44), 
      .S(n_0_1_212));
   FA_X1 i_0_1_45 (.A(n_0_451), .B(n_0_1_583), .CI(n_0_1_44), .CO(n_0_1_45), 
      .S(n_0_1_213));
   FA_X1 i_0_1_46 (.A(n_0_452), .B(n_0_1_595), .CI(n_0_1_45), .CO(n_0_1_46), 
      .S(n_0_1_214));
   FA_X1 i_0_1_47 (.A(n_0_453), .B(n_0_1_607), .CI(n_0_1_46), .CO(n_0_1_47), 
      .S(n_0_1_215));
   FA_X1 i_0_1_48 (.A(n_0_454), .B(n_0_1_619), .CI(n_0_1_47), .CO(n_0_1_48), 
      .S(n_0_1_216));
   FA_X1 i_0_1_49 (.A(n_0_455), .B(n_0_1_631), .CI(n_0_1_48), .CO(n_0_1_49), 
      .S(n_0_1_217));
   FA_X1 i_0_1_50 (.A(n_0_456), .B(n_0_1_643), .CI(n_0_1_49), .CO(n_0_1_50), 
      .S(n_0_1_218));
   FA_X1 i_0_1_51 (.A(n_0_457), .B(n_0_1_654), .CI(n_0_1_50), .CO(n_0_1_51), 
      .S(n_0_1_219));
   FA_X1 i_0_1_52 (.A(in_a[1]), .B(n_0_1_340), .CI(n_0_1_161), .CO(n_0_1_52), 
      .S(n_0_1_220));
   FA_X1 i_0_1_53 (.A(in_a[2]), .B(n_0_1_338), .CI(n_0_1_52), .CO(n_0_1_53), 
      .S(n_0_1_221));
   FA_X1 i_0_1_54 (.A(in_a[3]), .B(n_0_1_336), .CI(n_0_1_53), .CO(n_0_1_54), 
      .S(n_0_1_222));
   FA_X1 i_0_1_55 (.A(in_a[4]), .B(n_0_1_557), .CI(n_0_1_54), .CO(n_0_1_55), 
      .S(n_0_1_223));
   FA_X1 i_0_1_56 (.A(in_a[5]), .B(n_0_1_569), .CI(n_0_1_55), .CO(n_0_1_56), 
      .S(n_0_1_224));
   FA_X1 i_0_1_57 (.A(in_a[6]), .B(n_0_1_581), .CI(n_0_1_56), .CO(n_0_1_57), 
      .S(n_0_1_225));
   FA_X1 i_0_1_58 (.A(in_a[7]), .B(n_0_1_593), .CI(n_0_1_57), .CO(n_0_1_58), 
      .S(n_0_1_226));
   FA_X1 i_0_1_59 (.A(in_a[8]), .B(n_0_1_605), .CI(n_0_1_58), .CO(n_0_1_59), 
      .S(n_0_1_227));
   FA_X1 i_0_1_60 (.A(in_a[9]), .B(n_0_1_617), .CI(n_0_1_59), .CO(n_0_1_60), 
      .S(n_0_1_228));
   FA_X1 i_0_1_61 (.A(in_a[10]), .B(n_0_1_629), .CI(n_0_1_60), .CO(n_0_1_61), 
      .S(n_0_1_229));
   FA_X1 i_0_1_62 (.A(in_a[11]), .B(n_0_1_641), .CI(n_0_1_61), .CO(n_0_1_62), 
      .S(n_0_1_230));
   FA_X1 i_0_1_63 (.A(in_a[12]), .B(n_0_1_652), .CI(n_0_1_62), .CO(n_0_1_63), 
      .S(n_0_1_231));
   FA_X1 i_0_1_64 (.A(in_a[13]), .B(n_0_1_668), .CI(n_0_1_63), .CO(n_0_1_64), 
      .S(n_0_1_232));
   FA_X1 i_0_1_65 (.A(n_0_445), .B(n_0_1_340), .CI(n_0_1_161), .CO(n_0_1_65), 
      .S(n_0_1_233));
   FA_X1 i_0_1_66 (.A(n_0_446), .B(n_0_1_338), .CI(n_0_1_65), .CO(n_0_1_66), 
      .S(n_0_1_234));
   FA_X1 i_0_1_67 (.A(n_0_447), .B(n_0_1_336), .CI(n_0_1_66), .CO(n_0_1_67), 
      .S(n_0_1_235));
   FA_X1 i_0_1_68 (.A(n_0_448), .B(n_0_1_557), .CI(n_0_1_67), .CO(n_0_1_68), 
      .S(n_0_1_236));
   FA_X1 i_0_1_69 (.A(n_0_449), .B(n_0_1_569), .CI(n_0_1_68), .CO(n_0_1_69), 
      .S(n_0_1_237));
   FA_X1 i_0_1_70 (.A(n_0_450), .B(n_0_1_581), .CI(n_0_1_69), .CO(n_0_1_70), 
      .S(n_0_1_238));
   FA_X1 i_0_1_71 (.A(n_0_451), .B(n_0_1_593), .CI(n_0_1_70), .CO(n_0_1_71), 
      .S(n_0_1_239));
   FA_X1 i_0_1_72 (.A(n_0_452), .B(n_0_1_605), .CI(n_0_1_71), .CO(n_0_1_72), 
      .S(n_0_1_240));
   FA_X1 i_0_1_73 (.A(n_0_453), .B(n_0_1_617), .CI(n_0_1_72), .CO(n_0_1_73), 
      .S(n_0_1_241));
   FA_X1 i_0_1_74 (.A(n_0_454), .B(n_0_1_629), .CI(n_0_1_73), .CO(n_0_1_74), 
      .S(n_0_1_242));
   FA_X1 i_0_1_75 (.A(n_0_455), .B(n_0_1_641), .CI(n_0_1_74), .CO(n_0_1_75), 
      .S(n_0_1_243));
   FA_X1 i_0_1_76 (.A(n_0_456), .B(n_0_1_652), .CI(n_0_1_75), .CO(n_0_1_76), 
      .S(n_0_1_244));
   FA_X1 i_0_1_77 (.A(n_0_457), .B(n_0_1_668), .CI(n_0_1_76), .CO(n_0_1_77), 
      .S(n_0_1_245));
   FA_X1 i_0_1_78 (.A(in_a[1]), .B(n_0_1_332), .CI(n_0_1_163), .CO(n_0_1_78), 
      .S(n_0_1_246));
   FA_X1 i_0_1_79 (.A(in_a[2]), .B(n_0_1_330), .CI(n_0_1_78), .CO(n_0_1_79), 
      .S(n_0_1_247));
   FA_X1 i_0_1_80 (.A(in_a[3]), .B(n_0_1_555), .CI(n_0_1_79), .CO(n_0_1_80), 
      .S(n_0_1_248));
   FA_X1 i_0_1_81 (.A(in_a[4]), .B(n_0_1_567), .CI(n_0_1_80), .CO(n_0_1_81), 
      .S(n_0_1_249));
   FA_X1 i_0_1_82 (.A(in_a[5]), .B(n_0_1_579), .CI(n_0_1_81), .CO(n_0_1_82), 
      .S(n_0_1_250));
   FA_X1 i_0_1_83 (.A(in_a[6]), .B(n_0_1_591), .CI(n_0_1_82), .CO(n_0_1_83), 
      .S(n_0_1_251));
   FA_X1 i_0_1_84 (.A(in_a[7]), .B(n_0_1_603), .CI(n_0_1_83), .CO(n_0_1_84), 
      .S(n_0_1_252));
   FA_X1 i_0_1_85 (.A(in_a[8]), .B(n_0_1_615), .CI(n_0_1_84), .CO(n_0_1_85), 
      .S(n_0_1_253));
   FA_X1 i_0_1_86 (.A(in_a[9]), .B(n_0_1_627), .CI(n_0_1_85), .CO(n_0_1_86), 
      .S(n_0_1_254));
   FA_X1 i_0_1_87 (.A(in_a[10]), .B(n_0_1_639), .CI(n_0_1_86), .CO(n_0_1_87), 
      .S(n_0_1_255));
   FA_X1 i_0_1_88 (.A(in_a[11]), .B(n_0_1_650), .CI(n_0_1_87), .CO(n_0_1_88), 
      .S(n_0_1_256));
   FA_X1 i_0_1_89 (.A(in_a[12]), .B(n_0_1_666), .CI(n_0_1_88), .CO(n_0_1_89), 
      .S(n_0_1_257));
   FA_X1 i_0_1_90 (.A(in_a[13]), .B(n_0_1_679), .CI(n_0_1_89), .CO(n_0_1_90), 
      .S(n_0_1_258));
   FA_X1 i_0_1_91 (.A(n_0_445), .B(n_0_1_332), .CI(n_0_1_163), .CO(n_0_1_91), 
      .S(n_0_1_259));
   FA_X1 i_0_1_92 (.A(n_0_446), .B(n_0_1_330), .CI(n_0_1_91), .CO(n_0_1_92), 
      .S(n_0_1_260));
   FA_X1 i_0_1_93 (.A(n_0_447), .B(n_0_1_555), .CI(n_0_1_92), .CO(n_0_1_93), 
      .S(n_0_1_261));
   FA_X1 i_0_1_94 (.A(n_0_448), .B(n_0_1_567), .CI(n_0_1_93), .CO(n_0_1_94), 
      .S(n_0_1_262));
   FA_X1 i_0_1_95 (.A(n_0_449), .B(n_0_1_579), .CI(n_0_1_94), .CO(n_0_1_95), 
      .S(n_0_1_263));
   FA_X1 i_0_1_96 (.A(n_0_450), .B(n_0_1_591), .CI(n_0_1_95), .CO(n_0_1_96), 
      .S(n_0_1_264));
   FA_X1 i_0_1_97 (.A(n_0_451), .B(n_0_1_603), .CI(n_0_1_96), .CO(n_0_1_97), 
      .S(n_0_1_265));
   FA_X1 i_0_1_98 (.A(n_0_452), .B(n_0_1_615), .CI(n_0_1_97), .CO(n_0_1_98), 
      .S(n_0_1_266));
   FA_X1 i_0_1_99 (.A(n_0_453), .B(n_0_1_627), .CI(n_0_1_98), .CO(n_0_1_99), 
      .S(n_0_1_267));
   FA_X1 i_0_1_100 (.A(n_0_454), .B(n_0_1_639), .CI(n_0_1_99), .CO(n_0_1_100), 
      .S(n_0_1_268));
   FA_X1 i_0_1_101 (.A(n_0_455), .B(n_0_1_650), .CI(n_0_1_100), .CO(n_0_1_101), 
      .S(n_0_1_269));
   FA_X1 i_0_1_102 (.A(n_0_456), .B(n_0_1_666), .CI(n_0_1_101), .CO(n_0_1_102), 
      .S(n_0_1_270));
   FA_X1 i_0_1_103 (.A(n_0_457), .B(n_0_1_679), .CI(n_0_1_102), .CO(n_0_1_103), 
      .S(n_0_1_271));
   FA_X1 i_0_1_104 (.A(in_a[1]), .B(n_0_1_326), .CI(n_0_1_165), .CO(n_0_1_104), 
      .S(n_0_1_272));
   FA_X1 i_0_1_105 (.A(in_a[2]), .B(n_0_1_553), .CI(n_0_1_104), .CO(n_0_1_105), 
      .S(n_0_1_273));
   FA_X1 i_0_1_106 (.A(in_a[3]), .B(n_0_1_565), .CI(n_0_1_105), .CO(n_0_1_106), 
      .S(n_0_1_274));
   FA_X1 i_0_1_107 (.A(in_a[4]), .B(n_0_1_577), .CI(n_0_1_106), .CO(n_0_1_107), 
      .S(n_0_1_275));
   FA_X1 i_0_1_108 (.A(in_a[5]), .B(n_0_1_589), .CI(n_0_1_107), .CO(n_0_1_108), 
      .S(n_0_1_276));
   FA_X1 i_0_1_109 (.A(in_a[6]), .B(n_0_1_601), .CI(n_0_1_108), .CO(n_0_1_109), 
      .S(n_0_1_277));
   FA_X1 i_0_1_110 (.A(in_a[7]), .B(n_0_1_613), .CI(n_0_1_109), .CO(n_0_1_110), 
      .S(n_0_1_278));
   FA_X1 i_0_1_111 (.A(in_a[8]), .B(n_0_1_625), .CI(n_0_1_110), .CO(n_0_1_111), 
      .S(n_0_1_279));
   FA_X1 i_0_1_112 (.A(in_a[9]), .B(n_0_1_637), .CI(n_0_1_111), .CO(n_0_1_112), 
      .S(n_0_1_280));
   FA_X1 i_0_1_113 (.A(in_a[10]), .B(n_0_1_648), .CI(n_0_1_112), .CO(n_0_1_113), 
      .S(n_0_1_281));
   FA_X1 i_0_1_114 (.A(in_a[11]), .B(n_0_1_664), .CI(n_0_1_113), .CO(n_0_1_114), 
      .S(n_0_1_282));
   FA_X1 i_0_1_115 (.A(in_a[12]), .B(n_0_1_677), .CI(n_0_1_114), .CO(n_0_1_115), 
      .S(n_0_1_283));
   FA_X1 i_0_1_116 (.A(in_a[13]), .B(n_0_1_686), .CI(n_0_1_115), .CO(n_0_1_116), 
      .S(n_0_1_284));
   FA_X1 i_0_1_117 (.A(n_0_445), .B(n_0_1_326), .CI(n_0_1_165), .CO(n_0_1_117), 
      .S(n_0_1_285));
   FA_X1 i_0_1_118 (.A(n_0_446), .B(n_0_1_553), .CI(n_0_1_117), .CO(n_0_1_118), 
      .S(n_0_1_286));
   FA_X1 i_0_1_119 (.A(n_0_447), .B(n_0_1_565), .CI(n_0_1_118), .CO(n_0_1_119), 
      .S(n_0_1_287));
   FA_X1 i_0_1_120 (.A(n_0_448), .B(n_0_1_577), .CI(n_0_1_119), .CO(n_0_1_120), 
      .S(n_0_1_288));
   FA_X1 i_0_1_121 (.A(n_0_449), .B(n_0_1_589), .CI(n_0_1_120), .CO(n_0_1_121), 
      .S(n_0_1_289));
   FA_X1 i_0_1_122 (.A(n_0_450), .B(n_0_1_601), .CI(n_0_1_121), .CO(n_0_1_122), 
      .S(n_0_1_290));
   FA_X1 i_0_1_123 (.A(n_0_451), .B(n_0_1_613), .CI(n_0_1_122), .CO(n_0_1_123), 
      .S(n_0_1_291));
   FA_X1 i_0_1_124 (.A(n_0_452), .B(n_0_1_625), .CI(n_0_1_123), .CO(n_0_1_124), 
      .S(n_0_1_292));
   FA_X1 i_0_1_125 (.A(n_0_453), .B(n_0_1_637), .CI(n_0_1_124), .CO(n_0_1_125), 
      .S(n_0_1_293));
   FA_X1 i_0_1_126 (.A(n_0_454), .B(n_0_1_648), .CI(n_0_1_125), .CO(n_0_1_126), 
      .S(n_0_1_294));
   FA_X1 i_0_1_127 (.A(n_0_455), .B(n_0_1_664), .CI(n_0_1_126), .CO(n_0_1_127), 
      .S(n_0_1_295));
   FA_X1 i_0_1_128 (.A(n_0_456), .B(n_0_1_677), .CI(n_0_1_127), .CO(n_0_1_128), 
      .S(n_0_1_296));
   FA_X1 i_0_1_129 (.A(n_0_457), .B(n_0_1_686), .CI(n_0_1_128), .CO(n_0_1_129), 
      .S(n_0_1_297));
   FA_X1 i_0_1_130 (.A(in_a[1]), .B(n_0_1_551), .CI(n_0_1_167), .CO(n_0_1_130), 
      .S(n_0_1_298));
   FA_X1 i_0_1_131 (.A(in_a[2]), .B(n_0_1_563), .CI(n_0_1_130), .CO(n_0_1_131), 
      .S(n_0_1_299));
   FA_X1 i_0_1_132 (.A(in_a[3]), .B(n_0_1_575), .CI(n_0_1_131), .CO(n_0_1_132), 
      .S(n_0_1_300));
   FA_X1 i_0_1_133 (.A(in_a[4]), .B(n_0_1_587), .CI(n_0_1_132), .CO(n_0_1_133), 
      .S(n_0_1_301));
   FA_X1 i_0_1_134 (.A(in_a[5]), .B(n_0_1_599), .CI(n_0_1_133), .CO(n_0_1_134), 
      .S(n_0_1_302));
   FA_X1 i_0_1_135 (.A(in_a[6]), .B(n_0_1_611), .CI(n_0_1_134), .CO(n_0_1_135), 
      .S(n_0_1_303));
   FA_X1 i_0_1_136 (.A(in_a[7]), .B(n_0_1_623), .CI(n_0_1_135), .CO(n_0_1_136), 
      .S(n_0_1_304));
   FA_X1 i_0_1_137 (.A(in_a[8]), .B(n_0_1_635), .CI(n_0_1_136), .CO(n_0_1_137), 
      .S(n_0_1_305));
   FA_X1 i_0_1_138 (.A(in_a[9]), .B(n_0_1_646), .CI(n_0_1_137), .CO(n_0_1_138), 
      .S(n_0_1_306));
   FA_X1 i_0_1_139 (.A(in_a[10]), .B(n_0_1_662), .CI(n_0_1_138), .CO(n_0_1_139), 
      .S(n_0_1_307));
   FA_X1 i_0_1_140 (.A(in_a[11]), .B(n_0_1_675), .CI(n_0_1_139), .CO(n_0_1_140), 
      .S(n_0_1_308));
   FA_X1 i_0_1_141 (.A(in_a[12]), .B(n_0_1_684), .CI(n_0_1_140), .CO(n_0_1_141), 
      .S(n_0_1_309));
   FA_X1 i_0_1_142 (.A(in_a[13]), .B(n_0_1_691), .CI(n_0_1_141), .CO(n_0_1_142), 
      .S(n_0_1_310));
   FA_X1 i_0_1_143 (.A(n_0_445), .B(n_0_1_551), .CI(n_0_1_167), .CO(n_0_1_143), 
      .S(n_0_1_311));
   FA_X1 i_0_1_144 (.A(n_0_446), .B(n_0_1_563), .CI(n_0_1_143), .CO(n_0_1_144), 
      .S(n_0_1_312));
   FA_X1 i_0_1_145 (.A(n_0_447), .B(n_0_1_575), .CI(n_0_1_144), .CO(n_0_1_145), 
      .S(n_0_1_313));
   FA_X1 i_0_1_146 (.A(n_0_448), .B(n_0_1_587), .CI(n_0_1_145), .CO(n_0_1_146), 
      .S(n_0_1_314));
   FA_X1 i_0_1_147 (.A(n_0_449), .B(n_0_1_599), .CI(n_0_1_146), .CO(n_0_1_147), 
      .S(n_0_1_315));
   FA_X1 i_0_1_148 (.A(n_0_450), .B(n_0_1_611), .CI(n_0_1_147), .CO(n_0_1_148), 
      .S(n_0_1_316));
   FA_X1 i_0_1_149 (.A(n_0_451), .B(n_0_1_623), .CI(n_0_1_148), .CO(n_0_1_149), 
      .S(n_0_1_317));
   FA_X1 i_0_1_150 (.A(n_0_452), .B(n_0_1_635), .CI(n_0_1_149), .CO(n_0_1_150), 
      .S(n_0_1_318));
   FA_X1 i_0_1_151 (.A(n_0_453), .B(n_0_1_646), .CI(n_0_1_150), .CO(n_0_1_151), 
      .S(n_0_1_319));
   FA_X1 i_0_1_152 (.A(n_0_454), .B(n_0_1_662), .CI(n_0_1_151), .CO(n_0_1_152), 
      .S(n_0_1_320));
   FA_X1 i_0_1_153 (.A(n_0_455), .B(n_0_1_675), .CI(n_0_1_152), .CO(n_0_1_153), 
      .S(n_0_1_321));
   FA_X1 i_0_1_154 (.A(n_0_456), .B(n_0_1_684), .CI(n_0_1_153), .CO(n_0_1_154), 
      .S(n_0_1_322));
   FA_X1 i_0_1_155 (.A(n_0_457), .B(n_0_1_691), .CI(n_0_1_154), .CO(n_0_1_155), 
      .S(n_0_1_323));
   HA_X1 i_0_1_156 (.A(in_a[0]), .B(n_0_1_359), .CO(n_0_1_157), .S(n_0_1_156));
   HA_X1 i_0_1_157 (.A(in_a[0]), .B(n_0_1_352), .CO(n_0_1_159), .S(n_0_1_158));
   HA_X1 i_0_1_158 (.A(in_a[0]), .B(n_0_1_342), .CO(n_0_1_161), .S(n_0_1_160));
   HA_X1 i_0_1_159 (.A(in_a[0]), .B(n_0_1_334), .CO(n_0_1_163), .S(n_0_1_162));
   HA_X1 i_0_1_160 (.A(in_a[0]), .B(n_0_1_328), .CO(n_0_1_165), .S(n_0_1_164));
   HA_X1 i_0_1_161 (.A(in_a[0]), .B(n_0_1_324), .CO(n_0_1_167), .S(n_0_1_166));
   INV_X1 i_0_1_162 (.A(n_0_1_325), .ZN(n_0_1_324));
   AOI222_X1 i_0_1_163 (.A1(n_0_1_272), .A2(n_0_1_717), .B1(n_0_1_285), .B2(
      n_0_1_719), .C1(n_0_1_716), .C2(n_0_1_326), .ZN(n_0_1_325));
   INV_X1 i_0_1_164 (.A(n_0_1_327), .ZN(n_0_1_326));
   AOI222_X1 i_0_1_165 (.A1(n_0_1_247), .A2(n_0_1_730), .B1(n_0_1_260), .B2(
      n_0_1_728), .C1(n_0_1_727), .C2(n_0_1_330), .ZN(n_0_1_327));
   INV_X1 i_0_1_166 (.A(n_0_1_329), .ZN(n_0_1_328));
   AOI222_X1 i_0_1_167 (.A1(n_0_1_246), .A2(n_0_1_730), .B1(n_0_1_259), .B2(
      n_0_1_728), .C1(n_0_1_727), .C2(n_0_1_332), .ZN(n_0_1_329));
   INV_X1 i_0_1_168 (.A(n_0_1_331), .ZN(n_0_1_330));
   AOI222_X1 i_0_1_169 (.A1(n_0_1_222), .A2(n_0_1_739), .B1(n_0_1_235), .B2(
      n_0_1_741), .C1(n_0_1_738), .C2(n_0_1_336), .ZN(n_0_1_331));
   INV_X1 i_0_1_170 (.A(n_0_1_333), .ZN(n_0_1_332));
   AOI222_X1 i_0_1_171 (.A1(n_0_1_221), .A2(n_0_1_739), .B1(n_0_1_234), .B2(
      n_0_1_741), .C1(n_0_1_738), .C2(n_0_1_338), .ZN(n_0_1_333));
   INV_X1 i_0_1_172 (.A(n_0_1_335), .ZN(n_0_1_334));
   AOI222_X1 i_0_1_173 (.A1(n_0_1_220), .A2(n_0_1_739), .B1(n_0_1_233), .B2(
      n_0_1_741), .C1(n_0_1_738), .C2(n_0_1_340), .ZN(n_0_1_335));
   INV_X1 i_0_1_174 (.A(n_0_1_337), .ZN(n_0_1_336));
   AOI222_X1 i_0_1_175 (.A1(n_0_1_197), .A2(n_0_1_751), .B1(n_0_1_210), .B2(
      n_0_1_753), .C1(n_0_1_750), .C2(n_0_1_344), .ZN(n_0_1_337));
   INV_X1 i_0_1_176 (.A(n_0_1_339), .ZN(n_0_1_338));
   AOI222_X1 i_0_1_177 (.A1(n_0_1_196), .A2(n_0_1_751), .B1(n_0_1_209), .B2(
      n_0_1_753), .C1(n_0_1_750), .C2(n_0_1_346), .ZN(n_0_1_339));
   INV_X1 i_0_1_178 (.A(n_0_1_341), .ZN(n_0_1_340));
   AOI222_X1 i_0_1_179 (.A1(n_0_1_195), .A2(n_0_1_751), .B1(n_0_1_208), .B2(
      n_0_1_753), .C1(n_0_1_750), .C2(n_0_1_348), .ZN(n_0_1_341));
   INV_X1 i_0_1_180 (.A(n_0_1_343), .ZN(n_0_1_342));
   AOI222_X1 i_0_1_181 (.A1(n_0_1_194), .A2(n_0_1_751), .B1(n_0_1_207), .B2(
      n_0_1_753), .C1(n_0_1_750), .C2(n_0_1_350), .ZN(n_0_1_343));
   INV_X1 i_0_1_182 (.A(n_0_1_345), .ZN(n_0_1_344));
   AOI222_X1 i_0_1_183 (.A1(n_0_1_172), .A2(n_0_1_763), .B1(n_0_1_185), .B2(
      n_0_1_765), .C1(n_0_1_762), .C2(n_0_1_354), .ZN(n_0_1_345));
   INV_X1 i_0_1_184 (.A(n_0_1_347), .ZN(n_0_1_346));
   AOI222_X1 i_0_1_185 (.A1(n_0_1_171), .A2(n_0_1_763), .B1(n_0_1_184), .B2(
      n_0_1_765), .C1(n_0_1_762), .C2(n_0_1_355), .ZN(n_0_1_347));
   INV_X1 i_0_1_186 (.A(n_0_1_349), .ZN(n_0_1_348));
   AOI222_X1 i_0_1_187 (.A1(n_0_1_170), .A2(n_0_1_763), .B1(n_0_1_183), .B2(
      n_0_1_765), .C1(n_0_1_762), .C2(n_0_1_356), .ZN(n_0_1_349));
   INV_X1 i_0_1_188 (.A(n_0_1_351), .ZN(n_0_1_350));
   AOI222_X1 i_0_1_189 (.A1(n_0_1_169), .A2(n_0_1_763), .B1(n_0_1_182), .B2(
      n_0_1_765), .C1(n_0_1_762), .C2(n_0_1_357), .ZN(n_0_1_351));
   INV_X1 i_0_1_190 (.A(n_0_1_353), .ZN(n_0_1_352));
   AOI222_X1 i_0_1_191 (.A1(n_0_1_168), .A2(n_0_1_763), .B1(n_0_1_181), .B2(
      n_0_1_765), .C1(n_0_1_762), .C2(n_0_1_358), .ZN(n_0_1_353));
   AND2_X1 i_0_1_192 (.A1(in_b[0]), .A2(n_0_450), .ZN(n_0_1_354));
   AND2_X1 i_0_1_193 (.A1(in_b[0]), .A2(n_0_449), .ZN(n_0_1_355));
   AND2_X1 i_0_1_194 (.A1(in_b[0]), .A2(n_0_448), .ZN(n_0_1_356));
   AND2_X1 i_0_1_195 (.A1(in_b[0]), .A2(n_0_447), .ZN(n_0_1_357));
   AND2_X1 i_0_1_196 (.A1(in_b[0]), .A2(n_0_446), .ZN(n_0_1_358));
   AND2_X1 i_0_1_197 (.A1(in_b[0]), .A2(n_0_445), .ZN(n_0_1_359));
   AOI22_X1 i_0_1_198 (.A1(n_0_1_369), .A2(n_0_1_363), .B1(n_0_1_368), .B2(
      n_0_1_360), .ZN(n_0_291));
   NOR2_X1 i_0_1_199 (.A1(n_0_1_362), .A2(n_0_1_361), .ZN(n_0_1_360));
   NAND4_X1 i_0_1_200 (.A1(n_0_1_370), .A2(n_0_1_365), .A3(n_0_1_393), .A4(
      n_0_1_367), .ZN(n_0_1_361));
   NAND4_X1 i_0_1_201 (.A1(n_0_1_372), .A2(n_0_1_371), .A3(n_0_1_392), .A4(
      n_0_1_366), .ZN(n_0_1_362));
   AND3_X1 i_0_1_202 (.A1(\output ), .A2(n_0_309), .A3(n_0_1_364), .ZN(n_0_1_363));
   NOR4_X1 i_0_1_203 (.A1(n_0_1_368), .A2(n_0_1_367), .A3(n_0_1_366), .A4(
      n_0_1_365), .ZN(n_0_1_364));
   AOI222_X1 i_0_1_204 (.A1(n_0_283), .A2(n_0_1_396), .B1(n_0_267), .B2(
      n_0_1_397), .C1(n_0_320), .C2(n_0_1_395), .ZN(n_0_1_365));
   AOI221_X1 i_0_1_205 (.A(n_0_1_394), .B1(n_0_271), .B2(n_0_1_397), .C1(n_0_287), 
      .C2(n_0_1_396), .ZN(n_0_1_366));
   AOI222_X1 i_0_1_206 (.A1(n_0_281), .A2(n_0_1_396), .B1(n_0_265), .B2(
      n_0_1_397), .C1(n_0_318), .C2(n_0_1_395), .ZN(n_0_1_367));
   AOI222_X1 i_0_1_207 (.A1(n_0_269), .A2(n_0_1_397), .B1(n_0_285), .B2(
      n_0_1_396), .C1(n_0_322), .C2(n_0_1_395), .ZN(n_0_1_368));
   NOR3_X1 i_0_1_208 (.A1(n_0_1_371), .A2(n_0_1_370), .A3(n_0_1_372), .ZN(
      n_0_1_369));
   AOI222_X1 i_0_1_209 (.A1(n_0_284), .A2(n_0_1_396), .B1(n_0_268), .B2(
      n_0_1_397), .C1(n_0_321), .C2(n_0_1_395), .ZN(n_0_1_370));
   AOI222_X1 i_0_1_210 (.A1(n_0_286), .A2(n_0_1_396), .B1(n_0_270), .B2(
      n_0_1_397), .C1(n_0_323), .C2(n_0_1_395), .ZN(n_0_1_371));
   AOI222_X1 i_0_1_211 (.A1(n_0_282), .A2(n_0_1_396), .B1(n_0_266), .B2(
      n_0_1_397), .C1(n_0_319), .C2(n_0_1_395), .ZN(n_0_1_372));
   NOR2_X1 i_0_1_212 (.A1(n_0_302), .A2(n_0_293), .ZN(n_0_292));
   NOR4_X1 i_0_1_213 (.A1(n_0_304), .A2(n_0_1_374), .A3(n_0_305), .A4(n_0_1_373), 
      .ZN(n_0_293));
   NAND4_X1 i_0_1_214 (.A1(n_0_1_390), .A2(n_0_1_389), .A3(n_0_1_391), .A4(
      n_0_1_392), .ZN(n_0_1_373));
   NAND4_X1 i_0_1_215 (.A1(n_0_1_384), .A2(n_0_1_375), .A3(n_0_1_385), .A4(
      n_0_1_386), .ZN(n_0_1_374));
   AND4_X1 i_0_1_216 (.A1(n_0_1_381), .A2(n_0_1_376), .A3(n_0_1_382), .A4(
      n_0_1_383), .ZN(n_0_1_375));
   NOR4_X1 i_0_1_217 (.A1(n_0_295), .A2(n_0_294), .A3(n_0_296), .A4(n_0_297), 
      .ZN(n_0_1_376));
   INV_X1 i_0_1_218 (.A(n_0_1_377), .ZN(n_0_294));
   AOI222_X1 i_0_1_219 (.A1(n_0_0), .A2(n_0_1_548), .B1(n_0_17), .B2(n_0_1_549), 
      .C1(n_0_430), .C2(n_0_1_547), .ZN(n_0_1_377));
   INV_X1 i_0_1_220 (.A(n_0_1_378), .ZN(n_0_295));
   AOI222_X1 i_0_1_221 (.A1(n_0_33), .A2(n_0_1_529), .B1(n_0_49), .B2(n_0_1_530), 
      .C1(n_0_415), .C2(n_0_1_528), .ZN(n_0_1_378));
   INV_X1 i_0_1_222 (.A(n_0_1_379), .ZN(n_0_296));
   AOI222_X1 i_0_1_223 (.A1(n_0_65), .A2(n_0_1_510), .B1(n_0_81), .B2(n_0_1_511), 
      .C1(n_0_400), .C2(n_0_1_509), .ZN(n_0_1_379));
   INV_X1 i_0_1_224 (.A(n_0_1_380), .ZN(n_0_297));
   AOI222_X1 i_0_1_225 (.A1(n_0_97), .A2(n_0_1_491), .B1(n_0_113), .B2(n_0_1_492), 
      .C1(n_0_385), .C2(n_0_1_490), .ZN(n_0_1_380));
   INV_X1 i_0_1_226 (.A(n_0_1_381), .ZN(n_0_298));
   AOI222_X1 i_0_1_227 (.A1(n_0_129), .A2(n_0_1_472), .B1(n_0_145), .B2(
      n_0_1_473), .C1(n_0_370), .C2(n_0_1_471), .ZN(n_0_1_381));
   INV_X1 i_0_1_228 (.A(n_0_1_382), .ZN(n_0_299));
   AOI222_X1 i_0_1_229 (.A1(n_0_161), .A2(n_0_1_453), .B1(n_0_177), .B2(
      n_0_1_454), .C1(n_0_355), .C2(n_0_1_452), .ZN(n_0_1_382));
   INV_X1 i_0_1_230 (.A(n_0_1_383), .ZN(n_0_300));
   AOI222_X1 i_0_1_231 (.A1(n_0_193), .A2(n_0_1_434), .B1(n_0_209), .B2(
      n_0_1_435), .C1(n_0_340), .C2(n_0_1_433), .ZN(n_0_1_383));
   INV_X1 i_0_1_232 (.A(n_0_1_384), .ZN(n_0_301));
   AOI222_X1 i_0_1_233 (.A1(n_0_225), .A2(n_0_1_415), .B1(n_0_241), .B2(
      n_0_1_416), .C1(n_0_325), .C2(n_0_1_414), .ZN(n_0_1_384));
   INV_X1 i_0_1_234 (.A(n_0_1_385), .ZN(n_0_302));
   AOI222_X1 i_0_1_235 (.A1(n_0_257), .A2(n_0_1_397), .B1(n_0_273), .B2(
      n_0_1_396), .C1(n_0_310), .C2(n_0_1_395), .ZN(n_0_1_385));
   INV_X1 i_0_1_236 (.A(n_0_1_386), .ZN(n_0_303));
   AOI222_X1 i_0_1_237 (.A1(n_0_258), .A2(n_0_1_397), .B1(n_0_274), .B2(
      n_0_1_396), .C1(n_0_311), .C2(n_0_1_395), .ZN(n_0_1_386));
   INV_X1 i_0_1_238 (.A(n_0_1_387), .ZN(n_0_304));
   AOI222_X1 i_0_1_239 (.A1(n_0_259), .A2(n_0_1_397), .B1(n_0_275), .B2(
      n_0_1_396), .C1(n_0_312), .C2(n_0_1_395), .ZN(n_0_1_387));
   INV_X1 i_0_1_240 (.A(n_0_1_388), .ZN(n_0_305));
   AOI222_X1 i_0_1_241 (.A1(n_0_260), .A2(n_0_1_397), .B1(n_0_276), .B2(
      n_0_1_396), .C1(n_0_313), .C2(n_0_1_395), .ZN(n_0_1_388));
   INV_X1 i_0_1_242 (.A(n_0_1_389), .ZN(n_0_306));
   AOI222_X1 i_0_1_243 (.A1(n_0_277), .A2(n_0_1_396), .B1(n_0_261), .B2(
      n_0_1_397), .C1(n_0_314), .C2(n_0_1_395), .ZN(n_0_1_389));
   INV_X1 i_0_1_244 (.A(n_0_1_390), .ZN(n_0_307));
   AOI222_X1 i_0_1_245 (.A1(n_0_278), .A2(n_0_1_396), .B1(n_0_262), .B2(
      n_0_1_397), .C1(n_0_315), .C2(n_0_1_395), .ZN(n_0_1_390));
   INV_X1 i_0_1_246 (.A(n_0_1_391), .ZN(n_0_308));
   AOI222_X1 i_0_1_247 (.A1(n_0_279), .A2(n_0_1_396), .B1(n_0_263), .B2(
      n_0_1_397), .C1(n_0_316), .C2(n_0_1_395), .ZN(n_0_1_391));
   INV_X1 i_0_1_248 (.A(n_0_1_392), .ZN(n_0_309));
   AOI222_X1 i_0_1_249 (.A1(n_0_280), .A2(n_0_1_396), .B1(n_0_264), .B2(
      n_0_1_397), .C1(n_0_317), .C2(n_0_1_395), .ZN(n_0_1_392));
   INV_X1 i_0_1_250 (.A(n_0_1_393), .ZN(\output ));
   AOI221_X1 i_0_1_251 (.A(n_0_1_394), .B1(n_0_272), .B2(n_0_1_397), .C1(n_0_288), 
      .C2(n_0_1_396), .ZN(n_0_1_393));
   AND2_X1 i_0_1_252 (.A1(n_0_324), .A2(n_0_1_395), .ZN(n_0_1_394));
   NOR2_X1 i_0_1_253 (.A1(n_0_1_397), .A2(n_0_1_396), .ZN(n_0_1_395));
   AND2_X1 i_0_1_254 (.A1(in_b[15]), .A2(n_0_1_827), .ZN(n_0_1_396));
   NOR2_X1 i_0_1_255 (.A1(in_b[15]), .A2(n_0_1_827), .ZN(n_0_1_397));
   INV_X1 i_0_1_256 (.A(n_0_1_398), .ZN(n_0_310));
   AOI222_X1 i_0_1_257 (.A1(n_0_226), .A2(n_0_1_415), .B1(n_0_242), .B2(
      n_0_1_416), .C1(n_0_326), .C2(n_0_1_414), .ZN(n_0_1_398));
   INV_X1 i_0_1_258 (.A(n_0_1_399), .ZN(n_0_311));
   AOI222_X1 i_0_1_259 (.A1(n_0_227), .A2(n_0_1_415), .B1(n_0_243), .B2(
      n_0_1_416), .C1(n_0_327), .C2(n_0_1_414), .ZN(n_0_1_399));
   INV_X1 i_0_1_260 (.A(n_0_1_400), .ZN(n_0_312));
   AOI222_X1 i_0_1_261 (.A1(n_0_228), .A2(n_0_1_415), .B1(n_0_244), .B2(
      n_0_1_416), .C1(n_0_328), .C2(n_0_1_414), .ZN(n_0_1_400));
   INV_X1 i_0_1_262 (.A(n_0_1_401), .ZN(n_0_313));
   AOI222_X1 i_0_1_263 (.A1(n_0_229), .A2(n_0_1_415), .B1(n_0_245), .B2(
      n_0_1_416), .C1(n_0_329), .C2(n_0_1_414), .ZN(n_0_1_401));
   INV_X1 i_0_1_264 (.A(n_0_1_402), .ZN(n_0_314));
   AOI222_X1 i_0_1_265 (.A1(n_0_246), .A2(n_0_1_416), .B1(n_0_230), .B2(
      n_0_1_415), .C1(n_0_330), .C2(n_0_1_414), .ZN(n_0_1_402));
   INV_X1 i_0_1_266 (.A(n_0_1_403), .ZN(n_0_315));
   AOI222_X1 i_0_1_267 (.A1(n_0_247), .A2(n_0_1_416), .B1(n_0_231), .B2(
      n_0_1_415), .C1(n_0_331), .C2(n_0_1_414), .ZN(n_0_1_403));
   INV_X1 i_0_1_268 (.A(n_0_1_404), .ZN(n_0_316));
   AOI222_X1 i_0_1_269 (.A1(n_0_248), .A2(n_0_1_416), .B1(n_0_232), .B2(
      n_0_1_415), .C1(n_0_332), .C2(n_0_1_414), .ZN(n_0_1_404));
   INV_X1 i_0_1_270 (.A(n_0_1_405), .ZN(n_0_317));
   AOI222_X1 i_0_1_271 (.A1(n_0_249), .A2(n_0_1_416), .B1(n_0_233), .B2(
      n_0_1_415), .C1(n_0_333), .C2(n_0_1_414), .ZN(n_0_1_405));
   INV_X1 i_0_1_272 (.A(n_0_1_406), .ZN(n_0_318));
   AOI222_X1 i_0_1_273 (.A1(n_0_250), .A2(n_0_1_416), .B1(n_0_234), .B2(
      n_0_1_415), .C1(n_0_334), .C2(n_0_1_414), .ZN(n_0_1_406));
   INV_X1 i_0_1_274 (.A(n_0_1_407), .ZN(n_0_319));
   AOI222_X1 i_0_1_275 (.A1(n_0_251), .A2(n_0_1_416), .B1(n_0_235), .B2(
      n_0_1_415), .C1(n_0_335), .C2(n_0_1_414), .ZN(n_0_1_407));
   INV_X1 i_0_1_276 (.A(n_0_1_408), .ZN(n_0_320));
   AOI222_X1 i_0_1_277 (.A1(n_0_252), .A2(n_0_1_416), .B1(n_0_236), .B2(
      n_0_1_415), .C1(n_0_336), .C2(n_0_1_414), .ZN(n_0_1_408));
   INV_X1 i_0_1_278 (.A(n_0_1_409), .ZN(n_0_321));
   AOI222_X1 i_0_1_279 (.A1(n_0_253), .A2(n_0_1_416), .B1(n_0_237), .B2(
      n_0_1_415), .C1(n_0_337), .C2(n_0_1_414), .ZN(n_0_1_409));
   INV_X1 i_0_1_280 (.A(n_0_1_410), .ZN(n_0_322));
   AOI222_X1 i_0_1_281 (.A1(n_0_238), .A2(n_0_1_415), .B1(n_0_254), .B2(
      n_0_1_416), .C1(n_0_338), .C2(n_0_1_414), .ZN(n_0_1_410));
   INV_X1 i_0_1_282 (.A(n_0_1_411), .ZN(n_0_323));
   AOI221_X1 i_0_1_283 (.A(n_0_1_413), .B1(n_0_239), .B2(n_0_1_415), .C1(n_0_255), 
      .C2(n_0_1_416), .ZN(n_0_1_411));
   INV_X1 i_0_1_284 (.A(n_0_1_412), .ZN(n_0_324));
   AOI221_X1 i_0_1_285 (.A(n_0_1_413), .B1(n_0_240), .B2(n_0_1_415), .C1(n_0_256), 
      .C2(n_0_1_416), .ZN(n_0_1_412));
   AND2_X1 i_0_1_286 (.A1(n_0_339), .A2(n_0_1_414), .ZN(n_0_1_413));
   NOR2_X1 i_0_1_287 (.A1(n_0_1_416), .A2(n_0_1_415), .ZN(n_0_1_414));
   NOR2_X1 i_0_1_288 (.A1(in_b[14]), .A2(n_0_1_826), .ZN(n_0_1_415));
   NOR2_X1 i_0_1_289 (.A1(n_0_1_827), .A2(in_b[13]), .ZN(n_0_1_416));
   INV_X1 i_0_1_290 (.A(n_0_1_417), .ZN(n_0_325));
   AOI222_X1 i_0_1_291 (.A1(n_0_194), .A2(n_0_1_434), .B1(n_0_210), .B2(
      n_0_1_435), .C1(n_0_341), .C2(n_0_1_433), .ZN(n_0_1_417));
   INV_X1 i_0_1_292 (.A(n_0_1_418), .ZN(n_0_326));
   AOI222_X1 i_0_1_293 (.A1(n_0_195), .A2(n_0_1_434), .B1(n_0_211), .B2(
      n_0_1_435), .C1(n_0_342), .C2(n_0_1_433), .ZN(n_0_1_418));
   INV_X1 i_0_1_294 (.A(n_0_1_419), .ZN(n_0_327));
   AOI222_X1 i_0_1_295 (.A1(n_0_196), .A2(n_0_1_434), .B1(n_0_212), .B2(
      n_0_1_435), .C1(n_0_343), .C2(n_0_1_433), .ZN(n_0_1_419));
   INV_X1 i_0_1_296 (.A(n_0_1_420), .ZN(n_0_328));
   AOI222_X1 i_0_1_297 (.A1(n_0_197), .A2(n_0_1_434), .B1(n_0_213), .B2(
      n_0_1_435), .C1(n_0_344), .C2(n_0_1_433), .ZN(n_0_1_420));
   INV_X1 i_0_1_298 (.A(n_0_1_421), .ZN(n_0_329));
   AOI222_X1 i_0_1_299 (.A1(n_0_198), .A2(n_0_1_434), .B1(n_0_214), .B2(
      n_0_1_435), .C1(n_0_345), .C2(n_0_1_433), .ZN(n_0_1_421));
   INV_X1 i_0_1_300 (.A(n_0_1_422), .ZN(n_0_330));
   AOI222_X1 i_0_1_301 (.A1(n_0_215), .A2(n_0_1_435), .B1(n_0_199), .B2(
      n_0_1_434), .C1(n_0_346), .C2(n_0_1_433), .ZN(n_0_1_422));
   INV_X1 i_0_1_302 (.A(n_0_1_423), .ZN(n_0_331));
   AOI222_X1 i_0_1_303 (.A1(n_0_216), .A2(n_0_1_435), .B1(n_0_200), .B2(
      n_0_1_434), .C1(n_0_347), .C2(n_0_1_433), .ZN(n_0_1_423));
   INV_X1 i_0_1_304 (.A(n_0_1_424), .ZN(n_0_332));
   AOI222_X1 i_0_1_305 (.A1(n_0_217), .A2(n_0_1_435), .B1(n_0_201), .B2(
      n_0_1_434), .C1(n_0_348), .C2(n_0_1_433), .ZN(n_0_1_424));
   INV_X1 i_0_1_306 (.A(n_0_1_425), .ZN(n_0_333));
   AOI222_X1 i_0_1_307 (.A1(n_0_218), .A2(n_0_1_435), .B1(n_0_202), .B2(
      n_0_1_434), .C1(n_0_349), .C2(n_0_1_433), .ZN(n_0_1_425));
   INV_X1 i_0_1_308 (.A(n_0_1_426), .ZN(n_0_334));
   AOI222_X1 i_0_1_309 (.A1(n_0_219), .A2(n_0_1_435), .B1(n_0_203), .B2(
      n_0_1_434), .C1(n_0_350), .C2(n_0_1_433), .ZN(n_0_1_426));
   INV_X1 i_0_1_310 (.A(n_0_1_427), .ZN(n_0_335));
   AOI222_X1 i_0_1_311 (.A1(n_0_220), .A2(n_0_1_435), .B1(n_0_204), .B2(
      n_0_1_434), .C1(n_0_351), .C2(n_0_1_433), .ZN(n_0_1_427));
   INV_X1 i_0_1_312 (.A(n_0_1_428), .ZN(n_0_336));
   AOI222_X1 i_0_1_313 (.A1(n_0_221), .A2(n_0_1_435), .B1(n_0_205), .B2(
      n_0_1_434), .C1(n_0_352), .C2(n_0_1_433), .ZN(n_0_1_428));
   INV_X1 i_0_1_314 (.A(n_0_1_429), .ZN(n_0_337));
   AOI222_X1 i_0_1_315 (.A1(n_0_222), .A2(n_0_1_435), .B1(n_0_206), .B2(
      n_0_1_434), .C1(n_0_353), .C2(n_0_1_433), .ZN(n_0_1_429));
   INV_X1 i_0_1_316 (.A(n_0_1_430), .ZN(n_0_338));
   AOI221_X1 i_0_1_317 (.A(n_0_1_432), .B1(n_0_207), .B2(n_0_1_434), .C1(n_0_223), 
      .C2(n_0_1_435), .ZN(n_0_1_430));
   INV_X1 i_0_1_318 (.A(n_0_1_431), .ZN(n_0_339));
   AOI221_X1 i_0_1_319 (.A(n_0_1_432), .B1(n_0_208), .B2(n_0_1_434), .C1(n_0_224), 
      .C2(n_0_1_435), .ZN(n_0_1_431));
   AND2_X1 i_0_1_320 (.A1(n_0_354), .A2(n_0_1_433), .ZN(n_0_1_432));
   NOR2_X1 i_0_1_321 (.A1(n_0_1_435), .A2(n_0_1_434), .ZN(n_0_1_433));
   NOR2_X1 i_0_1_322 (.A1(in_b[13]), .A2(n_0_1_825), .ZN(n_0_1_434));
   NOR2_X1 i_0_1_323 (.A1(n_0_1_826), .A2(in_b[12]), .ZN(n_0_1_435));
   INV_X1 i_0_1_324 (.A(n_0_1_436), .ZN(n_0_340));
   AOI222_X1 i_0_1_325 (.A1(n_0_162), .A2(n_0_1_453), .B1(n_0_178), .B2(
      n_0_1_454), .C1(n_0_356), .C2(n_0_1_452), .ZN(n_0_1_436));
   INV_X1 i_0_1_326 (.A(n_0_1_437), .ZN(n_0_341));
   AOI222_X1 i_0_1_327 (.A1(n_0_163), .A2(n_0_1_453), .B1(n_0_179), .B2(
      n_0_1_454), .C1(n_0_357), .C2(n_0_1_452), .ZN(n_0_1_437));
   INV_X1 i_0_1_328 (.A(n_0_1_438), .ZN(n_0_342));
   AOI222_X1 i_0_1_329 (.A1(n_0_164), .A2(n_0_1_453), .B1(n_0_180), .B2(
      n_0_1_454), .C1(n_0_358), .C2(n_0_1_452), .ZN(n_0_1_438));
   INV_X1 i_0_1_330 (.A(n_0_1_439), .ZN(n_0_343));
   AOI222_X1 i_0_1_331 (.A1(n_0_165), .A2(n_0_1_453), .B1(n_0_181), .B2(
      n_0_1_454), .C1(n_0_359), .C2(n_0_1_452), .ZN(n_0_1_439));
   INV_X1 i_0_1_332 (.A(n_0_1_440), .ZN(n_0_344));
   AOI222_X1 i_0_1_333 (.A1(n_0_166), .A2(n_0_1_453), .B1(n_0_182), .B2(
      n_0_1_454), .C1(n_0_360), .C2(n_0_1_452), .ZN(n_0_1_440));
   INV_X1 i_0_1_334 (.A(n_0_1_441), .ZN(n_0_345));
   AOI222_X1 i_0_1_335 (.A1(n_0_167), .A2(n_0_1_453), .B1(n_0_183), .B2(
      n_0_1_454), .C1(n_0_361), .C2(n_0_1_452), .ZN(n_0_1_441));
   INV_X1 i_0_1_336 (.A(n_0_1_442), .ZN(n_0_346));
   AOI222_X1 i_0_1_337 (.A1(n_0_168), .A2(n_0_1_453), .B1(n_0_184), .B2(
      n_0_1_454), .C1(n_0_362), .C2(n_0_1_452), .ZN(n_0_1_442));
   INV_X1 i_0_1_338 (.A(n_0_1_443), .ZN(n_0_347));
   AOI222_X1 i_0_1_339 (.A1(n_0_185), .A2(n_0_1_454), .B1(n_0_169), .B2(
      n_0_1_453), .C1(n_0_363), .C2(n_0_1_452), .ZN(n_0_1_443));
   INV_X1 i_0_1_340 (.A(n_0_1_444), .ZN(n_0_348));
   AOI222_X1 i_0_1_341 (.A1(n_0_186), .A2(n_0_1_454), .B1(n_0_170), .B2(
      n_0_1_453), .C1(n_0_364), .C2(n_0_1_452), .ZN(n_0_1_444));
   INV_X1 i_0_1_342 (.A(n_0_1_445), .ZN(n_0_349));
   AOI222_X1 i_0_1_343 (.A1(n_0_187), .A2(n_0_1_454), .B1(n_0_171), .B2(
      n_0_1_453), .C1(n_0_365), .C2(n_0_1_452), .ZN(n_0_1_445));
   INV_X1 i_0_1_344 (.A(n_0_1_446), .ZN(n_0_350));
   AOI222_X1 i_0_1_345 (.A1(n_0_188), .A2(n_0_1_454), .B1(n_0_172), .B2(
      n_0_1_453), .C1(n_0_366), .C2(n_0_1_452), .ZN(n_0_1_446));
   INV_X1 i_0_1_346 (.A(n_0_1_447), .ZN(n_0_351));
   AOI222_X1 i_0_1_347 (.A1(n_0_189), .A2(n_0_1_454), .B1(n_0_173), .B2(
      n_0_1_453), .C1(n_0_367), .C2(n_0_1_452), .ZN(n_0_1_447));
   INV_X1 i_0_1_348 (.A(n_0_1_448), .ZN(n_0_352));
   AOI222_X1 i_0_1_349 (.A1(n_0_190), .A2(n_0_1_454), .B1(n_0_174), .B2(
      n_0_1_453), .C1(n_0_368), .C2(n_0_1_452), .ZN(n_0_1_448));
   INV_X1 i_0_1_350 (.A(n_0_1_449), .ZN(n_0_353));
   AOI221_X1 i_0_1_351 (.A(n_0_1_451), .B1(n_0_175), .B2(n_0_1_453), .C1(n_0_191), 
      .C2(n_0_1_454), .ZN(n_0_1_449));
   INV_X1 i_0_1_352 (.A(n_0_1_450), .ZN(n_0_354));
   AOI221_X1 i_0_1_353 (.A(n_0_1_451), .B1(n_0_176), .B2(n_0_1_453), .C1(n_0_192), 
      .C2(n_0_1_454), .ZN(n_0_1_450));
   AND2_X1 i_0_1_354 (.A1(n_0_369), .A2(n_0_1_452), .ZN(n_0_1_451));
   NOR2_X1 i_0_1_355 (.A1(n_0_1_454), .A2(n_0_1_453), .ZN(n_0_1_452));
   NOR2_X1 i_0_1_356 (.A1(in_b[12]), .A2(n_0_1_824), .ZN(n_0_1_453));
   NOR2_X1 i_0_1_357 (.A1(n_0_1_825), .A2(in_b[11]), .ZN(n_0_1_454));
   INV_X1 i_0_1_358 (.A(n_0_1_455), .ZN(n_0_355));
   AOI222_X1 i_0_1_359 (.A1(n_0_130), .A2(n_0_1_472), .B1(n_0_146), .B2(
      n_0_1_473), .C1(n_0_371), .C2(n_0_1_471), .ZN(n_0_1_455));
   INV_X1 i_0_1_360 (.A(n_0_1_456), .ZN(n_0_356));
   AOI222_X1 i_0_1_361 (.A1(n_0_131), .A2(n_0_1_472), .B1(n_0_147), .B2(
      n_0_1_473), .C1(n_0_372), .C2(n_0_1_471), .ZN(n_0_1_456));
   INV_X1 i_0_1_362 (.A(n_0_1_457), .ZN(n_0_357));
   AOI222_X1 i_0_1_363 (.A1(n_0_132), .A2(n_0_1_472), .B1(n_0_148), .B2(
      n_0_1_473), .C1(n_0_373), .C2(n_0_1_471), .ZN(n_0_1_457));
   INV_X1 i_0_1_364 (.A(n_0_1_458), .ZN(n_0_358));
   AOI222_X1 i_0_1_365 (.A1(n_0_133), .A2(n_0_1_472), .B1(n_0_149), .B2(
      n_0_1_473), .C1(n_0_374), .C2(n_0_1_471), .ZN(n_0_1_458));
   INV_X1 i_0_1_366 (.A(n_0_1_459), .ZN(n_0_359));
   AOI222_X1 i_0_1_367 (.A1(n_0_134), .A2(n_0_1_472), .B1(n_0_150), .B2(
      n_0_1_473), .C1(n_0_375), .C2(n_0_1_471), .ZN(n_0_1_459));
   INV_X1 i_0_1_368 (.A(n_0_1_460), .ZN(n_0_360));
   AOI222_X1 i_0_1_369 (.A1(n_0_135), .A2(n_0_1_472), .B1(n_0_151), .B2(
      n_0_1_473), .C1(n_0_376), .C2(n_0_1_471), .ZN(n_0_1_460));
   INV_X1 i_0_1_370 (.A(n_0_1_461), .ZN(n_0_361));
   AOI222_X1 i_0_1_371 (.A1(n_0_136), .A2(n_0_1_472), .B1(n_0_152), .B2(
      n_0_1_473), .C1(n_0_377), .C2(n_0_1_471), .ZN(n_0_1_461));
   INV_X1 i_0_1_372 (.A(n_0_1_462), .ZN(n_0_362));
   AOI222_X1 i_0_1_373 (.A1(n_0_137), .A2(n_0_1_472), .B1(n_0_153), .B2(
      n_0_1_473), .C1(n_0_378), .C2(n_0_1_471), .ZN(n_0_1_462));
   INV_X1 i_0_1_374 (.A(n_0_1_463), .ZN(n_0_363));
   AOI222_X1 i_0_1_375 (.A1(n_0_138), .A2(n_0_1_472), .B1(n_0_154), .B2(
      n_0_1_473), .C1(n_0_379), .C2(n_0_1_471), .ZN(n_0_1_463));
   INV_X1 i_0_1_376 (.A(n_0_1_464), .ZN(n_0_364));
   AOI222_X1 i_0_1_377 (.A1(n_0_155), .A2(n_0_1_473), .B1(n_0_139), .B2(
      n_0_1_472), .C1(n_0_380), .C2(n_0_1_471), .ZN(n_0_1_464));
   INV_X1 i_0_1_378 (.A(n_0_1_465), .ZN(n_0_365));
   AOI222_X1 i_0_1_379 (.A1(n_0_156), .A2(n_0_1_473), .B1(n_0_140), .B2(
      n_0_1_472), .C1(n_0_381), .C2(n_0_1_471), .ZN(n_0_1_465));
   INV_X1 i_0_1_380 (.A(n_0_1_466), .ZN(n_0_366));
   AOI222_X1 i_0_1_381 (.A1(n_0_157), .A2(n_0_1_473), .B1(n_0_141), .B2(
      n_0_1_472), .C1(n_0_382), .C2(n_0_1_471), .ZN(n_0_1_466));
   INV_X1 i_0_1_382 (.A(n_0_1_467), .ZN(n_0_367));
   AOI222_X1 i_0_1_383 (.A1(n_0_158), .A2(n_0_1_473), .B1(n_0_142), .B2(
      n_0_1_472), .C1(n_0_383), .C2(n_0_1_471), .ZN(n_0_1_467));
   INV_X1 i_0_1_384 (.A(n_0_1_468), .ZN(n_0_368));
   AOI221_X1 i_0_1_385 (.A(n_0_1_470), .B1(n_0_143), .B2(n_0_1_472), .C1(n_0_159), 
      .C2(n_0_1_473), .ZN(n_0_1_468));
   INV_X1 i_0_1_386 (.A(n_0_1_469), .ZN(n_0_369));
   AOI221_X1 i_0_1_387 (.A(n_0_1_470), .B1(n_0_144), .B2(n_0_1_472), .C1(n_0_160), 
      .C2(n_0_1_473), .ZN(n_0_1_469));
   AND2_X1 i_0_1_388 (.A1(n_0_384), .A2(n_0_1_471), .ZN(n_0_1_470));
   NOR2_X1 i_0_1_389 (.A1(n_0_1_473), .A2(n_0_1_472), .ZN(n_0_1_471));
   NOR2_X1 i_0_1_390 (.A1(in_b[11]), .A2(n_0_1_823), .ZN(n_0_1_472));
   NOR2_X1 i_0_1_391 (.A1(n_0_1_824), .A2(in_b[10]), .ZN(n_0_1_473));
   INV_X1 i_0_1_392 (.A(n_0_1_474), .ZN(n_0_370));
   AOI222_X1 i_0_1_393 (.A1(n_0_98), .A2(n_0_1_491), .B1(n_0_114), .B2(n_0_1_492), 
      .C1(n_0_386), .C2(n_0_1_490), .ZN(n_0_1_474));
   INV_X1 i_0_1_394 (.A(n_0_1_475), .ZN(n_0_371));
   AOI222_X1 i_0_1_395 (.A1(n_0_99), .A2(n_0_1_491), .B1(n_0_115), .B2(n_0_1_492), 
      .C1(n_0_387), .C2(n_0_1_490), .ZN(n_0_1_475));
   INV_X1 i_0_1_396 (.A(n_0_1_476), .ZN(n_0_372));
   AOI222_X1 i_0_1_397 (.A1(n_0_100), .A2(n_0_1_491), .B1(n_0_116), .B2(
      n_0_1_492), .C1(n_0_388), .C2(n_0_1_490), .ZN(n_0_1_476));
   INV_X1 i_0_1_398 (.A(n_0_1_477), .ZN(n_0_373));
   AOI222_X1 i_0_1_399 (.A1(n_0_101), .A2(n_0_1_491), .B1(n_0_117), .B2(
      n_0_1_492), .C1(n_0_389), .C2(n_0_1_490), .ZN(n_0_1_477));
   INV_X1 i_0_1_400 (.A(n_0_1_478), .ZN(n_0_374));
   AOI222_X1 i_0_1_401 (.A1(n_0_102), .A2(n_0_1_491), .B1(n_0_118), .B2(
      n_0_1_492), .C1(n_0_390), .C2(n_0_1_490), .ZN(n_0_1_478));
   INV_X1 i_0_1_402 (.A(n_0_1_479), .ZN(n_0_375));
   AOI222_X1 i_0_1_403 (.A1(n_0_103), .A2(n_0_1_491), .B1(n_0_119), .B2(
      n_0_1_492), .C1(n_0_391), .C2(n_0_1_490), .ZN(n_0_1_479));
   INV_X1 i_0_1_404 (.A(n_0_1_480), .ZN(n_0_376));
   AOI222_X1 i_0_1_405 (.A1(n_0_104), .A2(n_0_1_491), .B1(n_0_120), .B2(
      n_0_1_492), .C1(n_0_392), .C2(n_0_1_490), .ZN(n_0_1_480));
   INV_X1 i_0_1_406 (.A(n_0_1_481), .ZN(n_0_377));
   AOI222_X1 i_0_1_407 (.A1(n_0_105), .A2(n_0_1_491), .B1(n_0_121), .B2(
      n_0_1_492), .C1(n_0_393), .C2(n_0_1_490), .ZN(n_0_1_481));
   INV_X1 i_0_1_408 (.A(n_0_1_482), .ZN(n_0_378));
   AOI222_X1 i_0_1_409 (.A1(n_0_106), .A2(n_0_1_491), .B1(n_0_122), .B2(
      n_0_1_492), .C1(n_0_394), .C2(n_0_1_490), .ZN(n_0_1_482));
   INV_X1 i_0_1_410 (.A(n_0_1_483), .ZN(n_0_379));
   AOI222_X1 i_0_1_411 (.A1(n_0_107), .A2(n_0_1_491), .B1(n_0_123), .B2(
      n_0_1_492), .C1(n_0_395), .C2(n_0_1_490), .ZN(n_0_1_483));
   INV_X1 i_0_1_412 (.A(n_0_1_484), .ZN(n_0_380));
   AOI222_X1 i_0_1_413 (.A1(n_0_124), .A2(n_0_1_492), .B1(n_0_108), .B2(
      n_0_1_491), .C1(n_0_396), .C2(n_0_1_490), .ZN(n_0_1_484));
   INV_X1 i_0_1_414 (.A(n_0_1_485), .ZN(n_0_381));
   AOI222_X1 i_0_1_415 (.A1(n_0_125), .A2(n_0_1_492), .B1(n_0_109), .B2(
      n_0_1_491), .C1(n_0_397), .C2(n_0_1_490), .ZN(n_0_1_485));
   INV_X1 i_0_1_416 (.A(n_0_1_486), .ZN(n_0_382));
   AOI222_X1 i_0_1_417 (.A1(n_0_126), .A2(n_0_1_492), .B1(n_0_110), .B2(
      n_0_1_491), .C1(n_0_398), .C2(n_0_1_490), .ZN(n_0_1_486));
   INV_X1 i_0_1_418 (.A(n_0_1_487), .ZN(n_0_383));
   AOI221_X1 i_0_1_419 (.A(n_0_1_489), .B1(n_0_111), .B2(n_0_1_491), .C1(n_0_127), 
      .C2(n_0_1_492), .ZN(n_0_1_487));
   INV_X1 i_0_1_420 (.A(n_0_1_488), .ZN(n_0_384));
   AOI221_X1 i_0_1_421 (.A(n_0_1_489), .B1(n_0_112), .B2(n_0_1_491), .C1(n_0_128), 
      .C2(n_0_1_492), .ZN(n_0_1_488));
   AND2_X1 i_0_1_422 (.A1(n_0_399), .A2(n_0_1_490), .ZN(n_0_1_489));
   NOR2_X1 i_0_1_423 (.A1(n_0_1_492), .A2(n_0_1_491), .ZN(n_0_1_490));
   NOR2_X1 i_0_1_424 (.A1(in_b[10]), .A2(n_0_1_822), .ZN(n_0_1_491));
   NOR2_X1 i_0_1_425 (.A1(n_0_1_823), .A2(in_b[9]), .ZN(n_0_1_492));
   INV_X1 i_0_1_426 (.A(n_0_1_493), .ZN(n_0_385));
   AOI222_X1 i_0_1_427 (.A1(n_0_66), .A2(n_0_1_510), .B1(n_0_82), .B2(n_0_1_511), 
      .C1(n_0_401), .C2(n_0_1_509), .ZN(n_0_1_493));
   INV_X1 i_0_1_428 (.A(n_0_1_494), .ZN(n_0_386));
   AOI222_X1 i_0_1_429 (.A1(n_0_67), .A2(n_0_1_510), .B1(n_0_83), .B2(n_0_1_511), 
      .C1(n_0_402), .C2(n_0_1_509), .ZN(n_0_1_494));
   INV_X1 i_0_1_430 (.A(n_0_1_495), .ZN(n_0_387));
   AOI222_X1 i_0_1_431 (.A1(n_0_68), .A2(n_0_1_510), .B1(n_0_84), .B2(n_0_1_511), 
      .C1(n_0_403), .C2(n_0_1_509), .ZN(n_0_1_495));
   INV_X1 i_0_1_432 (.A(n_0_1_496), .ZN(n_0_388));
   AOI222_X1 i_0_1_433 (.A1(n_0_69), .A2(n_0_1_510), .B1(n_0_85), .B2(n_0_1_511), 
      .C1(n_0_404), .C2(n_0_1_509), .ZN(n_0_1_496));
   INV_X1 i_0_1_434 (.A(n_0_1_497), .ZN(n_0_389));
   AOI222_X1 i_0_1_435 (.A1(n_0_70), .A2(n_0_1_510), .B1(n_0_86), .B2(n_0_1_511), 
      .C1(n_0_405), .C2(n_0_1_509), .ZN(n_0_1_497));
   INV_X1 i_0_1_436 (.A(n_0_1_498), .ZN(n_0_390));
   AOI222_X1 i_0_1_437 (.A1(n_0_71), .A2(n_0_1_510), .B1(n_0_87), .B2(n_0_1_511), 
      .C1(n_0_406), .C2(n_0_1_509), .ZN(n_0_1_498));
   INV_X1 i_0_1_438 (.A(n_0_1_499), .ZN(n_0_391));
   AOI222_X1 i_0_1_439 (.A1(n_0_72), .A2(n_0_1_510), .B1(n_0_88), .B2(n_0_1_511), 
      .C1(n_0_407), .C2(n_0_1_509), .ZN(n_0_1_499));
   INV_X1 i_0_1_440 (.A(n_0_1_500), .ZN(n_0_392));
   AOI222_X1 i_0_1_441 (.A1(n_0_73), .A2(n_0_1_510), .B1(n_0_89), .B2(n_0_1_511), 
      .C1(n_0_408), .C2(n_0_1_509), .ZN(n_0_1_500));
   INV_X1 i_0_1_442 (.A(n_0_1_501), .ZN(n_0_393));
   AOI222_X1 i_0_1_443 (.A1(n_0_74), .A2(n_0_1_510), .B1(n_0_90), .B2(n_0_1_511), 
      .C1(n_0_409), .C2(n_0_1_509), .ZN(n_0_1_501));
   INV_X1 i_0_1_444 (.A(n_0_1_502), .ZN(n_0_394));
   AOI222_X1 i_0_1_445 (.A1(n_0_75), .A2(n_0_1_510), .B1(n_0_91), .B2(n_0_1_511), 
      .C1(n_0_410), .C2(n_0_1_509), .ZN(n_0_1_502));
   INV_X1 i_0_1_446 (.A(n_0_1_503), .ZN(n_0_395));
   AOI222_X1 i_0_1_447 (.A1(n_0_76), .A2(n_0_1_510), .B1(n_0_92), .B2(n_0_1_511), 
      .C1(n_0_411), .C2(n_0_1_509), .ZN(n_0_1_503));
   INV_X1 i_0_1_448 (.A(n_0_1_504), .ZN(n_0_396));
   AOI222_X1 i_0_1_449 (.A1(n_0_77), .A2(n_0_1_510), .B1(n_0_93), .B2(n_0_1_511), 
      .C1(n_0_412), .C2(n_0_1_509), .ZN(n_0_1_504));
   INV_X1 i_0_1_450 (.A(n_0_1_505), .ZN(n_0_397));
   AOI222_X1 i_0_1_451 (.A1(n_0_94), .A2(n_0_1_511), .B1(n_0_78), .B2(n_0_1_510), 
      .C1(n_0_413), .C2(n_0_1_509), .ZN(n_0_1_505));
   INV_X1 i_0_1_452 (.A(n_0_1_506), .ZN(n_0_398));
   AOI221_X1 i_0_1_453 (.A(n_0_1_508), .B1(n_0_79), .B2(n_0_1_510), .C1(n_0_95), 
      .C2(n_0_1_511), .ZN(n_0_1_506));
   INV_X1 i_0_1_454 (.A(n_0_1_507), .ZN(n_0_399));
   AOI221_X1 i_0_1_455 (.A(n_0_1_508), .B1(n_0_80), .B2(n_0_1_510), .C1(n_0_96), 
      .C2(n_0_1_511), .ZN(n_0_1_507));
   AND2_X1 i_0_1_456 (.A1(n_0_414), .A2(n_0_1_509), .ZN(n_0_1_508));
   NOR2_X1 i_0_1_457 (.A1(n_0_1_511), .A2(n_0_1_510), .ZN(n_0_1_509));
   NOR2_X1 i_0_1_458 (.A1(in_b[9]), .A2(n_0_1_821), .ZN(n_0_1_510));
   NOR2_X1 i_0_1_459 (.A1(n_0_1_822), .A2(in_b[8]), .ZN(n_0_1_511));
   INV_X1 i_0_1_460 (.A(n_0_1_512), .ZN(n_0_400));
   AOI222_X1 i_0_1_461 (.A1(n_0_34), .A2(n_0_1_529), .B1(n_0_50), .B2(n_0_1_530), 
      .C1(n_0_416), .C2(n_0_1_528), .ZN(n_0_1_512));
   INV_X1 i_0_1_462 (.A(n_0_1_513), .ZN(n_0_401));
   AOI222_X1 i_0_1_463 (.A1(n_0_35), .A2(n_0_1_529), .B1(n_0_51), .B2(n_0_1_530), 
      .C1(n_0_417), .C2(n_0_1_528), .ZN(n_0_1_513));
   INV_X1 i_0_1_464 (.A(n_0_1_514), .ZN(n_0_402));
   AOI222_X1 i_0_1_465 (.A1(n_0_36), .A2(n_0_1_529), .B1(n_0_52), .B2(n_0_1_530), 
      .C1(n_0_418), .C2(n_0_1_528), .ZN(n_0_1_514));
   INV_X1 i_0_1_466 (.A(n_0_1_515), .ZN(n_0_403));
   AOI222_X1 i_0_1_467 (.A1(n_0_37), .A2(n_0_1_529), .B1(n_0_53), .B2(n_0_1_530), 
      .C1(n_0_419), .C2(n_0_1_528), .ZN(n_0_1_515));
   INV_X1 i_0_1_468 (.A(n_0_1_516), .ZN(n_0_404));
   AOI222_X1 i_0_1_469 (.A1(n_0_38), .A2(n_0_1_529), .B1(n_0_54), .B2(n_0_1_530), 
      .C1(n_0_420), .C2(n_0_1_528), .ZN(n_0_1_516));
   INV_X1 i_0_1_470 (.A(n_0_1_517), .ZN(n_0_405));
   AOI222_X1 i_0_1_471 (.A1(n_0_39), .A2(n_0_1_529), .B1(n_0_55), .B2(n_0_1_530), 
      .C1(n_0_421), .C2(n_0_1_528), .ZN(n_0_1_517));
   INV_X1 i_0_1_472 (.A(n_0_1_518), .ZN(n_0_406));
   AOI222_X1 i_0_1_473 (.A1(n_0_40), .A2(n_0_1_529), .B1(n_0_56), .B2(n_0_1_530), 
      .C1(n_0_422), .C2(n_0_1_528), .ZN(n_0_1_518));
   INV_X1 i_0_1_474 (.A(n_0_1_519), .ZN(n_0_407));
   AOI222_X1 i_0_1_475 (.A1(n_0_41), .A2(n_0_1_529), .B1(n_0_57), .B2(n_0_1_530), 
      .C1(n_0_423), .C2(n_0_1_528), .ZN(n_0_1_519));
   INV_X1 i_0_1_476 (.A(n_0_1_520), .ZN(n_0_408));
   AOI222_X1 i_0_1_477 (.A1(n_0_42), .A2(n_0_1_529), .B1(n_0_58), .B2(n_0_1_530), 
      .C1(n_0_424), .C2(n_0_1_528), .ZN(n_0_1_520));
   INV_X1 i_0_1_478 (.A(n_0_1_521), .ZN(n_0_409));
   AOI222_X1 i_0_1_479 (.A1(n_0_43), .A2(n_0_1_529), .B1(n_0_59), .B2(n_0_1_530), 
      .C1(n_0_425), .C2(n_0_1_528), .ZN(n_0_1_521));
   INV_X1 i_0_1_480 (.A(n_0_1_522), .ZN(n_0_410));
   AOI222_X1 i_0_1_481 (.A1(n_0_44), .A2(n_0_1_529), .B1(n_0_60), .B2(n_0_1_530), 
      .C1(n_0_426), .C2(n_0_1_528), .ZN(n_0_1_522));
   INV_X1 i_0_1_482 (.A(n_0_1_523), .ZN(n_0_411));
   AOI222_X1 i_0_1_483 (.A1(n_0_45), .A2(n_0_1_529), .B1(n_0_61), .B2(n_0_1_530), 
      .C1(n_0_427), .C2(n_0_1_528), .ZN(n_0_1_523));
   INV_X1 i_0_1_484 (.A(n_0_1_524), .ZN(n_0_412));
   AOI222_X1 i_0_1_485 (.A1(n_0_46), .A2(n_0_1_529), .B1(n_0_62), .B2(n_0_1_530), 
      .C1(n_0_428), .C2(n_0_1_528), .ZN(n_0_1_524));
   INV_X1 i_0_1_486 (.A(n_0_1_525), .ZN(n_0_413));
   AOI221_X1 i_0_1_487 (.A(n_0_1_527), .B1(n_0_47), .B2(n_0_1_529), .C1(n_0_63), 
      .C2(n_0_1_530), .ZN(n_0_1_525));
   INV_X1 i_0_1_488 (.A(n_0_1_526), .ZN(n_0_414));
   AOI221_X1 i_0_1_489 (.A(n_0_1_527), .B1(n_0_48), .B2(n_0_1_529), .C1(n_0_64), 
      .C2(n_0_1_530), .ZN(n_0_1_526));
   AND2_X1 i_0_1_490 (.A1(n_0_429), .A2(n_0_1_528), .ZN(n_0_1_527));
   NOR2_X1 i_0_1_491 (.A1(n_0_1_530), .A2(n_0_1_529), .ZN(n_0_1_528));
   NOR2_X1 i_0_1_492 (.A1(in_b[8]), .A2(n_0_1_820), .ZN(n_0_1_529));
   NOR2_X1 i_0_1_493 (.A1(n_0_1_821), .A2(in_b[7]), .ZN(n_0_1_530));
   INV_X1 i_0_1_494 (.A(n_0_1_531), .ZN(n_0_415));
   AOI222_X1 i_0_1_495 (.A1(n_0_1), .A2(n_0_1_548), .B1(n_0_18), .B2(n_0_1_549), 
      .C1(n_0_431), .C2(n_0_1_547), .ZN(n_0_1_531));
   INV_X1 i_0_1_496 (.A(n_0_1_532), .ZN(n_0_416));
   AOI222_X1 i_0_1_497 (.A1(n_0_2), .A2(n_0_1_548), .B1(n_0_19), .B2(n_0_1_549), 
      .C1(n_0_432), .C2(n_0_1_547), .ZN(n_0_1_532));
   INV_X1 i_0_1_498 (.A(n_0_1_533), .ZN(n_0_417));
   AOI222_X1 i_0_1_499 (.A1(n_0_3), .A2(n_0_1_548), .B1(n_0_20), .B2(n_0_1_549), 
      .C1(n_0_433), .C2(n_0_1_547), .ZN(n_0_1_533));
   INV_X1 i_0_1_500 (.A(n_0_1_534), .ZN(n_0_418));
   AOI222_X1 i_0_1_501 (.A1(n_0_5), .A2(n_0_1_548), .B1(n_0_21), .B2(n_0_1_549), 
      .C1(n_0_434), .C2(n_0_1_547), .ZN(n_0_1_534));
   INV_X1 i_0_1_502 (.A(n_0_1_535), .ZN(n_0_419));
   AOI222_X1 i_0_1_503 (.A1(n_0_6), .A2(n_0_1_548), .B1(n_0_22), .B2(n_0_1_549), 
      .C1(n_0_435), .C2(n_0_1_547), .ZN(n_0_1_535));
   INV_X1 i_0_1_504 (.A(n_0_1_536), .ZN(n_0_420));
   AOI222_X1 i_0_1_505 (.A1(n_0_7), .A2(n_0_1_548), .B1(n_0_23), .B2(n_0_1_549), 
      .C1(n_0_436), .C2(n_0_1_547), .ZN(n_0_1_536));
   INV_X1 i_0_1_506 (.A(n_0_1_537), .ZN(n_0_421));
   AOI222_X1 i_0_1_507 (.A1(n_0_8), .A2(n_0_1_548), .B1(n_0_24), .B2(n_0_1_549), 
      .C1(n_0_437), .C2(n_0_1_547), .ZN(n_0_1_537));
   INV_X1 i_0_1_508 (.A(n_0_1_538), .ZN(n_0_422));
   AOI222_X1 i_0_1_509 (.A1(n_0_9), .A2(n_0_1_548), .B1(n_0_25), .B2(n_0_1_549), 
      .C1(n_0_438), .C2(n_0_1_547), .ZN(n_0_1_538));
   INV_X1 i_0_1_510 (.A(n_0_1_539), .ZN(n_0_423));
   AOI222_X1 i_0_1_511 (.A1(n_0_10), .A2(n_0_1_548), .B1(n_0_26), .B2(n_0_1_549), 
      .C1(n_0_439), .C2(n_0_1_547), .ZN(n_0_1_539));
   INV_X1 i_0_1_512 (.A(n_0_1_540), .ZN(n_0_424));
   AOI222_X1 i_0_1_513 (.A1(n_0_11), .A2(n_0_1_548), .B1(n_0_27), .B2(n_0_1_549), 
      .C1(n_0_440), .C2(n_0_1_547), .ZN(n_0_1_540));
   INV_X1 i_0_1_514 (.A(n_0_1_541), .ZN(n_0_425));
   AOI222_X1 i_0_1_515 (.A1(n_0_12), .A2(n_0_1_548), .B1(n_0_28), .B2(n_0_1_549), 
      .C1(n_0_441), .C2(n_0_1_547), .ZN(n_0_1_541));
   INV_X1 i_0_1_516 (.A(n_0_1_542), .ZN(n_0_426));
   AOI222_X1 i_0_1_517 (.A1(n_0_13), .A2(n_0_1_548), .B1(n_0_29), .B2(n_0_1_549), 
      .C1(n_0_442), .C2(n_0_1_547), .ZN(n_0_1_542));
   INV_X1 i_0_1_518 (.A(n_0_1_543), .ZN(n_0_427));
   AOI222_X1 i_0_1_519 (.A1(n_0_14), .A2(n_0_1_548), .B1(n_0_30), .B2(n_0_1_549), 
      .C1(n_0_443), .C2(n_0_1_547), .ZN(n_0_1_543));
   INV_X1 i_0_1_520 (.A(n_0_1_544), .ZN(n_0_428));
   AOI221_X1 i_0_1_521 (.A(n_0_1_546), .B1(n_0_15), .B2(n_0_1_548), .C1(n_0_31), 
      .C2(n_0_1_549), .ZN(n_0_1_544));
   INV_X1 i_0_1_522 (.A(n_0_1_545), .ZN(n_0_429));
   AOI221_X1 i_0_1_523 (.A(n_0_1_546), .B1(n_0_16), .B2(n_0_1_548), .C1(n_0_32), 
      .C2(n_0_1_549), .ZN(n_0_1_545));
   AND2_X1 i_0_1_524 (.A1(n_0_444), .A2(n_0_1_547), .ZN(n_0_1_546));
   NOR2_X1 i_0_1_525 (.A1(n_0_1_549), .A2(n_0_1_548), .ZN(n_0_1_547));
   NOR2_X1 i_0_1_526 (.A1(in_b[7]), .A2(n_0_1_819), .ZN(n_0_1_548));
   NOR2_X1 i_0_1_527 (.A1(n_0_1_820), .A2(in_b[6]), .ZN(n_0_1_549));
   INV_X1 i_0_1_528 (.A(n_0_1_550), .ZN(n_0_430));
   AOI222_X1 i_0_1_529 (.A1(n_0_1_298), .A2(n_0_1_705), .B1(n_0_1_311), .B2(
      n_0_1_707), .C1(n_0_1_704), .C2(n_0_1_551), .ZN(n_0_1_550));
   INV_X1 i_0_1_530 (.A(n_0_1_552), .ZN(n_0_1_551));
   AOI222_X1 i_0_1_531 (.A1(n_0_1_273), .A2(n_0_1_717), .B1(n_0_1_286), .B2(
      n_0_1_719), .C1(n_0_1_716), .C2(n_0_1_553), .ZN(n_0_1_552));
   INV_X1 i_0_1_532 (.A(n_0_1_554), .ZN(n_0_1_553));
   AOI222_X1 i_0_1_533 (.A1(n_0_1_248), .A2(n_0_1_730), .B1(n_0_1_261), .B2(
      n_0_1_728), .C1(n_0_1_727), .C2(n_0_1_555), .ZN(n_0_1_554));
   INV_X1 i_0_1_534 (.A(n_0_1_556), .ZN(n_0_1_555));
   AOI222_X1 i_0_1_535 (.A1(n_0_1_223), .A2(n_0_1_739), .B1(n_0_1_236), .B2(
      n_0_1_741), .C1(n_0_1_738), .C2(n_0_1_557), .ZN(n_0_1_556));
   INV_X1 i_0_1_536 (.A(n_0_1_558), .ZN(n_0_1_557));
   AOI222_X1 i_0_1_537 (.A1(n_0_1_198), .A2(n_0_1_751), .B1(n_0_1_211), .B2(
      n_0_1_753), .C1(n_0_1_750), .C2(n_0_1_559), .ZN(n_0_1_558));
   INV_X1 i_0_1_538 (.A(n_0_1_560), .ZN(n_0_1_559));
   AOI222_X1 i_0_1_539 (.A1(n_0_1_173), .A2(n_0_1_763), .B1(n_0_1_186), .B2(
      n_0_1_765), .C1(n_0_1_762), .C2(n_0_1_561), .ZN(n_0_1_560));
   AND2_X1 i_0_1_540 (.A1(in_b[0]), .A2(n_0_451), .ZN(n_0_1_561));
   INV_X1 i_0_1_541 (.A(n_0_1_562), .ZN(n_0_431));
   AOI222_X1 i_0_1_542 (.A1(n_0_1_299), .A2(n_0_1_705), .B1(n_0_1_312), .B2(
      n_0_1_707), .C1(n_0_1_704), .C2(n_0_1_563), .ZN(n_0_1_562));
   INV_X1 i_0_1_543 (.A(n_0_1_564), .ZN(n_0_1_563));
   AOI222_X1 i_0_1_544 (.A1(n_0_1_274), .A2(n_0_1_717), .B1(n_0_1_287), .B2(
      n_0_1_719), .C1(n_0_1_716), .C2(n_0_1_565), .ZN(n_0_1_564));
   INV_X1 i_0_1_545 (.A(n_0_1_566), .ZN(n_0_1_565));
   AOI222_X1 i_0_1_546 (.A1(n_0_1_249), .A2(n_0_1_730), .B1(n_0_1_262), .B2(
      n_0_1_728), .C1(n_0_1_727), .C2(n_0_1_567), .ZN(n_0_1_566));
   INV_X1 i_0_1_547 (.A(n_0_1_568), .ZN(n_0_1_567));
   AOI222_X1 i_0_1_548 (.A1(n_0_1_224), .A2(n_0_1_739), .B1(n_0_1_237), .B2(
      n_0_1_741), .C1(n_0_1_738), .C2(n_0_1_569), .ZN(n_0_1_568));
   INV_X1 i_0_1_549 (.A(n_0_1_570), .ZN(n_0_1_569));
   AOI222_X1 i_0_1_550 (.A1(n_0_1_199), .A2(n_0_1_751), .B1(n_0_1_212), .B2(
      n_0_1_753), .C1(n_0_1_750), .C2(n_0_1_571), .ZN(n_0_1_570));
   INV_X1 i_0_1_551 (.A(n_0_1_572), .ZN(n_0_1_571));
   AOI222_X1 i_0_1_552 (.A1(n_0_1_174), .A2(n_0_1_763), .B1(n_0_1_187), .B2(
      n_0_1_765), .C1(n_0_1_762), .C2(n_0_1_573), .ZN(n_0_1_572));
   AND2_X1 i_0_1_553 (.A1(in_b[0]), .A2(n_0_452), .ZN(n_0_1_573));
   INV_X1 i_0_1_554 (.A(n_0_1_574), .ZN(n_0_432));
   AOI222_X1 i_0_1_555 (.A1(n_0_1_300), .A2(n_0_1_705), .B1(n_0_1_313), .B2(
      n_0_1_707), .C1(n_0_1_704), .C2(n_0_1_575), .ZN(n_0_1_574));
   INV_X1 i_0_1_556 (.A(n_0_1_576), .ZN(n_0_1_575));
   AOI222_X1 i_0_1_557 (.A1(n_0_1_275), .A2(n_0_1_717), .B1(n_0_1_288), .B2(
      n_0_1_719), .C1(n_0_1_716), .C2(n_0_1_577), .ZN(n_0_1_576));
   INV_X1 i_0_1_558 (.A(n_0_1_578), .ZN(n_0_1_577));
   AOI222_X1 i_0_1_559 (.A1(n_0_1_250), .A2(n_0_1_730), .B1(n_0_1_263), .B2(
      n_0_1_728), .C1(n_0_1_727), .C2(n_0_1_579), .ZN(n_0_1_578));
   INV_X1 i_0_1_560 (.A(n_0_1_580), .ZN(n_0_1_579));
   AOI222_X1 i_0_1_561 (.A1(n_0_1_225), .A2(n_0_1_739), .B1(n_0_1_238), .B2(
      n_0_1_741), .C1(n_0_1_738), .C2(n_0_1_581), .ZN(n_0_1_580));
   INV_X1 i_0_1_562 (.A(n_0_1_582), .ZN(n_0_1_581));
   AOI222_X1 i_0_1_563 (.A1(n_0_1_200), .A2(n_0_1_751), .B1(n_0_1_213), .B2(
      n_0_1_753), .C1(n_0_1_750), .C2(n_0_1_583), .ZN(n_0_1_582));
   INV_X1 i_0_1_564 (.A(n_0_1_584), .ZN(n_0_1_583));
   AOI222_X1 i_0_1_565 (.A1(n_0_1_175), .A2(n_0_1_763), .B1(n_0_1_188), .B2(
      n_0_1_765), .C1(n_0_1_762), .C2(n_0_1_585), .ZN(n_0_1_584));
   AND2_X1 i_0_1_566 (.A1(in_b[0]), .A2(n_0_453), .ZN(n_0_1_585));
   INV_X1 i_0_1_567 (.A(n_0_1_586), .ZN(n_0_433));
   AOI222_X1 i_0_1_568 (.A1(n_0_1_301), .A2(n_0_1_705), .B1(n_0_1_314), .B2(
      n_0_1_707), .C1(n_0_1_704), .C2(n_0_1_587), .ZN(n_0_1_586));
   INV_X1 i_0_1_569 (.A(n_0_1_588), .ZN(n_0_1_587));
   AOI222_X1 i_0_1_570 (.A1(n_0_1_276), .A2(n_0_1_717), .B1(n_0_1_289), .B2(
      n_0_1_719), .C1(n_0_1_716), .C2(n_0_1_589), .ZN(n_0_1_588));
   INV_X1 i_0_1_571 (.A(n_0_1_590), .ZN(n_0_1_589));
   AOI222_X1 i_0_1_572 (.A1(n_0_1_251), .A2(n_0_1_730), .B1(n_0_1_264), .B2(
      n_0_1_728), .C1(n_0_1_727), .C2(n_0_1_591), .ZN(n_0_1_590));
   INV_X1 i_0_1_573 (.A(n_0_1_592), .ZN(n_0_1_591));
   AOI222_X1 i_0_1_574 (.A1(n_0_1_226), .A2(n_0_1_739), .B1(n_0_1_239), .B2(
      n_0_1_741), .C1(n_0_1_738), .C2(n_0_1_593), .ZN(n_0_1_592));
   INV_X1 i_0_1_575 (.A(n_0_1_594), .ZN(n_0_1_593));
   AOI222_X1 i_0_1_576 (.A1(n_0_1_201), .A2(n_0_1_751), .B1(n_0_1_214), .B2(
      n_0_1_753), .C1(n_0_1_750), .C2(n_0_1_595), .ZN(n_0_1_594));
   INV_X1 i_0_1_577 (.A(n_0_1_596), .ZN(n_0_1_595));
   AOI222_X1 i_0_1_578 (.A1(n_0_1_176), .A2(n_0_1_763), .B1(n_0_1_189), .B2(
      n_0_1_765), .C1(n_0_1_762), .C2(n_0_1_597), .ZN(n_0_1_596));
   AND2_X1 i_0_1_579 (.A1(in_b[0]), .A2(n_0_454), .ZN(n_0_1_597));
   INV_X1 i_0_1_580 (.A(n_0_1_598), .ZN(n_0_434));
   AOI222_X1 i_0_1_581 (.A1(n_0_1_302), .A2(n_0_1_705), .B1(n_0_1_315), .B2(
      n_0_1_707), .C1(n_0_1_704), .C2(n_0_1_599), .ZN(n_0_1_598));
   INV_X1 i_0_1_582 (.A(n_0_1_600), .ZN(n_0_1_599));
   AOI222_X1 i_0_1_583 (.A1(n_0_1_277), .A2(n_0_1_717), .B1(n_0_1_290), .B2(
      n_0_1_719), .C1(n_0_1_716), .C2(n_0_1_601), .ZN(n_0_1_600));
   INV_X1 i_0_1_584 (.A(n_0_1_602), .ZN(n_0_1_601));
   AOI222_X1 i_0_1_585 (.A1(n_0_1_252), .A2(n_0_1_730), .B1(n_0_1_265), .B2(
      n_0_1_728), .C1(n_0_1_727), .C2(n_0_1_603), .ZN(n_0_1_602));
   INV_X1 i_0_1_586 (.A(n_0_1_604), .ZN(n_0_1_603));
   AOI222_X1 i_0_1_587 (.A1(n_0_1_227), .A2(n_0_1_739), .B1(n_0_1_240), .B2(
      n_0_1_741), .C1(n_0_1_738), .C2(n_0_1_605), .ZN(n_0_1_604));
   INV_X1 i_0_1_588 (.A(n_0_1_606), .ZN(n_0_1_605));
   AOI222_X1 i_0_1_589 (.A1(n_0_1_202), .A2(n_0_1_751), .B1(n_0_1_215), .B2(
      n_0_1_753), .C1(n_0_1_750), .C2(n_0_1_607), .ZN(n_0_1_606));
   INV_X1 i_0_1_590 (.A(n_0_1_608), .ZN(n_0_1_607));
   AOI222_X1 i_0_1_591 (.A1(n_0_1_177), .A2(n_0_1_763), .B1(n_0_1_190), .B2(
      n_0_1_765), .C1(n_0_1_762), .C2(n_0_1_609), .ZN(n_0_1_608));
   AND2_X1 i_0_1_592 (.A1(in_b[0]), .A2(n_0_455), .ZN(n_0_1_609));
   INV_X1 i_0_1_593 (.A(n_0_1_610), .ZN(n_0_435));
   AOI222_X1 i_0_1_594 (.A1(n_0_1_303), .A2(n_0_1_705), .B1(n_0_1_316), .B2(
      n_0_1_707), .C1(n_0_1_704), .C2(n_0_1_611), .ZN(n_0_1_610));
   INV_X1 i_0_1_595 (.A(n_0_1_612), .ZN(n_0_1_611));
   AOI222_X1 i_0_1_596 (.A1(n_0_1_278), .A2(n_0_1_717), .B1(n_0_1_291), .B2(
      n_0_1_719), .C1(n_0_1_716), .C2(n_0_1_613), .ZN(n_0_1_612));
   INV_X1 i_0_1_597 (.A(n_0_1_614), .ZN(n_0_1_613));
   AOI222_X1 i_0_1_598 (.A1(n_0_1_253), .A2(n_0_1_730), .B1(n_0_1_266), .B2(
      n_0_1_728), .C1(n_0_1_727), .C2(n_0_1_615), .ZN(n_0_1_614));
   INV_X1 i_0_1_599 (.A(n_0_1_616), .ZN(n_0_1_615));
   AOI222_X1 i_0_1_600 (.A1(n_0_1_228), .A2(n_0_1_739), .B1(n_0_1_241), .B2(
      n_0_1_741), .C1(n_0_1_738), .C2(n_0_1_617), .ZN(n_0_1_616));
   INV_X1 i_0_1_601 (.A(n_0_1_618), .ZN(n_0_1_617));
   AOI222_X1 i_0_1_602 (.A1(n_0_1_203), .A2(n_0_1_751), .B1(n_0_1_216), .B2(
      n_0_1_753), .C1(n_0_1_750), .C2(n_0_1_619), .ZN(n_0_1_618));
   INV_X1 i_0_1_603 (.A(n_0_1_620), .ZN(n_0_1_619));
   AOI222_X1 i_0_1_604 (.A1(n_0_1_178), .A2(n_0_1_763), .B1(n_0_1_191), .B2(
      n_0_1_765), .C1(n_0_1_762), .C2(n_0_1_621), .ZN(n_0_1_620));
   AND2_X1 i_0_1_605 (.A1(in_b[0]), .A2(n_0_456), .ZN(n_0_1_621));
   INV_X1 i_0_1_606 (.A(n_0_1_622), .ZN(n_0_436));
   AOI222_X1 i_0_1_607 (.A1(n_0_1_304), .A2(n_0_1_705), .B1(n_0_1_317), .B2(
      n_0_1_707), .C1(n_0_1_704), .C2(n_0_1_623), .ZN(n_0_1_622));
   INV_X1 i_0_1_608 (.A(n_0_1_624), .ZN(n_0_1_623));
   AOI222_X1 i_0_1_609 (.A1(n_0_1_279), .A2(n_0_1_717), .B1(n_0_1_292), .B2(
      n_0_1_719), .C1(n_0_1_716), .C2(n_0_1_625), .ZN(n_0_1_624));
   INV_X1 i_0_1_610 (.A(n_0_1_626), .ZN(n_0_1_625));
   AOI222_X1 i_0_1_611 (.A1(n_0_1_254), .A2(n_0_1_730), .B1(n_0_1_267), .B2(
      n_0_1_728), .C1(n_0_1_727), .C2(n_0_1_627), .ZN(n_0_1_626));
   INV_X1 i_0_1_612 (.A(n_0_1_628), .ZN(n_0_1_627));
   AOI222_X1 i_0_1_613 (.A1(n_0_1_229), .A2(n_0_1_739), .B1(n_0_1_242), .B2(
      n_0_1_741), .C1(n_0_1_738), .C2(n_0_1_629), .ZN(n_0_1_628));
   INV_X1 i_0_1_614 (.A(n_0_1_630), .ZN(n_0_1_629));
   AOI222_X1 i_0_1_615 (.A1(n_0_1_204), .A2(n_0_1_751), .B1(n_0_1_217), .B2(
      n_0_1_753), .C1(n_0_1_750), .C2(n_0_1_631), .ZN(n_0_1_630));
   INV_X1 i_0_1_616 (.A(n_0_1_632), .ZN(n_0_1_631));
   AOI222_X1 i_0_1_617 (.A1(n_0_1_179), .A2(n_0_1_763), .B1(n_0_1_192), .B2(
      n_0_1_765), .C1(n_0_1_762), .C2(n_0_1_633), .ZN(n_0_1_632));
   AND2_X1 i_0_1_618 (.A1(in_b[0]), .A2(n_0_457), .ZN(n_0_1_633));
   INV_X1 i_0_1_619 (.A(n_0_1_634), .ZN(n_0_437));
   AOI222_X1 i_0_1_620 (.A1(n_0_1_305), .A2(n_0_1_705), .B1(n_0_1_318), .B2(
      n_0_1_707), .C1(n_0_1_704), .C2(n_0_1_635), .ZN(n_0_1_634));
   INV_X1 i_0_1_621 (.A(n_0_1_636), .ZN(n_0_1_635));
   AOI222_X1 i_0_1_622 (.A1(n_0_1_280), .A2(n_0_1_717), .B1(n_0_1_293), .B2(
      n_0_1_719), .C1(n_0_1_716), .C2(n_0_1_637), .ZN(n_0_1_636));
   INV_X1 i_0_1_623 (.A(n_0_1_638), .ZN(n_0_1_637));
   AOI222_X1 i_0_1_624 (.A1(n_0_1_255), .A2(n_0_1_730), .B1(n_0_1_268), .B2(
      n_0_1_728), .C1(n_0_1_727), .C2(n_0_1_639), .ZN(n_0_1_638));
   INV_X1 i_0_1_625 (.A(n_0_1_640), .ZN(n_0_1_639));
   AOI222_X1 i_0_1_626 (.A1(n_0_1_230), .A2(n_0_1_739), .B1(n_0_1_243), .B2(
      n_0_1_741), .C1(n_0_1_738), .C2(n_0_1_641), .ZN(n_0_1_640));
   INV_X1 i_0_1_627 (.A(n_0_1_642), .ZN(n_0_1_641));
   AOI222_X1 i_0_1_628 (.A1(n_0_1_205), .A2(n_0_1_751), .B1(n_0_1_218), .B2(
      n_0_1_753), .C1(n_0_1_750), .C2(n_0_1_643), .ZN(n_0_1_642));
   INV_X1 i_0_1_629 (.A(n_0_1_644), .ZN(n_0_1_643));
   AOI222_X1 i_0_1_630 (.A1(n_0_1_180), .A2(n_0_1_763), .B1(n_0_1_193), .B2(
      n_0_1_765), .C1(n_0_1_769), .C2(n_0_1_762), .ZN(n_0_1_644));
   INV_X1 i_0_1_631 (.A(n_0_1_645), .ZN(n_0_438));
   AOI222_X1 i_0_1_632 (.A1(n_0_1_306), .A2(n_0_1_705), .B1(n_0_1_319), .B2(
      n_0_1_707), .C1(n_0_1_704), .C2(n_0_1_646), .ZN(n_0_1_645));
   INV_X1 i_0_1_633 (.A(n_0_1_647), .ZN(n_0_1_646));
   AOI222_X1 i_0_1_634 (.A1(n_0_1_281), .A2(n_0_1_717), .B1(n_0_1_294), .B2(
      n_0_1_719), .C1(n_0_1_716), .C2(n_0_1_648), .ZN(n_0_1_647));
   INV_X1 i_0_1_635 (.A(n_0_1_649), .ZN(n_0_1_648));
   AOI222_X1 i_0_1_636 (.A1(n_0_1_256), .A2(n_0_1_730), .B1(n_0_1_269), .B2(
      n_0_1_728), .C1(n_0_1_727), .C2(n_0_1_650), .ZN(n_0_1_649));
   INV_X1 i_0_1_637 (.A(n_0_1_651), .ZN(n_0_1_650));
   AOI222_X1 i_0_1_638 (.A1(n_0_1_231), .A2(n_0_1_739), .B1(n_0_1_244), .B2(
      n_0_1_741), .C1(n_0_1_738), .C2(n_0_1_652), .ZN(n_0_1_651));
   INV_X1 i_0_1_639 (.A(n_0_1_653), .ZN(n_0_1_652));
   AOI222_X1 i_0_1_640 (.A1(n_0_1_206), .A2(n_0_1_751), .B1(n_0_1_219), .B2(
      n_0_1_753), .C1(n_0_1_750), .C2(n_0_1_654), .ZN(n_0_1_653));
   OAI21_X1 i_0_1_641 (.A(n_0_1_655), .B1(n_0_1_766), .B2(n_0_1_658), .ZN(
      n_0_1_654));
   AOI21_X1 i_0_1_642 (.A(n_0_1_761), .B1(n_0_1_763), .B2(n_0_1_656), .ZN(
      n_0_1_655));
   XOR2_X1 i_0_1_643 (.A(n_0_1_771), .B(n_0_1_657), .Z(n_0_1_656));
   OAI22_X1 i_0_1_644 (.A1(in_a[14]), .A2(n_0_1_812), .B1(n_0_1_813), .B2(
      n_0_1_15), .ZN(n_0_1_657));
   OAI21_X1 i_0_1_645 (.A(n_0_1_659), .B1(n_0_1_25), .B2(n_0_1_660), .ZN(
      n_0_1_658));
   NAND2_X1 i_0_1_646 (.A1(n_0_1_25), .A2(n_0_1_660), .ZN(n_0_1_659));
   AOI21_X1 i_0_1_647 (.A(n_0_1_770), .B1(n_0_459), .B2(n_0_1_769), .ZN(
      n_0_1_660));
   INV_X1 i_0_1_648 (.A(n_0_1_661), .ZN(n_0_439));
   AOI222_X1 i_0_1_649 (.A1(n_0_1_307), .A2(n_0_1_705), .B1(n_0_1_320), .B2(
      n_0_1_707), .C1(n_0_1_704), .C2(n_0_1_662), .ZN(n_0_1_661));
   INV_X1 i_0_1_650 (.A(n_0_1_663), .ZN(n_0_1_662));
   AOI222_X1 i_0_1_651 (.A1(n_0_1_282), .A2(n_0_1_717), .B1(n_0_1_295), .B2(
      n_0_1_719), .C1(n_0_1_716), .C2(n_0_1_664), .ZN(n_0_1_663));
   INV_X1 i_0_1_652 (.A(n_0_1_665), .ZN(n_0_1_664));
   AOI222_X1 i_0_1_653 (.A1(n_0_1_257), .A2(n_0_1_730), .B1(n_0_1_270), .B2(
      n_0_1_728), .C1(n_0_1_727), .C2(n_0_1_666), .ZN(n_0_1_665));
   INV_X1 i_0_1_654 (.A(n_0_1_667), .ZN(n_0_1_666));
   AOI222_X1 i_0_1_655 (.A1(n_0_1_232), .A2(n_0_1_739), .B1(n_0_1_245), .B2(
      n_0_1_741), .C1(n_0_1_738), .C2(n_0_1_668), .ZN(n_0_1_667));
   INV_X1 i_0_1_656 (.A(n_0_1_669), .ZN(n_0_1_668));
   AOI221_X1 i_0_1_657 (.A(n_0_1_749), .B1(n_0_1_751), .B2(n_0_1_670), .C1(
      n_0_1_753), .C2(n_0_1_672), .ZN(n_0_1_669));
   XOR2_X1 i_0_1_658 (.A(n_0_1_756), .B(n_0_1_671), .Z(n_0_1_670));
   OAI22_X1 i_0_1_659 (.A1(in_a[14]), .A2(n_0_1_811), .B1(n_0_1_813), .B2(
      n_0_1_38), .ZN(n_0_1_671));
   XOR2_X1 i_0_1_660 (.A(n_0_1_756), .B(n_0_1_673), .Z(n_0_1_672));
   OAI22_X1 i_0_1_661 (.A1(n_0_1_810), .A2(n_0_458), .B1(n_0_1_51), .B2(
      n_0_1_774), .ZN(n_0_1_673));
   INV_X1 i_0_1_662 (.A(n_0_1_674), .ZN(n_0_440));
   AOI222_X1 i_0_1_663 (.A1(n_0_1_308), .A2(n_0_1_705), .B1(n_0_1_321), .B2(
      n_0_1_707), .C1(n_0_1_704), .C2(n_0_1_675), .ZN(n_0_1_674));
   INV_X1 i_0_1_664 (.A(n_0_1_676), .ZN(n_0_1_675));
   AOI222_X1 i_0_1_665 (.A1(n_0_1_283), .A2(n_0_1_717), .B1(n_0_1_296), .B2(
      n_0_1_719), .C1(n_0_1_716), .C2(n_0_1_677), .ZN(n_0_1_676));
   INV_X1 i_0_1_666 (.A(n_0_1_678), .ZN(n_0_1_677));
   AOI222_X1 i_0_1_667 (.A1(n_0_1_258), .A2(n_0_1_730), .B1(n_0_1_271), .B2(
      n_0_1_728), .C1(n_0_1_727), .C2(n_0_1_679), .ZN(n_0_1_678));
   XOR2_X1 i_0_1_668 (.A(n_0_1_745), .B(n_0_1_680), .Z(n_0_1_679));
   AOI22_X1 i_0_1_669 (.A1(n_0_1_739), .A2(n_0_1_682), .B1(n_0_1_741), .B2(
      n_0_1_681), .ZN(n_0_1_680));
   OAI22_X1 i_0_1_670 (.A1(n_0_1_808), .A2(n_0_458), .B1(n_0_1_77), .B2(
      n_0_1_774), .ZN(n_0_1_681));
   OAI22_X1 i_0_1_671 (.A1(in_a[14]), .A2(n_0_1_809), .B1(n_0_1_813), .B2(
      n_0_1_64), .ZN(n_0_1_682));
   INV_X1 i_0_1_672 (.A(n_0_1_683), .ZN(n_0_441));
   AOI222_X1 i_0_1_673 (.A1(n_0_1_309), .A2(n_0_1_705), .B1(n_0_1_322), .B2(
      n_0_1_707), .C1(n_0_1_704), .C2(n_0_1_684), .ZN(n_0_1_683));
   INV_X1 i_0_1_674 (.A(n_0_1_685), .ZN(n_0_1_684));
   AOI222_X1 i_0_1_675 (.A1(n_0_1_284), .A2(n_0_1_717), .B1(n_0_1_297), .B2(
      n_0_1_719), .C1(n_0_1_716), .C2(n_0_1_686), .ZN(n_0_1_685));
   XNOR2_X1 i_0_1_676 (.A(n_0_1_733), .B(n_0_1_687), .ZN(n_0_1_686));
   AOI22_X1 i_0_1_677 (.A1(n_0_1_730), .A2(n_0_1_689), .B1(n_0_1_728), .B2(
      n_0_1_688), .ZN(n_0_1_687));
   OAI22_X1 i_0_1_678 (.A1(n_0_1_806), .A2(n_0_458), .B1(n_0_1_103), .B2(
      n_0_1_774), .ZN(n_0_1_688));
   OAI22_X1 i_0_1_679 (.A1(in_a[14]), .A2(n_0_1_807), .B1(n_0_1_813), .B2(
      n_0_1_90), .ZN(n_0_1_689));
   INV_X1 i_0_1_680 (.A(n_0_1_690), .ZN(n_0_442));
   AOI222_X1 i_0_1_681 (.A1(n_0_1_310), .A2(n_0_1_705), .B1(n_0_1_323), .B2(
      n_0_1_707), .C1(n_0_1_704), .C2(n_0_1_691), .ZN(n_0_1_690));
   INV_X1 i_0_1_682 (.A(n_0_1_692), .ZN(n_0_1_691));
   AOI221_X1 i_0_1_683 (.A(n_0_1_715), .B1(n_0_1_717), .B2(n_0_1_693), .C1(
      n_0_1_719), .C2(n_0_1_695), .ZN(n_0_1_692));
   XOR2_X1 i_0_1_684 (.A(n_0_1_722), .B(n_0_1_694), .Z(n_0_1_693));
   OAI22_X1 i_0_1_685 (.A1(in_a[14]), .A2(n_0_1_805), .B1(n_0_1_813), .B2(
      n_0_1_116), .ZN(n_0_1_694));
   XOR2_X1 i_0_1_686 (.A(n_0_1_722), .B(n_0_1_696), .Z(n_0_1_695));
   OAI22_X1 i_0_1_687 (.A1(n_0_1_804), .A2(n_0_458), .B1(n_0_1_129), .B2(
      n_0_1_774), .ZN(n_0_1_696));
   XOR2_X1 i_0_1_688 (.A(n_0_1_711), .B(n_0_1_697), .Z(n_0_443));
   AOI22_X1 i_0_1_689 (.A1(n_0_1_705), .A2(n_0_1_699), .B1(n_0_1_707), .B2(
      n_0_1_698), .ZN(n_0_1_697));
   OAI22_X1 i_0_1_690 (.A1(n_0_1_802), .A2(n_0_458), .B1(n_0_1_155), .B2(
      n_0_1_774), .ZN(n_0_1_698));
   OAI22_X1 i_0_1_691 (.A1(in_a[14]), .A2(n_0_1_803), .B1(n_0_1_813), .B2(
      n_0_1_142), .ZN(n_0_1_699));
   INV_X1 i_0_1_692 (.A(n_0_1_700), .ZN(n_0_444));
   AOI222_X1 i_0_1_693 (.A1(n_0_1_710), .A2(n_0_1_704), .B1(n_0_1_705), .B2(
      n_0_1_701), .C1(n_0_1_707), .C2(n_0_1_706), .ZN(n_0_1_700));
   XOR2_X1 i_0_1_694 (.A(n_0_1_772), .B(n_0_1_702), .Z(n_0_1_701));
   AOI21_X1 i_0_1_695 (.A(n_0_1_703), .B1(n_0_1_813), .B2(n_0_1_142), .ZN(
      n_0_1_702));
   AOI21_X1 i_0_1_696 (.A(n_0_1_710), .B1(in_a[14]), .B2(n_0_1_803), .ZN(
      n_0_1_703));
   NOR2_X1 i_0_1_697 (.A1(n_0_1_707), .A2(n_0_1_705), .ZN(n_0_1_704));
   NOR2_X1 i_0_1_698 (.A1(in_b[6]), .A2(n_0_1_818), .ZN(n_0_1_705));
   XOR2_X1 i_0_1_699 (.A(n_0_1_773), .B(n_0_1_708), .Z(n_0_1_706));
   NOR2_X1 i_0_1_700 (.A1(n_0_1_819), .A2(in_b[5]), .ZN(n_0_1_707));
   AOI21_X1 i_0_1_701 (.A(n_0_1_709), .B1(n_0_1_155), .B2(n_0_1_774), .ZN(
      n_0_1_708));
   AOI21_X1 i_0_1_702 (.A(n_0_1_710), .B1(n_0_1_802), .B2(n_0_458), .ZN(
      n_0_1_709));
   INV_X1 i_0_1_703 (.A(n_0_1_711), .ZN(n_0_1_710));
   AOI221_X1 i_0_1_704 (.A(n_0_1_715), .B1(n_0_1_717), .B2(n_0_1_712), .C1(
      n_0_1_719), .C2(n_0_1_718), .ZN(n_0_1_711));
   XOR2_X1 i_0_1_705 (.A(n_0_1_772), .B(n_0_1_713), .Z(n_0_1_712));
   AOI21_X1 i_0_1_706 (.A(n_0_1_714), .B1(n_0_1_813), .B2(n_0_1_116), .ZN(
      n_0_1_713));
   AOI21_X1 i_0_1_707 (.A(n_0_1_722), .B1(in_a[14]), .B2(n_0_1_805), .ZN(
      n_0_1_714));
   AND2_X1 i_0_1_708 (.A1(n_0_1_722), .A2(n_0_1_716), .ZN(n_0_1_715));
   NOR2_X1 i_0_1_709 (.A1(n_0_1_719), .A2(n_0_1_717), .ZN(n_0_1_716));
   NOR2_X1 i_0_1_710 (.A1(in_b[5]), .A2(n_0_1_817), .ZN(n_0_1_717));
   XOR2_X1 i_0_1_711 (.A(n_0_1_773), .B(n_0_1_720), .Z(n_0_1_718));
   NOR2_X1 i_0_1_712 (.A1(n_0_1_818), .A2(in_b[4]), .ZN(n_0_1_719));
   AOI21_X1 i_0_1_713 (.A(n_0_1_721), .B1(n_0_1_129), .B2(n_0_1_774), .ZN(
      n_0_1_720));
   AOI21_X1 i_0_1_714 (.A(n_0_1_722), .B1(n_0_1_804), .B2(n_0_458), .ZN(
      n_0_1_721));
   INV_X1 i_0_1_715 (.A(n_0_1_723), .ZN(n_0_1_722));
   AOI222_X1 i_0_1_716 (.A1(n_0_1_733), .A2(n_0_1_727), .B1(n_0_1_728), .B2(
      n_0_1_724), .C1(n_0_1_730), .C2(n_0_1_729), .ZN(n_0_1_723));
   XOR2_X1 i_0_1_717 (.A(n_0_1_773), .B(n_0_1_725), .Z(n_0_1_724));
   AOI21_X1 i_0_1_718 (.A(n_0_1_726), .B1(n_0_1_103), .B2(n_0_1_774), .ZN(
      n_0_1_725));
   AOI21_X1 i_0_1_719 (.A(n_0_1_733), .B1(n_0_1_806), .B2(n_0_458), .ZN(
      n_0_1_726));
   NOR2_X1 i_0_1_720 (.A1(n_0_1_730), .A2(n_0_1_728), .ZN(n_0_1_727));
   NOR2_X1 i_0_1_721 (.A1(n_0_1_817), .A2(in_b[3]), .ZN(n_0_1_728));
   XOR2_X1 i_0_1_722 (.A(n_0_1_772), .B(n_0_1_731), .Z(n_0_1_729));
   NOR2_X1 i_0_1_723 (.A1(in_b[4]), .A2(n_0_1_816), .ZN(n_0_1_730));
   AOI21_X1 i_0_1_724 (.A(n_0_1_732), .B1(n_0_1_813), .B2(n_0_1_90), .ZN(
      n_0_1_731));
   AOI21_X1 i_0_1_725 (.A(n_0_1_733), .B1(in_a[14]), .B2(n_0_1_807), .ZN(
      n_0_1_732));
   INV_X1 i_0_1_726 (.A(n_0_1_734), .ZN(n_0_1_733));
   AOI222_X1 i_0_1_727 (.A1(n_0_1_744), .A2(n_0_1_738), .B1(n_0_1_739), .B2(
      n_0_1_735), .C1(n_0_1_741), .C2(n_0_1_740), .ZN(n_0_1_734));
   XOR2_X1 i_0_1_728 (.A(n_0_1_772), .B(n_0_1_736), .Z(n_0_1_735));
   AOI21_X1 i_0_1_729 (.A(n_0_1_737), .B1(n_0_1_813), .B2(n_0_1_64), .ZN(
      n_0_1_736));
   AOI21_X1 i_0_1_730 (.A(n_0_1_744), .B1(in_a[14]), .B2(n_0_1_809), .ZN(
      n_0_1_737));
   NOR2_X1 i_0_1_731 (.A1(n_0_1_741), .A2(n_0_1_739), .ZN(n_0_1_738));
   NOR2_X1 i_0_1_732 (.A1(in_b[3]), .A2(n_0_1_815), .ZN(n_0_1_739));
   XOR2_X1 i_0_1_733 (.A(n_0_1_773), .B(n_0_1_742), .Z(n_0_1_740));
   NOR2_X1 i_0_1_734 (.A1(n_0_1_816), .A2(in_b[2]), .ZN(n_0_1_741));
   AOI21_X1 i_0_1_735 (.A(n_0_1_743), .B1(n_0_1_77), .B2(n_0_1_774), .ZN(
      n_0_1_742));
   AOI21_X1 i_0_1_736 (.A(n_0_1_744), .B1(n_0_1_808), .B2(n_0_458), .ZN(
      n_0_1_743));
   INV_X1 i_0_1_737 (.A(n_0_1_745), .ZN(n_0_1_744));
   AOI221_X1 i_0_1_738 (.A(n_0_1_749), .B1(n_0_1_751), .B2(n_0_1_746), .C1(
      n_0_1_753), .C2(n_0_1_752), .ZN(n_0_1_745));
   XOR2_X1 i_0_1_739 (.A(n_0_1_772), .B(n_0_1_747), .Z(n_0_1_746));
   AOI21_X1 i_0_1_740 (.A(n_0_1_748), .B1(n_0_1_813), .B2(n_0_1_38), .ZN(
      n_0_1_747));
   AOI21_X1 i_0_1_741 (.A(n_0_1_756), .B1(in_a[14]), .B2(n_0_1_811), .ZN(
      n_0_1_748));
   AND2_X1 i_0_1_742 (.A1(n_0_1_756), .A2(n_0_1_750), .ZN(n_0_1_749));
   NOR2_X1 i_0_1_743 (.A1(n_0_1_753), .A2(n_0_1_751), .ZN(n_0_1_750));
   AND2_X1 i_0_1_744 (.A1(n_0_1_815), .A2(in_b[1]), .ZN(n_0_1_751));
   XOR2_X1 i_0_1_745 (.A(n_0_1_773), .B(n_0_1_754), .Z(n_0_1_752));
   NOR2_X1 i_0_1_746 (.A1(n_0_1_815), .A2(in_b[1]), .ZN(n_0_1_753));
   AOI21_X1 i_0_1_747 (.A(n_0_1_755), .B1(n_0_1_51), .B2(n_0_1_774), .ZN(
      n_0_1_754));
   AOI21_X1 i_0_1_748 (.A(n_0_1_756), .B1(n_0_1_810), .B2(n_0_458), .ZN(
      n_0_1_755));
   INV_X1 i_0_1_749 (.A(n_0_1_757), .ZN(n_0_1_756));
   AOI221_X1 i_0_1_750 (.A(n_0_1_761), .B1(n_0_1_763), .B2(n_0_1_758), .C1(
      n_0_1_765), .C2(n_0_1_764), .ZN(n_0_1_757));
   XOR2_X1 i_0_1_751 (.A(n_0_1_772), .B(n_0_1_759), .Z(n_0_1_758));
   OAI21_X1 i_0_1_752 (.A(n_0_1_760), .B1(n_0_1_813), .B2(n_0_1_15), .ZN(
      n_0_1_759));
   OAI21_X1 i_0_1_753 (.A(n_0_1_771), .B1(in_a[14]), .B2(n_0_1_812), .ZN(
      n_0_1_760));
   AND2_X1 i_0_1_754 (.A1(n_0_1_771), .A2(n_0_1_762), .ZN(n_0_1_761));
   NOR2_X1 i_0_1_755 (.A1(n_0_1_765), .A2(n_0_1_763), .ZN(n_0_1_762));
   NOR2_X1 i_0_1_756 (.A1(in_b[1]), .A2(n_0_1_814), .ZN(n_0_1_763));
   XOR2_X1 i_0_1_757 (.A(n_0_1_773), .B(n_0_1_767), .Z(n_0_1_764));
   INV_X1 i_0_1_758 (.A(n_0_1_766), .ZN(n_0_1_765));
   NAND2_X1 i_0_1_759 (.A1(in_b[1]), .A2(n_0_1_814), .ZN(n_0_1_766));
   AOI21_X1 i_0_1_760 (.A(n_0_1_770), .B1(n_0_1_25), .B2(n_0_1_768), .ZN(
      n_0_1_767));
   NAND2_X1 i_0_1_761 (.A1(n_0_459), .A2(n_0_1_769), .ZN(n_0_1_768));
   NOR2_X1 i_0_1_762 (.A1(n_0_1_814), .A2(n_0_1_774), .ZN(n_0_1_769));
   NOR2_X1 i_0_1_763 (.A1(n_0_458), .A2(n_0_1_771), .ZN(n_0_1_770));
   AND2_X1 i_0_1_764 (.A1(in_b[0]), .A2(n_0_459), .ZN(n_0_1_771));
   XNOR2_X1 i_0_1_765 (.A(in_a[15]), .B(n_0_1_813), .ZN(n_0_1_772));
   XNOR2_X1 i_0_1_766 (.A(in_a[15]), .B(n_0_1_775), .ZN(n_0_1_773));
   AOI21_X1 i_0_1_767 (.A(n_0_1_801), .B1(in_a[1]), .B2(in_a[0]), .ZN(n_0_445));
   AOI21_X1 i_0_1_768 (.A(n_0_1_799), .B1(in_a[2]), .B2(n_0_1_800), .ZN(n_0_446));
   AOI21_X1 i_0_1_769 (.A(n_0_1_797), .B1(in_a[3]), .B2(n_0_1_798), .ZN(n_0_447));
   AOI21_X1 i_0_1_770 (.A(n_0_1_795), .B1(in_a[4]), .B2(n_0_1_796), .ZN(n_0_448));
   AOI21_X1 i_0_1_771 (.A(n_0_1_793), .B1(in_a[5]), .B2(n_0_1_794), .ZN(n_0_449));
   AOI21_X1 i_0_1_772 (.A(n_0_1_791), .B1(in_a[6]), .B2(n_0_1_792), .ZN(n_0_450));
   AOI21_X1 i_0_1_773 (.A(n_0_1_789), .B1(in_a[7]), .B2(n_0_1_790), .ZN(n_0_451));
   AOI21_X1 i_0_1_774 (.A(n_0_1_787), .B1(in_a[8]), .B2(n_0_1_788), .ZN(n_0_452));
   AOI21_X1 i_0_1_775 (.A(n_0_1_785), .B1(in_a[9]), .B2(n_0_1_786), .ZN(n_0_453));
   AOI21_X1 i_0_1_776 (.A(n_0_1_783), .B1(in_a[10]), .B2(n_0_1_784), .ZN(n_0_454));
   AOI21_X1 i_0_1_777 (.A(n_0_1_781), .B1(in_a[11]), .B2(n_0_1_782), .ZN(n_0_455));
   AOI21_X1 i_0_1_778 (.A(n_0_1_779), .B1(in_a[12]), .B2(n_0_1_780), .ZN(n_0_456));
   AOI21_X1 i_0_1_779 (.A(n_0_1_777), .B1(in_a[13]), .B2(n_0_1_778), .ZN(n_0_457));
   INV_X1 i_0_1_780 (.A(n_0_1_774), .ZN(n_0_458));
   NAND2_X1 i_0_1_781 (.A1(n_0_1_776), .A2(n_0_1_775), .ZN(n_0_1_774));
   OAI21_X1 i_0_1_782 (.A(in_a[14]), .B1(in_a[13]), .B2(n_0_1_778), .ZN(
      n_0_1_775));
   XOR2_X1 i_0_1_783 (.A(in_a[15]), .B(n_0_1_776), .Z(n_0_459));
   NAND2_X1 i_0_1_784 (.A1(n_0_1_813), .A2(n_0_1_777), .ZN(n_0_1_776));
   NOR2_X1 i_0_1_785 (.A1(in_a[13]), .A2(n_0_1_778), .ZN(n_0_1_777));
   INV_X1 i_0_1_786 (.A(n_0_1_779), .ZN(n_0_1_778));
   NOR2_X1 i_0_1_787 (.A1(in_a[12]), .A2(n_0_1_780), .ZN(n_0_1_779));
   INV_X1 i_0_1_788 (.A(n_0_1_781), .ZN(n_0_1_780));
   NOR2_X1 i_0_1_789 (.A1(in_a[11]), .A2(n_0_1_782), .ZN(n_0_1_781));
   INV_X1 i_0_1_790 (.A(n_0_1_783), .ZN(n_0_1_782));
   NOR2_X1 i_0_1_791 (.A1(in_a[10]), .A2(n_0_1_784), .ZN(n_0_1_783));
   INV_X1 i_0_1_792 (.A(n_0_1_785), .ZN(n_0_1_784));
   NOR2_X1 i_0_1_793 (.A1(in_a[9]), .A2(n_0_1_786), .ZN(n_0_1_785));
   INV_X1 i_0_1_794 (.A(n_0_1_787), .ZN(n_0_1_786));
   NOR2_X1 i_0_1_795 (.A1(in_a[8]), .A2(n_0_1_788), .ZN(n_0_1_787));
   INV_X1 i_0_1_796 (.A(n_0_1_789), .ZN(n_0_1_788));
   NOR2_X1 i_0_1_797 (.A1(in_a[7]), .A2(n_0_1_790), .ZN(n_0_1_789));
   INV_X1 i_0_1_798 (.A(n_0_1_791), .ZN(n_0_1_790));
   NOR2_X1 i_0_1_799 (.A1(in_a[6]), .A2(n_0_1_792), .ZN(n_0_1_791));
   INV_X1 i_0_1_800 (.A(n_0_1_793), .ZN(n_0_1_792));
   NOR2_X1 i_0_1_801 (.A1(in_a[5]), .A2(n_0_1_794), .ZN(n_0_1_793));
   INV_X1 i_0_1_802 (.A(n_0_1_795), .ZN(n_0_1_794));
   NOR2_X1 i_0_1_803 (.A1(in_a[4]), .A2(n_0_1_796), .ZN(n_0_1_795));
   INV_X1 i_0_1_804 (.A(n_0_1_797), .ZN(n_0_1_796));
   NOR2_X1 i_0_1_805 (.A1(in_a[3]), .A2(n_0_1_798), .ZN(n_0_1_797));
   INV_X1 i_0_1_806 (.A(n_0_1_799), .ZN(n_0_1_798));
   NOR2_X1 i_0_1_807 (.A1(in_a[2]), .A2(n_0_1_800), .ZN(n_0_1_799));
   INV_X1 i_0_1_808 (.A(n_0_1_801), .ZN(n_0_1_800));
   NOR2_X1 i_0_1_809 (.A1(in_a[1]), .A2(in_a[0]), .ZN(n_0_1_801));
   INV_X1 i_0_1_810 (.A(n_0_1_155), .ZN(n_0_1_802));
   INV_X1 i_0_1_811 (.A(n_0_1_142), .ZN(n_0_1_803));
   INV_X1 i_0_1_812 (.A(n_0_1_129), .ZN(n_0_1_804));
   INV_X1 i_0_1_813 (.A(n_0_1_116), .ZN(n_0_1_805));
   INV_X1 i_0_1_814 (.A(n_0_1_103), .ZN(n_0_1_806));
   INV_X1 i_0_1_815 (.A(n_0_1_90), .ZN(n_0_1_807));
   INV_X1 i_0_1_816 (.A(n_0_1_77), .ZN(n_0_1_808));
   INV_X1 i_0_1_817 (.A(n_0_1_64), .ZN(n_0_1_809));
   INV_X1 i_0_1_818 (.A(n_0_1_51), .ZN(n_0_1_810));
   INV_X1 i_0_1_819 (.A(n_0_1_38), .ZN(n_0_1_811));
   INV_X1 i_0_1_820 (.A(n_0_1_15), .ZN(n_0_1_812));
   INV_X1 i_0_1_821 (.A(in_a[14]), .ZN(n_0_1_813));
   INV_X1 i_0_1_822 (.A(in_b[0]), .ZN(n_0_1_814));
   INV_X1 i_0_1_823 (.A(in_b[2]), .ZN(n_0_1_815));
   INV_X1 i_0_1_824 (.A(in_b[3]), .ZN(n_0_1_816));
   INV_X1 i_0_1_825 (.A(in_b[4]), .ZN(n_0_1_817));
   INV_X1 i_0_1_826 (.A(in_b[5]), .ZN(n_0_1_818));
   INV_X1 i_0_1_827 (.A(in_b[6]), .ZN(n_0_1_819));
   INV_X1 i_0_1_828 (.A(in_b[7]), .ZN(n_0_1_820));
   INV_X1 i_0_1_829 (.A(in_b[8]), .ZN(n_0_1_821));
   INV_X1 i_0_1_830 (.A(in_b[9]), .ZN(n_0_1_822));
   INV_X1 i_0_1_831 (.A(in_b[10]), .ZN(n_0_1_823));
   INV_X1 i_0_1_832 (.A(in_b[11]), .ZN(n_0_1_824));
   INV_X1 i_0_1_833 (.A(in_b[12]), .ZN(n_0_1_825));
   INV_X1 i_0_1_834 (.A(in_b[13]), .ZN(n_0_1_826));
   INV_X1 i_0_1_835 (.A(in_b[14]), .ZN(n_0_1_827));
   NOR2_X1 i_0_2_0 (.A1(n_0_2_0), .A2(error), .ZN(n_0_460));
   AOI21_X1 i_0_2_1 (.A(rst), .B1(n_0_464), .B2(n_0_2_0), .ZN(n_0_463));
   NOR2_X1 i_0_2_2 (.A1(n_0_2_0), .A2(rst), .ZN(n_0_462));
   OR2_X1 i_0_2_3 (.A1(n_0_464), .A2(n_0_461), .ZN(n_0_465));
   OR2_X1 i_0_2_4 (.A1(rst), .A2(enbl), .ZN(n_0_461));
   INV_X1 i_0_2_5 (.A(enbl), .ZN(n_0_2_0));
   INV_X1 i_0_2_6 (.A(error), .ZN(n_0_464));
endmodule
